magic
tech sky130A
magscale 1 2
timestamp 1636369236
<< error_p >>
rect -907 562 -761 600
rect -907 536 -857 562
rect -907 530 1025 536
rect -927 494 989 500
rect -1147 -380 -1025 -346
rect -1147 -490 -599 -380
rect -1147 -500 989 -490
rect -1147 -514 -599 -500
rect -1025 -526 -599 -514
rect -1025 -536 985 -526
rect -1025 -552 -857 -536
rect -853 -552 -685 -536
rect -1025 -600 -685 -552
rect 1025 -562 1153 -358
rect -979 -634 -853 -600
rect -941 -667 -883 -661
rect -941 -701 -929 -667
rect -941 -707 -883 -701
rect -853 -720 -811 -634
<< nwell >>
rect -929 562 -907 600
rect -1025 530 -907 562
rect -1025 -514 1025 530
rect -1025 -600 -979 -514
rect -853 -526 1025 -514
rect -853 -600 -785 -526
rect 985 -562 1025 -526
rect -979 -720 -853 -634
<< pmos >>
rect -927 -500 -897 500
rect -831 -500 -801 500
rect -735 -500 -705 500
rect -639 -500 -609 500
rect -543 -500 -513 500
rect -447 -500 -417 500
rect -351 -500 -321 500
rect -255 -500 -225 500
rect -159 -500 -129 500
rect -63 -500 -33 500
rect 33 -500 63 500
rect 129 -500 159 500
rect 225 -500 255 500
rect 321 -500 351 500
rect 417 -500 447 500
rect 513 -500 543 500
rect 609 -500 639 500
rect 705 -500 735 500
rect 801 -500 831 500
rect 897 -500 927 500
<< pdiff >>
rect -989 488 -927 500
rect -989 -488 -977 488
rect -943 -488 -927 488
rect -989 -500 -927 -488
rect -897 488 -831 500
rect -897 -488 -881 488
rect -847 -488 -831 488
rect -897 -500 -831 -488
rect -801 488 -735 500
rect -801 -488 -785 488
rect -751 -488 -735 488
rect -801 -500 -735 -488
rect -705 488 -639 500
rect -705 -488 -689 488
rect -655 -488 -639 488
rect -705 -500 -639 -488
rect -609 488 -543 500
rect -609 -488 -593 488
rect -559 -488 -543 488
rect -609 -500 -543 -488
rect -513 488 -447 500
rect -513 -488 -497 488
rect -463 -488 -447 488
rect -513 -500 -447 -488
rect -417 488 -351 500
rect -417 -488 -401 488
rect -367 -488 -351 488
rect -417 -500 -351 -488
rect -321 488 -255 500
rect -321 -488 -305 488
rect -271 -488 -255 488
rect -321 -500 -255 -488
rect -225 488 -159 500
rect -225 -488 -209 488
rect -175 -488 -159 488
rect -225 -500 -159 -488
rect -129 488 -63 500
rect -129 -488 -113 488
rect -79 -488 -63 488
rect -129 -500 -63 -488
rect -33 488 33 500
rect -33 -488 -17 488
rect 17 -488 33 488
rect -33 -500 33 -488
rect 63 488 129 500
rect 63 -488 79 488
rect 113 -488 129 488
rect 63 -500 129 -488
rect 159 488 225 500
rect 159 -488 175 488
rect 209 -488 225 488
rect 159 -500 225 -488
rect 255 488 321 500
rect 255 -488 271 488
rect 305 -488 321 488
rect 255 -500 321 -488
rect 351 488 417 500
rect 351 -488 367 488
rect 401 -488 417 488
rect 351 -500 417 -488
rect 447 488 513 500
rect 447 -488 463 488
rect 497 -488 513 488
rect 447 -500 513 -488
rect 543 488 609 500
rect 543 -488 559 488
rect 593 -488 609 488
rect 543 -500 609 -488
rect 639 488 705 500
rect 639 -488 655 488
rect 689 -488 705 488
rect 639 -500 705 -488
rect 735 488 801 500
rect 735 -488 751 488
rect 785 -488 801 488
rect 735 -500 801 -488
rect 831 488 897 500
rect 831 -488 847 488
rect 881 -488 897 488
rect 831 -500 897 -488
rect 927 488 989 500
rect 927 -488 943 488
rect 977 -488 989 488
rect 927 -500 989 -488
<< pdiffc >>
rect -977 -488 -943 488
rect -881 -488 -847 488
rect -785 -488 -751 488
rect -689 -488 -655 488
rect -593 -488 -559 488
rect -497 -488 -463 488
rect -401 -488 -367 488
rect -305 -488 -271 488
rect -209 -488 -175 488
rect -113 -488 -79 488
rect -17 -488 17 488
rect 79 -488 113 488
rect 175 -488 209 488
rect 271 -488 305 488
rect 367 -488 401 488
rect 463 -488 497 488
rect 559 -488 593 488
rect 655 -488 689 488
rect 751 -488 785 488
rect 847 -488 881 488
rect 943 -488 977 488
<< poly >>
rect -927 500 -897 526
rect -831 500 -801 530
rect -735 500 -705 526
rect -639 500 -609 530
rect -543 500 -513 526
rect -447 500 -417 530
rect -351 500 -321 526
rect -255 500 -225 530
rect -159 500 -129 526
rect -63 500 -33 530
rect 33 500 63 526
rect 129 500 159 530
rect 225 500 255 526
rect 321 500 351 530
rect 417 500 447 526
rect 513 500 543 530
rect 609 500 639 526
rect 705 500 735 530
rect 801 500 831 526
rect 897 500 927 530
rect -927 -651 -897 -500
rect -831 -526 -801 -500
rect -735 -526 -705 -500
rect -639 -526 -609 -500
rect -543 -526 -513 -500
rect -447 -526 -417 -500
rect -351 -526 -321 -500
rect -255 -526 -225 -500
rect -159 -526 -129 -500
rect -63 -526 -33 -500
rect 33 -526 63 -500
rect 129 -526 159 -500
rect 225 -526 255 -500
rect 321 -526 351 -500
rect 417 -526 447 -500
rect 513 -526 543 -500
rect 609 -526 639 -500
rect 705 -526 735 -500
rect 801 -526 831 -500
rect 897 -526 927 -500
rect -945 -667 -879 -651
rect -945 -701 -929 -667
rect -895 -701 -879 -667
rect -945 -717 -879 -701
<< polycont >>
rect -929 -701 -895 -667
<< locali >>
rect -977 558 977 592
rect -977 488 -943 558
rect -977 -504 -943 -488
rect -881 488 -847 504
rect -881 -550 -847 -488
rect -785 488 -751 558
rect -785 -504 -751 -488
rect -689 488 -655 504
rect -689 -550 -655 -488
rect -593 488 -559 558
rect -593 -504 -559 -488
rect -497 488 -463 504
rect -497 -550 -463 -488
rect -401 488 -367 558
rect -401 -504 -367 -488
rect -305 488 -271 504
rect -305 -550 -271 -488
rect -209 488 -175 558
rect -209 -504 -175 -488
rect -113 488 -79 504
rect -113 -550 -79 -488
rect -17 488 17 558
rect -17 -504 17 -488
rect 79 488 113 504
rect 79 -550 113 -488
rect 175 488 209 558
rect 175 -504 209 -488
rect 271 488 305 504
rect 271 -550 305 -488
rect 367 488 401 558
rect 367 -504 401 -488
rect 463 488 497 504
rect 463 -550 497 -488
rect 559 488 593 558
rect 559 -504 593 -488
rect 655 488 689 504
rect 655 -550 689 -488
rect 751 488 785 558
rect 751 -504 785 -488
rect 847 488 881 504
rect 847 -550 881 -488
rect 943 488 977 558
rect 943 -504 977 -488
rect -881 -584 881 -550
rect -945 -701 -929 -667
rect -895 -701 -879 -667
<< viali >>
rect -977 -488 -943 488
rect -881 -488 -847 488
rect -785 -488 -751 488
rect -689 -488 -655 488
rect -593 -488 -559 488
rect -497 -488 -463 488
rect -401 -488 -367 488
rect -305 -488 -271 488
rect -209 -488 -175 488
rect -113 -488 -79 488
rect -17 -488 17 488
rect 79 -488 113 488
rect 175 -488 209 488
rect 271 -488 305 488
rect 367 -488 401 488
rect 463 -488 497 488
rect 559 -488 593 488
rect 655 -488 689 488
rect 751 -488 785 488
rect 847 -488 881 488
rect 943 -488 977 488
rect -929 -701 -895 -667
<< metal1 >>
rect -983 488 -937 500
rect -983 -488 -977 488
rect -943 -488 -937 488
rect -983 -500 -937 -488
rect -887 488 -841 500
rect -887 -488 -881 488
rect -847 -488 -841 488
rect -887 -500 -841 -488
rect -791 488 -745 500
rect -791 -488 -785 488
rect -751 -488 -745 488
rect -791 -500 -745 -488
rect -695 488 -649 500
rect -695 -488 -689 488
rect -655 -488 -649 488
rect -695 -500 -649 -488
rect -599 488 -553 500
rect -599 -488 -593 488
rect -559 -488 -553 488
rect -599 -500 -553 -488
rect -503 488 -457 500
rect -503 -488 -497 488
rect -463 -488 -457 488
rect -503 -500 -457 -488
rect -407 488 -361 500
rect -407 -488 -401 488
rect -367 -488 -361 488
rect -407 -500 -361 -488
rect -311 488 -265 500
rect -311 -488 -305 488
rect -271 -488 -265 488
rect -311 -500 -265 -488
rect -215 488 -169 500
rect -215 -488 -209 488
rect -175 -488 -169 488
rect -215 -500 -169 -488
rect -119 488 -73 500
rect -119 -488 -113 488
rect -79 -488 -73 488
rect -119 -500 -73 -488
rect -23 488 23 500
rect -23 -488 -17 488
rect 17 -488 23 488
rect -23 -500 23 -488
rect 73 488 119 500
rect 73 -488 79 488
rect 113 -488 119 488
rect 73 -500 119 -488
rect 169 488 215 500
rect 169 -488 175 488
rect 209 -488 215 488
rect 169 -500 215 -488
rect 265 488 311 500
rect 265 -488 271 488
rect 305 -488 311 488
rect 265 -500 311 -488
rect 361 488 407 500
rect 361 -488 367 488
rect 401 -488 407 488
rect 361 -500 407 -488
rect 457 488 503 500
rect 457 -488 463 488
rect 497 -488 503 488
rect 457 -500 503 -488
rect 553 488 599 500
rect 553 -488 559 488
rect 593 -488 599 488
rect 553 -500 599 -488
rect 649 488 695 500
rect 649 -488 655 488
rect 689 -488 695 488
rect 649 -500 695 -488
rect 745 488 791 500
rect 745 -488 751 488
rect 785 -488 791 488
rect 745 -500 791 -488
rect 841 488 887 500
rect 841 -488 847 488
rect 881 -488 887 488
rect 841 -500 887 -488
rect 937 488 983 500
rect 937 -488 943 488
rect 977 -488 983 488
rect 937 -500 983 -488
rect -941 -667 -883 -661
rect -941 -701 -929 -667
rect -895 -701 -883 -667
rect -941 -707 -883 -701
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string parameters w 5 l 0.15 m 1 nf 20 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
