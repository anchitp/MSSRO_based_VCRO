magic
tech sky130A
magscale 1 2
timestamp 1636291015
<< error_p >>
rect -221 -687 -163 -681
rect -221 -721 -209 -687
rect -221 -727 -163 -721
<< nwell >>
rect -305 -750 305 600
<< pmos >>
rect -207 -500 -177 500
rect -111 -500 -81 500
rect -15 -500 15 500
rect 81 -500 111 500
rect 177 -500 207 500
<< pdiff >>
rect -269 488 -207 500
rect -269 -488 -257 488
rect -223 -488 -207 488
rect -269 -500 -207 -488
rect -177 488 -111 500
rect -177 -488 -161 488
rect -127 -488 -111 488
rect -177 -500 -111 -488
rect -81 488 -15 500
rect -81 -488 -65 488
rect -31 -488 -15 488
rect -81 -500 -15 -488
rect 15 488 81 500
rect 15 -488 31 488
rect 65 -488 81 488
rect 15 -500 81 -488
rect 111 488 177 500
rect 111 -488 127 488
rect 161 -488 177 488
rect 111 -500 177 -488
rect 207 488 269 500
rect 207 -488 223 488
rect 257 -488 269 488
rect 207 -500 269 -488
<< pdiffc >>
rect -257 -488 -223 488
rect -161 -488 -127 488
rect -65 -488 -31 488
rect 31 -488 65 488
rect 127 -488 161 488
rect 223 -488 257 488
<< poly >>
rect -207 500 -177 526
rect -111 500 -81 528
rect -15 500 15 526
rect 81 500 111 528
rect 177 500 207 526
rect -207 -516 -177 -500
rect -111 -516 -81 -500
rect -15 -516 15 -500
rect 81 -516 111 -500
rect 177 -516 207 -500
rect -207 -546 207 -516
rect -207 -671 -177 -546
rect -225 -687 -159 -671
rect -225 -721 -209 -687
rect -175 -721 -159 -687
rect -225 -737 -159 -721
<< polycont >>
rect -209 -721 -175 -687
<< locali >>
rect -257 544 161 578
rect -257 488 -223 544
rect -257 -504 -223 -488
rect -161 488 -127 504
rect -161 -556 -127 -488
rect -65 488 -31 544
rect -65 -504 -31 -488
rect 31 488 65 504
rect 31 -556 65 -488
rect 127 488 161 544
rect 127 -504 161 -488
rect 223 488 257 504
rect 223 -556 257 -488
rect -163 -590 257 -556
rect -225 -721 -209 -687
rect -175 -721 -159 -687
<< viali >>
rect -257 -488 -223 488
rect -161 -488 -127 488
rect -65 -488 -31 488
rect 31 -488 65 488
rect 127 -488 161 488
rect 223 -488 257 488
rect -209 -721 -175 -687
<< metal1 >>
rect -263 488 -217 500
rect -263 -488 -257 488
rect -223 -488 -217 488
rect -263 -500 -217 -488
rect -167 488 -121 500
rect -167 -488 -161 488
rect -127 -488 -121 488
rect -167 -500 -121 -488
rect -71 488 -25 500
rect -71 -488 -65 488
rect -31 -488 -25 488
rect -71 -500 -25 -488
rect 25 488 71 500
rect 25 -488 31 488
rect 65 -488 71 488
rect 25 -500 71 -488
rect 121 488 167 500
rect 121 -488 127 488
rect 161 -488 167 488
rect 121 -500 167 -488
rect 217 488 263 500
rect 217 -488 223 488
rect 257 -488 263 488
rect 217 -500 263 -488
rect -221 -687 -163 -681
rect -221 -721 -209 -687
rect -175 -721 -163 -687
rect -221 -727 -163 -721
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string parameters w 5 l 0.15 m 1 nf 5 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
