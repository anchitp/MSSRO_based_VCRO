magic
tech sky130A
magscale 1 2
timestamp 1636292965
<< error_p >>
rect -447 562 -281 600
rect -447 536 -377 562
rect -447 526 509 536
rect 545 526 677 600
rect -483 490 509 500
rect -673 -392 -545 -358
rect -673 -490 -93 -392
rect -673 -500 507 -490
rect -673 -526 -93 -500
rect -545 -536 471 -526
rect -545 -552 -377 -536
rect -347 -552 -179 -536
rect -545 -600 -179 -552
rect 545 -562 639 -358
rect -505 -646 -347 -600
rect -461 -667 -403 -661
rect -461 -701 -449 -667
rect -461 -707 -403 -701
rect -347 -720 -337 -646
<< nwell >>
rect -449 562 -447 600
rect -545 526 -447 562
rect 509 526 545 600
rect -545 -526 545 526
rect -545 -600 -505 -526
rect -347 -600 -299 -526
rect 471 -562 545 -526
rect -505 -720 -347 -646
<< pmos >>
rect -447 -500 -417 500
rect -351 -500 -321 500
rect -255 -500 -225 500
rect -159 -500 -129 500
rect -63 -500 -33 500
rect 33 -500 63 500
rect 129 -500 159 500
rect 225 -500 255 500
rect 321 -500 351 500
rect 417 -500 447 500
<< pdiff >>
rect -509 488 -447 500
rect -509 -488 -497 488
rect -463 -488 -447 488
rect -509 -500 -447 -488
rect -417 488 -351 500
rect -417 -488 -401 488
rect -367 -488 -351 488
rect -417 -500 -351 -488
rect -321 488 -255 500
rect -321 -488 -305 488
rect -271 -488 -255 488
rect -321 -500 -255 -488
rect -225 488 -159 500
rect -225 -488 -209 488
rect -175 -488 -159 488
rect -225 -500 -159 -488
rect -129 488 -63 500
rect -129 -488 -113 488
rect -79 -488 -63 488
rect -129 -500 -63 -488
rect -33 488 33 500
rect -33 -488 -17 488
rect 17 -488 33 488
rect -33 -500 33 -488
rect 63 488 129 500
rect 63 -488 79 488
rect 113 -488 129 488
rect 63 -500 129 -488
rect 159 488 225 500
rect 159 -488 175 488
rect 209 -488 225 488
rect 159 -500 225 -488
rect 255 488 321 500
rect 255 -488 271 488
rect 305 -488 321 488
rect 255 -500 321 -488
rect 351 488 417 500
rect 351 -488 367 488
rect 401 -488 417 488
rect 351 -500 417 -488
rect 447 488 509 500
rect 447 -488 463 488
rect 497 -488 509 488
rect 447 -500 509 -488
<< pdiffc >>
rect -497 -488 -463 488
rect -401 -488 -367 488
rect -305 -488 -271 488
rect -209 -488 -175 488
rect -113 -488 -79 488
rect -17 -488 17 488
rect 79 -488 113 488
rect 175 -488 209 488
rect 271 -488 305 488
rect 367 -488 401 488
rect 463 -488 497 488
<< poly >>
rect -447 500 -417 526
rect -351 500 -321 526
rect -255 500 -225 526
rect -159 500 -129 526
rect -63 500 -33 526
rect 33 500 63 526
rect 129 500 159 526
rect 225 500 255 526
rect 321 500 351 526
rect 417 500 447 526
rect -447 -524 -417 -500
rect -351 -524 -321 -500
rect -255 -524 -225 -500
rect -159 -524 -129 -500
rect -63 -524 -33 -500
rect 33 -524 63 -500
rect 129 -524 159 -500
rect 225 -524 255 -500
rect 321 -524 351 -500
rect 417 -524 447 -500
rect -447 -554 447 -524
rect -447 -651 -417 -554
rect -465 -667 -399 -651
rect -465 -701 -449 -667
rect -415 -701 -399 -667
rect -465 -717 -399 -701
<< polycont >>
rect -449 -701 -415 -667
<< locali >>
rect -497 544 497 578
rect -497 488 -463 544
rect -497 -504 -463 -488
rect -401 488 -367 504
rect -401 -562 -367 -488
rect -305 488 -271 544
rect -305 -504 -271 -488
rect -209 488 -175 504
rect -209 -562 -175 -488
rect -113 488 -79 544
rect -113 -504 -79 -488
rect -17 488 17 504
rect -17 -562 17 -488
rect 79 488 113 544
rect 79 -504 113 -488
rect 175 488 209 504
rect 175 -562 209 -488
rect 271 488 305 544
rect 271 -504 305 -488
rect 367 488 401 504
rect 367 -562 401 -488
rect 463 488 497 544
rect 463 -504 497 -488
rect -401 -596 401 -562
rect -465 -701 -449 -667
rect -415 -701 -399 -667
<< viali >>
rect -497 -488 -463 488
rect -401 -488 -367 488
rect -305 -488 -271 488
rect -209 -488 -175 488
rect -113 -488 -79 488
rect -17 -488 17 488
rect 79 -488 113 488
rect 175 -488 209 488
rect 271 -488 305 488
rect 367 -488 401 488
rect 463 -488 497 488
rect -449 -701 -415 -667
<< metal1 >>
rect -503 488 -457 500
rect -503 -488 -497 488
rect -463 -488 -457 488
rect -503 -500 -457 -488
rect -407 488 -361 500
rect -407 -488 -401 488
rect -367 -488 -361 488
rect -407 -500 -361 -488
rect -311 488 -265 500
rect -311 -488 -305 488
rect -271 -488 -265 488
rect -311 -500 -265 -488
rect -215 488 -169 500
rect -215 -488 -209 488
rect -175 -488 -169 488
rect -215 -500 -169 -488
rect -119 488 -73 500
rect -119 -488 -113 488
rect -79 -488 -73 488
rect -119 -500 -73 -488
rect -23 488 23 500
rect -23 -488 -17 488
rect 17 -488 23 488
rect -23 -500 23 -488
rect 73 488 119 500
rect 73 -488 79 488
rect 113 -488 119 488
rect 73 -500 119 -488
rect 169 488 215 500
rect 169 -488 175 488
rect 209 -488 215 488
rect 169 -500 215 -488
rect 265 488 311 500
rect 265 -488 271 488
rect 305 -488 311 488
rect 265 -500 311 -488
rect 361 488 407 500
rect 361 -488 367 488
rect 401 -488 407 488
rect 361 -500 407 -488
rect 457 488 503 500
rect 457 -488 463 488
rect 497 -488 503 488
rect 457 -500 503 -488
rect -461 -667 -403 -661
rect -461 -701 -449 -667
rect -415 -701 -403 -667
rect -461 -707 -403 -701
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string parameters w 5 l 0.15 m 1 nf 10 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
