magic
tech sky130A
magscale 1 2
timestamp 1636296519
<< error_p >>
rect -605 672 -547 678
rect -605 638 -593 672
rect -605 632 -547 638
<< nmos >>
rect -687 -500 -657 500
rect -591 -500 -561 500
rect -495 -500 -465 500
rect -399 -500 -369 500
rect -303 -500 -273 500
rect -207 -500 -177 500
rect -111 -500 -81 500
rect -15 -500 15 500
rect 81 -500 111 500
rect 177 -500 207 500
rect 273 -500 303 500
rect 369 -500 399 500
rect 465 -500 495 500
rect 561 -500 591 500
rect 657 -500 687 500
<< ndiff >>
rect -749 488 -687 500
rect -749 -488 -737 488
rect -703 -488 -687 488
rect -749 -500 -687 -488
rect -657 488 -591 500
rect -657 -488 -641 488
rect -607 -488 -591 488
rect -657 -500 -591 -488
rect -561 488 -495 500
rect -561 -488 -545 488
rect -511 -488 -495 488
rect -561 -500 -495 -488
rect -465 488 -399 500
rect -465 -488 -449 488
rect -415 -488 -399 488
rect -465 -500 -399 -488
rect -369 488 -303 500
rect -369 -488 -353 488
rect -319 -488 -303 488
rect -369 -500 -303 -488
rect -273 488 -207 500
rect -273 -488 -257 488
rect -223 -488 -207 488
rect -273 -500 -207 -488
rect -177 488 -111 500
rect -177 -488 -161 488
rect -127 -488 -111 488
rect -177 -500 -111 -488
rect -81 488 -15 500
rect -81 -488 -65 488
rect -31 -488 -15 488
rect -81 -500 -15 -488
rect 15 488 81 500
rect 15 -488 31 488
rect 65 -488 81 488
rect 15 -500 81 -488
rect 111 488 177 500
rect 111 -488 127 488
rect 161 -488 177 488
rect 111 -500 177 -488
rect 207 488 273 500
rect 207 -488 223 488
rect 257 -488 273 488
rect 207 -500 273 -488
rect 303 488 369 500
rect 303 -488 319 488
rect 353 -488 369 488
rect 303 -500 369 -488
rect 399 488 465 500
rect 399 -488 415 488
rect 449 -488 465 488
rect 399 -500 465 -488
rect 495 488 561 500
rect 495 -488 511 488
rect 545 -488 561 488
rect 495 -500 561 -488
rect 591 488 657 500
rect 591 -488 607 488
rect 641 -488 657 488
rect 591 -500 657 -488
rect 687 488 749 500
rect 687 -488 703 488
rect 737 -488 749 488
rect 687 -500 749 -488
<< ndiffc >>
rect -737 -488 -703 488
rect -641 -488 -607 488
rect -545 -488 -511 488
rect -449 -488 -415 488
rect -353 -488 -319 488
rect -257 -488 -223 488
rect -161 -488 -127 488
rect -65 -488 -31 488
rect 31 -488 65 488
rect 127 -488 161 488
rect 223 -488 257 488
rect 319 -488 353 488
rect 415 -488 449 488
rect 511 -488 545 488
rect 607 -488 641 488
rect 703 -488 737 488
<< poly >>
rect -609 672 -543 688
rect -609 638 -593 672
rect -559 638 -543 672
rect -609 622 -543 638
rect -591 550 -561 622
rect -687 518 687 550
rect -687 500 -657 518
rect -591 500 -561 518
rect -495 500 -465 518
rect -399 500 -369 518
rect -303 500 -273 518
rect -207 500 -177 518
rect -111 500 -81 518
rect -15 500 15 518
rect 81 500 111 518
rect 177 500 207 518
rect 273 500 303 518
rect 369 500 399 518
rect 465 500 495 518
rect 561 500 591 518
rect 657 500 687 518
rect -687 -526 -657 -500
rect -591 -526 -561 -500
rect -495 -526 -465 -500
rect -399 -526 -369 -500
rect -303 -526 -273 -500
rect -207 -526 -177 -500
rect -111 -526 -81 -500
rect -15 -526 15 -500
rect 81 -526 111 -500
rect 177 -526 207 -500
rect 273 -526 303 -500
rect 369 -526 399 -500
rect 465 -526 495 -500
rect 561 -526 591 -500
rect 657 -526 687 -500
<< polycont >>
rect -593 638 -559 672
<< locali >>
rect -609 638 -593 672
rect -559 638 -543 672
rect -641 554 737 588
rect -737 488 -703 504
rect -737 -546 -703 -488
rect -641 488 -607 554
rect -641 -504 -607 -488
rect -545 488 -511 504
rect -545 -546 -511 -488
rect -449 488 -415 554
rect -449 -504 -415 -488
rect -353 488 -319 504
rect -353 -546 -319 -488
rect -257 488 -223 554
rect -257 -504 -223 -488
rect -161 488 -127 504
rect -161 -546 -127 -488
rect -65 488 -31 554
rect -65 -504 -31 -488
rect 31 488 65 504
rect 31 -546 65 -488
rect 127 488 161 554
rect 127 -504 161 -488
rect 223 488 257 504
rect 223 -546 257 -488
rect 319 488 353 554
rect 319 -504 353 -488
rect 415 488 449 504
rect 415 -546 449 -488
rect 511 488 545 554
rect 511 -504 545 -488
rect 607 488 641 504
rect 607 -546 641 -488
rect 703 488 737 554
rect 703 -504 737 -488
rect -737 -580 653 -546
<< viali >>
rect -593 638 -559 672
rect -737 -488 -703 488
rect -641 -488 -607 488
rect -545 -488 -511 488
rect -449 -488 -415 488
rect -353 -488 -319 488
rect -257 -488 -223 488
rect -161 -488 -127 488
rect -65 -488 -31 488
rect 31 -488 65 488
rect 127 -488 161 488
rect 223 -488 257 488
rect 319 -488 353 488
rect 415 -488 449 488
rect 511 -488 545 488
rect 607 -488 641 488
rect 703 -488 737 488
<< metal1 >>
rect -605 672 -547 678
rect -605 638 -593 672
rect -559 638 -547 672
rect -605 632 -547 638
rect -743 488 -697 500
rect -743 -488 -737 488
rect -703 -488 -697 488
rect -743 -500 -697 -488
rect -647 488 -601 500
rect -647 -488 -641 488
rect -607 -488 -601 488
rect -647 -500 -601 -488
rect -551 488 -505 500
rect -551 -488 -545 488
rect -511 -488 -505 488
rect -551 -500 -505 -488
rect -455 488 -409 500
rect -455 -488 -449 488
rect -415 -488 -409 488
rect -455 -500 -409 -488
rect -359 488 -313 500
rect -359 -488 -353 488
rect -319 -488 -313 488
rect -359 -500 -313 -488
rect -263 488 -217 500
rect -263 -488 -257 488
rect -223 -488 -217 488
rect -263 -500 -217 -488
rect -167 488 -121 500
rect -167 -488 -161 488
rect -127 -488 -121 488
rect -167 -500 -121 -488
rect -71 488 -25 500
rect -71 -488 -65 488
rect -31 -488 -25 488
rect -71 -500 -25 -488
rect 25 488 71 500
rect 25 -488 31 488
rect 65 -488 71 488
rect 25 -500 71 -488
rect 121 488 167 500
rect 121 -488 127 488
rect 161 -488 167 488
rect 121 -500 167 -488
rect 217 488 263 500
rect 217 -488 223 488
rect 257 -488 263 488
rect 217 -500 263 -488
rect 313 488 359 500
rect 313 -488 319 488
rect 353 -488 359 488
rect 313 -500 359 -488
rect 409 488 455 500
rect 409 -488 415 488
rect 449 -488 455 488
rect 409 -500 455 -488
rect 505 488 551 500
rect 505 -488 511 488
rect 545 -488 551 488
rect 505 -500 551 -488
rect 601 488 647 500
rect 601 -488 607 488
rect 641 -488 647 488
rect 601 -500 647 -488
rect 697 488 743 500
rect 697 -488 703 488
rect 737 -488 743 488
rect 697 -500 743 -488
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string parameters w 5 l 0.150 m 1 nf 15 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
