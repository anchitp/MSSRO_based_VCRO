magic
tech sky130A
magscale 1 2
timestamp 1639056503
<< nwell >>
rect -23776 4274 29034 9480
rect -23774 3876 29034 4274
rect -23774 3582 16042 3876
rect -23774 3580 -230 3582
rect 14938 3580 16030 3582
rect -23774 3190 -4672 3580
<< pwell >>
rect 16604 3554 23726 3558
rect 16604 3314 29010 3554
rect -2244 2982 29010 3314
rect -23760 -2308 29010 2982
rect -2244 -2310 29010 -2308
rect -2244 -2312 15906 -2310
<< nmos >>
rect -23442 1854 -23412 2854
rect -23346 1854 -23316 2854
rect -23250 1854 -23220 2854
rect -23154 1854 -23124 2854
rect -23058 1854 -23028 2854
rect -22962 1854 -22932 2854
rect -22866 1854 -22836 2854
rect -22770 1854 -22740 2854
rect -22674 1854 -22644 2854
rect -22578 1854 -22548 2854
rect -22482 1854 -22452 2854
rect -22386 1854 -22356 2854
rect -22290 1854 -22260 2854
rect -22194 1854 -22164 2854
rect -22098 1854 -22068 2854
rect -22002 1854 -21972 2854
rect -21906 1854 -21876 2854
rect -21810 1854 -21780 2854
rect -21714 1854 -21684 2854
rect -21618 1854 -21588 2854
rect -21294 1846 -21264 2846
rect -21198 1846 -21168 2846
rect -21102 1846 -21072 2846
rect -21006 1846 -20976 2846
rect -20910 1846 -20880 2846
rect -20814 1846 -20784 2846
rect -20718 1846 -20688 2846
rect -20622 1846 -20592 2846
rect -20526 1846 -20496 2846
rect -20430 1846 -20400 2846
rect -20334 1846 -20304 2846
rect -20238 1846 -20208 2846
rect -20142 1846 -20112 2846
rect -20046 1846 -20016 2846
rect -19950 1846 -19920 2846
rect -19616 1850 -19586 2850
rect -19520 1850 -19490 2850
rect -19424 1850 -19394 2850
rect -19328 1850 -19298 2850
rect -19232 1850 -19202 2850
rect -19136 1850 -19106 2850
rect -19040 1850 -19010 2850
rect -18944 1850 -18914 2850
rect -18848 1850 -18818 2850
rect -18752 1850 -18722 2850
rect -18444 1860 -18414 2860
rect -18348 1860 -18318 2860
rect -18252 1860 -18222 2860
rect -18156 1860 -18126 2860
rect -18060 1860 -18030 2860
rect -16612 1866 -16582 2866
rect -16516 1866 -16486 2866
rect -16420 1866 -16390 2866
rect -16324 1866 -16294 2866
rect -16228 1866 -16198 2866
rect -16132 1866 -16102 2866
rect -16036 1866 -16006 2866
rect -15940 1866 -15910 2866
rect -15844 1866 -15814 2866
rect -15748 1866 -15718 2866
rect -15652 1866 -15622 2866
rect -15556 1866 -15526 2866
rect -15460 1866 -15430 2866
rect -15364 1866 -15334 2866
rect -15268 1866 -15238 2866
rect -15172 1866 -15142 2866
rect -15076 1866 -15046 2866
rect -14980 1866 -14950 2866
rect -14884 1866 -14854 2866
rect -14788 1866 -14758 2866
rect -14464 1858 -14434 2858
rect -14368 1858 -14338 2858
rect -14272 1858 -14242 2858
rect -14176 1858 -14146 2858
rect -14080 1858 -14050 2858
rect -13984 1858 -13954 2858
rect -13888 1858 -13858 2858
rect -13792 1858 -13762 2858
rect -13696 1858 -13666 2858
rect -13600 1858 -13570 2858
rect -13504 1858 -13474 2858
rect -13408 1858 -13378 2858
rect -13312 1858 -13282 2858
rect -13216 1858 -13186 2858
rect -13120 1858 -13090 2858
rect -12786 1862 -12756 2862
rect -12690 1862 -12660 2862
rect -12594 1862 -12564 2862
rect -12498 1862 -12468 2862
rect -12402 1862 -12372 2862
rect -12306 1862 -12276 2862
rect -12210 1862 -12180 2862
rect -12114 1862 -12084 2862
rect -12018 1862 -11988 2862
rect -11922 1862 -11892 2862
rect -11614 1872 -11584 2872
rect -11518 1872 -11488 2872
rect -11422 1872 -11392 2872
rect -11326 1872 -11296 2872
rect -11230 1872 -11200 2872
rect -10146 1864 -10116 2864
rect -10050 1864 -10020 2864
rect -9954 1864 -9924 2864
rect -9858 1864 -9828 2864
rect -9762 1864 -9732 2864
rect -9666 1864 -9636 2864
rect -9570 1864 -9540 2864
rect -9474 1864 -9444 2864
rect -9378 1864 -9348 2864
rect -9282 1864 -9252 2864
rect -9186 1864 -9156 2864
rect -9090 1864 -9060 2864
rect -8994 1864 -8964 2864
rect -8898 1864 -8868 2864
rect -8802 1864 -8772 2864
rect -8706 1864 -8676 2864
rect -8610 1864 -8580 2864
rect -8514 1864 -8484 2864
rect -8418 1864 -8388 2864
rect -8322 1864 -8292 2864
rect -7998 1856 -7968 2856
rect -7902 1856 -7872 2856
rect -7806 1856 -7776 2856
rect -7710 1856 -7680 2856
rect -7614 1856 -7584 2856
rect -7518 1856 -7488 2856
rect -7422 1856 -7392 2856
rect -7326 1856 -7296 2856
rect -7230 1856 -7200 2856
rect -7134 1856 -7104 2856
rect -7038 1856 -7008 2856
rect -6942 1856 -6912 2856
rect -6846 1856 -6816 2856
rect -6750 1856 -6720 2856
rect -6654 1856 -6624 2856
rect -6320 1860 -6290 2860
rect -6224 1860 -6194 2860
rect -6128 1860 -6098 2860
rect -6032 1860 -6002 2860
rect -5936 1860 -5906 2860
rect -5840 1860 -5810 2860
rect -5744 1860 -5714 2860
rect -5648 1860 -5618 2860
rect -5552 1860 -5522 2860
rect -5456 1860 -5426 2860
rect -5148 1870 -5118 2870
rect -5052 1870 -5022 2870
rect -4956 1870 -4926 2870
rect -4860 1870 -4830 2870
rect -4764 1870 -4734 2870
rect -1636 2236 -1606 3236
rect -1540 2236 -1510 3236
rect -1444 2236 -1414 3236
rect -1348 2236 -1318 3236
rect -1252 2236 -1222 3236
rect -1156 2236 -1126 3236
rect -1060 2236 -1030 3236
rect -964 2236 -934 3236
rect 1532 1830 1562 2830
rect 1628 1830 1658 2830
rect 1724 1830 1754 2830
rect 1820 1830 1850 2830
rect 2546 2076 2646 2276
rect 4488 1814 4518 2814
rect 4584 1814 4614 2814
rect 4680 1814 4710 2814
rect 4776 1814 4806 2814
rect 5546 2076 5646 2276
rect 7518 1814 7548 2814
rect 7614 1814 7644 2814
rect 7710 1814 7740 2814
rect 7806 1814 7836 2814
rect 8546 2076 8646 2276
rect 10606 1812 10636 2812
rect 10702 1812 10732 2812
rect 10798 1812 10828 2812
rect 10894 1812 10924 2812
rect 11546 2076 11646 2276
rect 13762 1786 13792 2786
rect 13858 1786 13888 2786
rect 13954 1786 13984 2786
rect 14050 1786 14080 2786
rect 16736 2534 16766 3534
rect 16832 2534 16862 3534
rect 16928 2534 16958 3534
rect 17024 2534 17054 3534
rect 17120 2534 17150 3534
rect 17428 2524 17458 3524
rect 17524 2524 17554 3524
rect 17620 2524 17650 3524
rect 17716 2524 17746 3524
rect 17812 2524 17842 3524
rect 17908 2524 17938 3524
rect 18004 2524 18034 3524
rect 18100 2524 18130 3524
rect 18196 2524 18226 3524
rect 18292 2524 18322 3524
rect 18626 2520 18656 3520
rect 18722 2520 18752 3520
rect 18818 2520 18848 3520
rect 18914 2520 18944 3520
rect 19010 2520 19040 3520
rect 19106 2520 19136 3520
rect 19202 2520 19232 3520
rect 19298 2520 19328 3520
rect 19394 2520 19424 3520
rect 19490 2520 19520 3520
rect 19586 2520 19616 3520
rect 19682 2520 19712 3520
rect 19778 2520 19808 3520
rect 19874 2520 19904 3520
rect 19970 2520 20000 3520
rect 20294 2528 20324 3528
rect 20390 2528 20420 3528
rect 20486 2528 20516 3528
rect 20582 2528 20612 3528
rect 20678 2528 20708 3528
rect 20774 2528 20804 3528
rect 20870 2528 20900 3528
rect 20966 2528 20996 3528
rect 21062 2528 21092 3528
rect 21158 2528 21188 3528
rect 21254 2528 21284 3528
rect 21350 2528 21380 3528
rect 21446 2528 21476 3528
rect 21542 2528 21572 3528
rect 21638 2528 21668 3528
rect 21734 2528 21764 3528
rect 21830 2528 21860 3528
rect 21926 2528 21956 3528
rect 22022 2528 22052 3528
rect 22118 2528 22148 3528
rect 23224 2532 23254 3532
rect 23320 2532 23350 3532
rect 23416 2532 23446 3532
rect 23512 2532 23542 3532
rect 23608 2532 23638 3532
rect 23916 2522 23946 3522
rect 24012 2522 24042 3522
rect 24108 2522 24138 3522
rect 24204 2522 24234 3522
rect 24300 2522 24330 3522
rect 24396 2522 24426 3522
rect 24492 2522 24522 3522
rect 24588 2522 24618 3522
rect 24684 2522 24714 3522
rect 24780 2522 24810 3522
rect 25114 2518 25144 3518
rect 25210 2518 25240 3518
rect 25306 2518 25336 3518
rect 25402 2518 25432 3518
rect 25498 2518 25528 3518
rect 25594 2518 25624 3518
rect 25690 2518 25720 3518
rect 25786 2518 25816 3518
rect 25882 2518 25912 3518
rect 25978 2518 26008 3518
rect 26074 2518 26104 3518
rect 26170 2518 26200 3518
rect 26266 2518 26296 3518
rect 26362 2518 26392 3518
rect 26458 2518 26488 3518
rect 26782 2526 26812 3526
rect 26878 2526 26908 3526
rect 26974 2526 27004 3526
rect 27070 2526 27100 3526
rect 27166 2526 27196 3526
rect 27262 2526 27292 3526
rect 27358 2526 27388 3526
rect 27454 2526 27484 3526
rect 27550 2526 27580 3526
rect 27646 2526 27676 3526
rect 27742 2526 27772 3526
rect 27838 2526 27868 3526
rect 27934 2526 27964 3526
rect 28030 2526 28060 3526
rect 28126 2526 28156 3526
rect 28222 2526 28252 3526
rect 28318 2526 28348 3526
rect 28414 2526 28444 3526
rect 28510 2526 28540 3526
rect 28606 2526 28636 3526
rect 14546 2076 14646 2276
rect -1640 66 -1600 1066
rect -1542 66 -1502 1066
rect -1444 66 -1404 1066
rect -1346 66 -1306 1066
rect -1248 66 -1208 1066
rect -1150 66 -1110 1066
rect -1052 66 -1012 1066
rect -954 66 -914 1066
rect 208 268 238 1268
rect 304 268 334 1268
rect 400 268 430 1268
rect 496 268 526 1268
rect 592 268 622 1268
rect 688 268 718 1268
rect 784 268 814 1268
rect 880 268 910 1268
rect 976 268 1006 1268
rect 1072 268 1102 1268
rect 1168 268 1198 1268
rect 1264 268 1294 1268
rect 1976 268 2006 1268
rect 2072 268 2102 1268
rect 2168 268 2198 1268
rect 2264 268 2294 1268
rect 2360 268 2390 1268
rect 2456 268 2486 1268
rect 2552 268 2582 1268
rect 2648 268 2678 1268
rect 2744 268 2774 1268
rect 2840 268 2870 1268
rect 2936 268 2966 1268
rect 3164 252 3194 1252
rect 3260 252 3290 1252
rect 3356 252 3386 1252
rect 3452 252 3482 1252
rect 3548 252 3578 1252
rect 3644 252 3674 1252
rect 3740 252 3770 1252
rect 3836 252 3866 1252
rect 3932 252 3962 1252
rect 4028 252 4058 1252
rect 4124 252 4154 1252
rect 4220 252 4250 1252
rect 4932 252 4962 1252
rect 5028 252 5058 1252
rect 5124 252 5154 1252
rect 5220 252 5250 1252
rect 5316 252 5346 1252
rect 5412 252 5442 1252
rect 5508 252 5538 1252
rect 5604 252 5634 1252
rect 5700 252 5730 1252
rect 5796 252 5826 1252
rect 5892 252 5922 1252
rect 6194 252 6224 1252
rect 6290 252 6320 1252
rect 6386 252 6416 1252
rect 6482 252 6512 1252
rect 6578 252 6608 1252
rect 6674 252 6704 1252
rect 6770 252 6800 1252
rect 6866 252 6896 1252
rect 6962 252 6992 1252
rect 7058 252 7088 1252
rect 7154 252 7184 1252
rect 7250 252 7280 1252
rect 7962 252 7992 1252
rect 8058 252 8088 1252
rect 8154 252 8184 1252
rect 8250 252 8280 1252
rect 8346 252 8376 1252
rect 8442 252 8472 1252
rect 8538 252 8568 1252
rect 8634 252 8664 1252
rect 8730 252 8760 1252
rect 8826 252 8856 1252
rect 8922 252 8952 1252
rect 9282 250 9312 1250
rect 9378 250 9408 1250
rect 9474 250 9504 1250
rect 9570 250 9600 1250
rect 9666 250 9696 1250
rect 9762 250 9792 1250
rect 9858 250 9888 1250
rect 9954 250 9984 1250
rect 10050 250 10080 1250
rect 10146 250 10176 1250
rect 10242 250 10272 1250
rect 10338 250 10368 1250
rect 11050 250 11080 1250
rect 11146 250 11176 1250
rect 11242 250 11272 1250
rect 11338 250 11368 1250
rect 11434 250 11464 1250
rect 11530 250 11560 1250
rect 11626 250 11656 1250
rect 11722 250 11752 1250
rect 11818 250 11848 1250
rect 11914 250 11944 1250
rect 12010 250 12040 1250
rect 12438 224 12468 1224
rect 12534 224 12564 1224
rect 12630 224 12660 1224
rect 12726 224 12756 1224
rect 12822 224 12852 1224
rect 12918 224 12948 1224
rect 13014 224 13044 1224
rect 13110 224 13140 1224
rect 13206 224 13236 1224
rect 13302 224 13332 1224
rect 13398 224 13428 1224
rect 13494 224 13524 1224
rect 14206 224 14236 1224
rect 14302 224 14332 1224
rect 14398 224 14428 1224
rect 14494 224 14524 1224
rect 14590 224 14620 1224
rect 14686 224 14716 1224
rect 14782 224 14812 1224
rect 14878 224 14908 1224
rect 14974 224 15004 1224
rect 15070 224 15100 1224
rect 15166 224 15196 1224
rect 15468 100 15498 1300
<< pmos >>
rect -1606 4936 -1566 5936
rect -1508 4936 -1468 5936
rect -1410 4936 -1370 5936
rect -1312 4936 -1272 5936
rect -1214 4936 -1174 5936
rect -1116 4936 -1076 5936
rect -1018 4936 -978 5936
rect -920 4936 -880 5936
rect 244 5606 274 6606
rect 340 5606 370 6606
rect 436 5606 466 6606
rect 532 5606 562 6606
rect 628 5606 658 6606
rect 724 5606 754 6606
rect 820 5606 850 6606
rect 916 5606 946 6606
rect 1012 5606 1042 6606
rect 1108 5606 1138 6606
rect 1204 5606 1234 6606
rect 1300 5606 1330 6606
rect 2010 5602 2040 6602
rect 2106 5602 2136 6602
rect 2202 5602 2232 6602
rect 2298 5602 2328 6602
rect 2394 5602 2424 6602
rect 2490 5602 2520 6602
rect 2586 5602 2616 6602
rect 2682 5602 2712 6602
rect 3200 5590 3230 6590
rect 3296 5590 3326 6590
rect 3392 5590 3422 6590
rect 3488 5590 3518 6590
rect 3584 5590 3614 6590
rect 3680 5590 3710 6590
rect 3776 5590 3806 6590
rect 3872 5590 3902 6590
rect 3968 5590 3998 6590
rect 4064 5590 4094 6590
rect 4160 5590 4190 6590
rect 4256 5590 4286 6590
rect 4966 5586 4996 6586
rect 5062 5586 5092 6586
rect 5158 5586 5188 6586
rect 5254 5586 5284 6586
rect 5350 5586 5380 6586
rect 5446 5586 5476 6586
rect 5542 5586 5572 6586
rect 5638 5586 5668 6586
rect 6230 5590 6260 6590
rect 6326 5590 6356 6590
rect 6422 5590 6452 6590
rect 6518 5590 6548 6590
rect 6614 5590 6644 6590
rect 6710 5590 6740 6590
rect 6806 5590 6836 6590
rect 6902 5590 6932 6590
rect 6998 5590 7028 6590
rect 7094 5590 7124 6590
rect 7190 5590 7220 6590
rect 7286 5590 7316 6590
rect 7996 5586 8026 6586
rect 8092 5586 8122 6586
rect 8188 5586 8218 6586
rect 8284 5586 8314 6586
rect 8380 5586 8410 6586
rect 8476 5586 8506 6586
rect 8572 5586 8602 6586
rect 8668 5586 8698 6586
rect 9318 5588 9348 6588
rect 9414 5588 9444 6588
rect 9510 5588 9540 6588
rect 9606 5588 9636 6588
rect 9702 5588 9732 6588
rect 9798 5588 9828 6588
rect 9894 5588 9924 6588
rect 9990 5588 10020 6588
rect 10086 5588 10116 6588
rect 10182 5588 10212 6588
rect 10278 5588 10308 6588
rect 10374 5588 10404 6588
rect 11084 5584 11114 6584
rect 11180 5584 11210 6584
rect 11276 5584 11306 6584
rect 11372 5584 11402 6584
rect 11468 5584 11498 6584
rect 11564 5584 11594 6584
rect 11660 5584 11690 6584
rect 11756 5584 11786 6584
rect 12474 5562 12504 6562
rect 12570 5562 12600 6562
rect 12666 5562 12696 6562
rect 12762 5562 12792 6562
rect 12858 5562 12888 6562
rect 12954 5562 12984 6562
rect 13050 5562 13080 6562
rect 13146 5562 13176 6562
rect 13242 5562 13272 6562
rect 13338 5562 13368 6562
rect 13434 5562 13464 6562
rect 13530 5562 13560 6562
rect 14240 5558 14270 6558
rect 14336 5558 14366 6558
rect 14432 5558 14462 6558
rect 14528 5558 14558 6558
rect 14624 5558 14654 6558
rect 14720 5558 14750 6558
rect 14816 5558 14846 6558
rect 14912 5558 14942 6558
rect -23536 3442 -23506 4442
rect -23440 3442 -23410 4442
rect -23344 3442 -23314 4442
rect -23248 3442 -23218 4442
rect -23152 3442 -23122 4442
rect -23056 3442 -23026 4442
rect -22960 3442 -22930 4442
rect -22864 3442 -22834 4442
rect -22768 3442 -22738 4442
rect -22672 3442 -22642 4442
rect -22576 3442 -22546 4442
rect -22480 3442 -22450 4442
rect -22384 3442 -22354 4442
rect -22288 3442 -22258 4442
rect -22192 3442 -22162 4442
rect -22096 3442 -22066 4442
rect -22000 3442 -21970 4442
rect -21904 3442 -21874 4442
rect -21808 3442 -21778 4442
rect -21712 3442 -21682 4442
rect -21392 3448 -21362 4448
rect -21296 3448 -21266 4448
rect -21200 3448 -21170 4448
rect -21104 3448 -21074 4448
rect -21008 3448 -20978 4448
rect -20912 3448 -20882 4448
rect -20816 3448 -20786 4448
rect -20720 3448 -20690 4448
rect -20624 3448 -20594 4448
rect -20528 3448 -20498 4448
rect -20432 3448 -20402 4448
rect -20336 3448 -20306 4448
rect -20240 3448 -20210 4448
rect -20144 3448 -20114 4448
rect -20048 3448 -20018 4448
rect -19708 3454 -19678 4454
rect -19612 3454 -19582 4454
rect -19516 3454 -19486 4454
rect -19420 3454 -19390 4454
rect -19324 3454 -19294 4454
rect -19228 3454 -19198 4454
rect -19132 3454 -19102 4454
rect -19036 3454 -19006 4454
rect -18940 3454 -18910 4454
rect -18844 3454 -18814 4454
rect -18540 3456 -18510 4456
rect -18444 3456 -18414 4456
rect -18348 3456 -18318 4456
rect -18252 3456 -18222 4456
rect -18156 3456 -18126 4456
rect -16706 3454 -16676 4454
rect -16610 3454 -16580 4454
rect -16514 3454 -16484 4454
rect -16418 3454 -16388 4454
rect -16322 3454 -16292 4454
rect -16226 3454 -16196 4454
rect -16130 3454 -16100 4454
rect -16034 3454 -16004 4454
rect -15938 3454 -15908 4454
rect -15842 3454 -15812 4454
rect -15746 3454 -15716 4454
rect -15650 3454 -15620 4454
rect -15554 3454 -15524 4454
rect -15458 3454 -15428 4454
rect -15362 3454 -15332 4454
rect -15266 3454 -15236 4454
rect -15170 3454 -15140 4454
rect -15074 3454 -15044 4454
rect -14978 3454 -14948 4454
rect -14882 3454 -14852 4454
rect -14562 3460 -14532 4460
rect -14466 3460 -14436 4460
rect -14370 3460 -14340 4460
rect -14274 3460 -14244 4460
rect -14178 3460 -14148 4460
rect -14082 3460 -14052 4460
rect -13986 3460 -13956 4460
rect -13890 3460 -13860 4460
rect -13794 3460 -13764 4460
rect -13698 3460 -13668 4460
rect -13602 3460 -13572 4460
rect -13506 3460 -13476 4460
rect -13410 3460 -13380 4460
rect -13314 3460 -13284 4460
rect -13218 3460 -13188 4460
rect -12878 3466 -12848 4466
rect -12782 3466 -12752 4466
rect -12686 3466 -12656 4466
rect -12590 3466 -12560 4466
rect -12494 3466 -12464 4466
rect -12398 3466 -12368 4466
rect -12302 3466 -12272 4466
rect -12206 3466 -12176 4466
rect -12110 3466 -12080 4466
rect -12014 3466 -11984 4466
rect -11710 3468 -11680 4468
rect -11614 3468 -11584 4468
rect -11518 3468 -11488 4468
rect -11422 3468 -11392 4468
rect -11326 3468 -11296 4468
rect -10240 3452 -10210 4452
rect -10144 3452 -10114 4452
rect -10048 3452 -10018 4452
rect -9952 3452 -9922 4452
rect -9856 3452 -9826 4452
rect -9760 3452 -9730 4452
rect -9664 3452 -9634 4452
rect -9568 3452 -9538 4452
rect -9472 3452 -9442 4452
rect -9376 3452 -9346 4452
rect -9280 3452 -9250 4452
rect -9184 3452 -9154 4452
rect -9088 3452 -9058 4452
rect -8992 3452 -8962 4452
rect -8896 3452 -8866 4452
rect -8800 3452 -8770 4452
rect -8704 3452 -8674 4452
rect -8608 3452 -8578 4452
rect -8512 3452 -8482 4452
rect -8416 3452 -8386 4452
rect -8096 3458 -8066 4458
rect -8000 3458 -7970 4458
rect -7904 3458 -7874 4458
rect -7808 3458 -7778 4458
rect -7712 3458 -7682 4458
rect -7616 3458 -7586 4458
rect -7520 3458 -7490 4458
rect -7424 3458 -7394 4458
rect -7328 3458 -7298 4458
rect -7232 3458 -7202 4458
rect -7136 3458 -7106 4458
rect -7040 3458 -7010 4458
rect -6944 3458 -6914 4458
rect -6848 3458 -6818 4458
rect -6752 3458 -6722 4458
rect -6412 3464 -6382 4464
rect -6316 3464 -6286 4464
rect -6220 3464 -6190 4464
rect -6124 3464 -6094 4464
rect -6028 3464 -5998 4464
rect -5932 3464 -5902 4464
rect -5836 3464 -5806 4464
rect -5740 3464 -5710 4464
rect -5644 3464 -5614 4464
rect -5548 3464 -5518 4464
rect -5244 3466 -5214 4466
rect -5148 3466 -5118 4466
rect -5052 3466 -5022 4466
rect -4956 3466 -4926 4466
rect -4860 3466 -4830 4466
rect 1534 3944 1564 4944
rect 1630 3944 1660 4944
rect 1726 3944 1756 4944
rect 1822 3944 1852 4944
rect 4490 3928 4520 4928
rect 4586 3928 4616 4928
rect 4682 3928 4712 4928
rect 4778 3928 4808 4928
rect 7520 3928 7550 4928
rect 7616 3928 7646 4928
rect 7712 3928 7742 4928
rect 7808 3928 7838 4928
rect 10608 3926 10638 4926
rect 10704 3926 10734 4926
rect 10800 3926 10830 4926
rect 10896 3926 10926 4926
rect 13764 3900 13794 4900
rect 13860 3900 13890 4900
rect 13956 3900 13986 4900
rect 14052 3900 14082 4900
rect 15568 3926 15598 5926
rect 15664 3926 15694 5926
rect 16832 4130 16862 5130
rect 16928 4130 16958 5130
rect 17024 4130 17054 5130
rect 17120 4130 17150 5130
rect 17216 4130 17246 5130
rect 17520 4128 17550 5128
rect 17616 4128 17646 5128
rect 17712 4128 17742 5128
rect 17808 4128 17838 5128
rect 17904 4128 17934 5128
rect 18000 4128 18030 5128
rect 18096 4128 18126 5128
rect 18192 4128 18222 5128
rect 18288 4128 18318 5128
rect 18384 4128 18414 5128
rect 18724 4122 18754 5122
rect 18820 4122 18850 5122
rect 18916 4122 18946 5122
rect 19012 4122 19042 5122
rect 19108 4122 19138 5122
rect 19204 4122 19234 5122
rect 19300 4122 19330 5122
rect 19396 4122 19426 5122
rect 19492 4122 19522 5122
rect 19588 4122 19618 5122
rect 19684 4122 19714 5122
rect 19780 4122 19810 5122
rect 19876 4122 19906 5122
rect 19972 4122 20002 5122
rect 20068 4122 20098 5122
rect 20388 4116 20418 5116
rect 20484 4116 20514 5116
rect 20580 4116 20610 5116
rect 20676 4116 20706 5116
rect 20772 4116 20802 5116
rect 20868 4116 20898 5116
rect 20964 4116 20994 5116
rect 21060 4116 21090 5116
rect 21156 4116 21186 5116
rect 21252 4116 21282 5116
rect 21348 4116 21378 5116
rect 21444 4116 21474 5116
rect 21540 4116 21570 5116
rect 21636 4116 21666 5116
rect 21732 4116 21762 5116
rect 21828 4116 21858 5116
rect 21924 4116 21954 5116
rect 22020 4116 22050 5116
rect 22116 4116 22146 5116
rect 22212 4116 22242 5116
rect 23320 4128 23350 5128
rect 23416 4128 23446 5128
rect 23512 4128 23542 5128
rect 23608 4128 23638 5128
rect 23704 4128 23734 5128
rect 24008 4126 24038 5126
rect 24104 4126 24134 5126
rect 24200 4126 24230 5126
rect 24296 4126 24326 5126
rect 24392 4126 24422 5126
rect 24488 4126 24518 5126
rect 24584 4126 24614 5126
rect 24680 4126 24710 5126
rect 24776 4126 24806 5126
rect 24872 4126 24902 5126
rect 25212 4120 25242 5120
rect 25308 4120 25338 5120
rect 25404 4120 25434 5120
rect 25500 4120 25530 5120
rect 25596 4120 25626 5120
rect 25692 4120 25722 5120
rect 25788 4120 25818 5120
rect 25884 4120 25914 5120
rect 25980 4120 26010 5120
rect 26076 4120 26106 5120
rect 26172 4120 26202 5120
rect 26268 4120 26298 5120
rect 26364 4120 26394 5120
rect 26460 4120 26490 5120
rect 26556 4120 26586 5120
rect 26876 4114 26906 5114
rect 26972 4114 27002 5114
rect 27068 4114 27098 5114
rect 27164 4114 27194 5114
rect 27260 4114 27290 5114
rect 27356 4114 27386 5114
rect 27452 4114 27482 5114
rect 27548 4114 27578 5114
rect 27644 4114 27674 5114
rect 27740 4114 27770 5114
rect 27836 4114 27866 5114
rect 27932 4114 27962 5114
rect 28028 4114 28058 5114
rect 28124 4114 28154 5114
rect 28220 4114 28250 5114
rect 28316 4114 28346 5114
rect 28412 4114 28442 5114
rect 28508 4114 28538 5114
rect 28604 4114 28634 5114
rect 28700 4114 28730 5114
<< ndiff >>
rect 16674 3493 16736 3534
rect 16674 3459 16686 3493
rect 16720 3459 16736 3493
rect 16674 3425 16736 3459
rect 16674 3391 16686 3425
rect 16720 3391 16736 3425
rect 16674 3357 16736 3391
rect 16674 3323 16686 3357
rect 16720 3323 16736 3357
rect 16674 3289 16736 3323
rect 16674 3255 16686 3289
rect 16720 3255 16736 3289
rect -1698 3195 -1636 3236
rect -1698 3161 -1686 3195
rect -1652 3161 -1636 3195
rect -1698 3127 -1636 3161
rect -1698 3093 -1686 3127
rect -1652 3093 -1636 3127
rect -23504 2813 -23442 2854
rect -23504 2779 -23492 2813
rect -23458 2779 -23442 2813
rect -23504 2745 -23442 2779
rect -23504 2711 -23492 2745
rect -23458 2711 -23442 2745
rect -23504 2677 -23442 2711
rect -23504 2643 -23492 2677
rect -23458 2643 -23442 2677
rect -23504 2609 -23442 2643
rect -23504 2575 -23492 2609
rect -23458 2575 -23442 2609
rect -23504 2541 -23442 2575
rect -23504 2507 -23492 2541
rect -23458 2507 -23442 2541
rect -23504 2473 -23442 2507
rect -23504 2439 -23492 2473
rect -23458 2439 -23442 2473
rect -23504 2405 -23442 2439
rect -23504 2371 -23492 2405
rect -23458 2371 -23442 2405
rect -23504 2337 -23442 2371
rect -23504 2303 -23492 2337
rect -23458 2303 -23442 2337
rect -23504 2269 -23442 2303
rect -23504 2235 -23492 2269
rect -23458 2235 -23442 2269
rect -23504 2201 -23442 2235
rect -23504 2167 -23492 2201
rect -23458 2167 -23442 2201
rect -23504 2133 -23442 2167
rect -23504 2099 -23492 2133
rect -23458 2099 -23442 2133
rect -23504 2065 -23442 2099
rect -23504 2031 -23492 2065
rect -23458 2031 -23442 2065
rect -23504 1997 -23442 2031
rect -23504 1963 -23492 1997
rect -23458 1963 -23442 1997
rect -23504 1929 -23442 1963
rect -23504 1895 -23492 1929
rect -23458 1895 -23442 1929
rect -23504 1854 -23442 1895
rect -23412 2813 -23346 2854
rect -23412 2779 -23396 2813
rect -23362 2779 -23346 2813
rect -23412 2745 -23346 2779
rect -23412 2711 -23396 2745
rect -23362 2711 -23346 2745
rect -23412 2677 -23346 2711
rect -23412 2643 -23396 2677
rect -23362 2643 -23346 2677
rect -23412 2609 -23346 2643
rect -23412 2575 -23396 2609
rect -23362 2575 -23346 2609
rect -23412 2541 -23346 2575
rect -23412 2507 -23396 2541
rect -23362 2507 -23346 2541
rect -23412 2473 -23346 2507
rect -23412 2439 -23396 2473
rect -23362 2439 -23346 2473
rect -23412 2405 -23346 2439
rect -23412 2371 -23396 2405
rect -23362 2371 -23346 2405
rect -23412 2337 -23346 2371
rect -23412 2303 -23396 2337
rect -23362 2303 -23346 2337
rect -23412 2269 -23346 2303
rect -23412 2235 -23396 2269
rect -23362 2235 -23346 2269
rect -23412 2201 -23346 2235
rect -23412 2167 -23396 2201
rect -23362 2167 -23346 2201
rect -23412 2133 -23346 2167
rect -23412 2099 -23396 2133
rect -23362 2099 -23346 2133
rect -23412 2065 -23346 2099
rect -23412 2031 -23396 2065
rect -23362 2031 -23346 2065
rect -23412 1997 -23346 2031
rect -23412 1963 -23396 1997
rect -23362 1963 -23346 1997
rect -23412 1929 -23346 1963
rect -23412 1895 -23396 1929
rect -23362 1895 -23346 1929
rect -23412 1854 -23346 1895
rect -23316 2813 -23250 2854
rect -23316 2779 -23300 2813
rect -23266 2779 -23250 2813
rect -23316 2745 -23250 2779
rect -23316 2711 -23300 2745
rect -23266 2711 -23250 2745
rect -23316 2677 -23250 2711
rect -23316 2643 -23300 2677
rect -23266 2643 -23250 2677
rect -23316 2609 -23250 2643
rect -23316 2575 -23300 2609
rect -23266 2575 -23250 2609
rect -23316 2541 -23250 2575
rect -23316 2507 -23300 2541
rect -23266 2507 -23250 2541
rect -23316 2473 -23250 2507
rect -23316 2439 -23300 2473
rect -23266 2439 -23250 2473
rect -23316 2405 -23250 2439
rect -23316 2371 -23300 2405
rect -23266 2371 -23250 2405
rect -23316 2337 -23250 2371
rect -23316 2303 -23300 2337
rect -23266 2303 -23250 2337
rect -23316 2269 -23250 2303
rect -23316 2235 -23300 2269
rect -23266 2235 -23250 2269
rect -23316 2201 -23250 2235
rect -23316 2167 -23300 2201
rect -23266 2167 -23250 2201
rect -23316 2133 -23250 2167
rect -23316 2099 -23300 2133
rect -23266 2099 -23250 2133
rect -23316 2065 -23250 2099
rect -23316 2031 -23300 2065
rect -23266 2031 -23250 2065
rect -23316 1997 -23250 2031
rect -23316 1963 -23300 1997
rect -23266 1963 -23250 1997
rect -23316 1929 -23250 1963
rect -23316 1895 -23300 1929
rect -23266 1895 -23250 1929
rect -23316 1854 -23250 1895
rect -23220 2813 -23154 2854
rect -23220 2779 -23204 2813
rect -23170 2779 -23154 2813
rect -23220 2745 -23154 2779
rect -23220 2711 -23204 2745
rect -23170 2711 -23154 2745
rect -23220 2677 -23154 2711
rect -23220 2643 -23204 2677
rect -23170 2643 -23154 2677
rect -23220 2609 -23154 2643
rect -23220 2575 -23204 2609
rect -23170 2575 -23154 2609
rect -23220 2541 -23154 2575
rect -23220 2507 -23204 2541
rect -23170 2507 -23154 2541
rect -23220 2473 -23154 2507
rect -23220 2439 -23204 2473
rect -23170 2439 -23154 2473
rect -23220 2405 -23154 2439
rect -23220 2371 -23204 2405
rect -23170 2371 -23154 2405
rect -23220 2337 -23154 2371
rect -23220 2303 -23204 2337
rect -23170 2303 -23154 2337
rect -23220 2269 -23154 2303
rect -23220 2235 -23204 2269
rect -23170 2235 -23154 2269
rect -23220 2201 -23154 2235
rect -23220 2167 -23204 2201
rect -23170 2167 -23154 2201
rect -23220 2133 -23154 2167
rect -23220 2099 -23204 2133
rect -23170 2099 -23154 2133
rect -23220 2065 -23154 2099
rect -23220 2031 -23204 2065
rect -23170 2031 -23154 2065
rect -23220 1997 -23154 2031
rect -23220 1963 -23204 1997
rect -23170 1963 -23154 1997
rect -23220 1929 -23154 1963
rect -23220 1895 -23204 1929
rect -23170 1895 -23154 1929
rect -23220 1854 -23154 1895
rect -23124 2813 -23058 2854
rect -23124 2779 -23108 2813
rect -23074 2779 -23058 2813
rect -23124 2745 -23058 2779
rect -23124 2711 -23108 2745
rect -23074 2711 -23058 2745
rect -23124 2677 -23058 2711
rect -23124 2643 -23108 2677
rect -23074 2643 -23058 2677
rect -23124 2609 -23058 2643
rect -23124 2575 -23108 2609
rect -23074 2575 -23058 2609
rect -23124 2541 -23058 2575
rect -23124 2507 -23108 2541
rect -23074 2507 -23058 2541
rect -23124 2473 -23058 2507
rect -23124 2439 -23108 2473
rect -23074 2439 -23058 2473
rect -23124 2405 -23058 2439
rect -23124 2371 -23108 2405
rect -23074 2371 -23058 2405
rect -23124 2337 -23058 2371
rect -23124 2303 -23108 2337
rect -23074 2303 -23058 2337
rect -23124 2269 -23058 2303
rect -23124 2235 -23108 2269
rect -23074 2235 -23058 2269
rect -23124 2201 -23058 2235
rect -23124 2167 -23108 2201
rect -23074 2167 -23058 2201
rect -23124 2133 -23058 2167
rect -23124 2099 -23108 2133
rect -23074 2099 -23058 2133
rect -23124 2065 -23058 2099
rect -23124 2031 -23108 2065
rect -23074 2031 -23058 2065
rect -23124 1997 -23058 2031
rect -23124 1963 -23108 1997
rect -23074 1963 -23058 1997
rect -23124 1929 -23058 1963
rect -23124 1895 -23108 1929
rect -23074 1895 -23058 1929
rect -23124 1854 -23058 1895
rect -23028 2813 -22962 2854
rect -23028 2779 -23012 2813
rect -22978 2779 -22962 2813
rect -23028 2745 -22962 2779
rect -23028 2711 -23012 2745
rect -22978 2711 -22962 2745
rect -23028 2677 -22962 2711
rect -23028 2643 -23012 2677
rect -22978 2643 -22962 2677
rect -23028 2609 -22962 2643
rect -23028 2575 -23012 2609
rect -22978 2575 -22962 2609
rect -23028 2541 -22962 2575
rect -23028 2507 -23012 2541
rect -22978 2507 -22962 2541
rect -23028 2473 -22962 2507
rect -23028 2439 -23012 2473
rect -22978 2439 -22962 2473
rect -23028 2405 -22962 2439
rect -23028 2371 -23012 2405
rect -22978 2371 -22962 2405
rect -23028 2337 -22962 2371
rect -23028 2303 -23012 2337
rect -22978 2303 -22962 2337
rect -23028 2269 -22962 2303
rect -23028 2235 -23012 2269
rect -22978 2235 -22962 2269
rect -23028 2201 -22962 2235
rect -23028 2167 -23012 2201
rect -22978 2167 -22962 2201
rect -23028 2133 -22962 2167
rect -23028 2099 -23012 2133
rect -22978 2099 -22962 2133
rect -23028 2065 -22962 2099
rect -23028 2031 -23012 2065
rect -22978 2031 -22962 2065
rect -23028 1997 -22962 2031
rect -23028 1963 -23012 1997
rect -22978 1963 -22962 1997
rect -23028 1929 -22962 1963
rect -23028 1895 -23012 1929
rect -22978 1895 -22962 1929
rect -23028 1854 -22962 1895
rect -22932 2813 -22866 2854
rect -22932 2779 -22916 2813
rect -22882 2779 -22866 2813
rect -22932 2745 -22866 2779
rect -22932 2711 -22916 2745
rect -22882 2711 -22866 2745
rect -22932 2677 -22866 2711
rect -22932 2643 -22916 2677
rect -22882 2643 -22866 2677
rect -22932 2609 -22866 2643
rect -22932 2575 -22916 2609
rect -22882 2575 -22866 2609
rect -22932 2541 -22866 2575
rect -22932 2507 -22916 2541
rect -22882 2507 -22866 2541
rect -22932 2473 -22866 2507
rect -22932 2439 -22916 2473
rect -22882 2439 -22866 2473
rect -22932 2405 -22866 2439
rect -22932 2371 -22916 2405
rect -22882 2371 -22866 2405
rect -22932 2337 -22866 2371
rect -22932 2303 -22916 2337
rect -22882 2303 -22866 2337
rect -22932 2269 -22866 2303
rect -22932 2235 -22916 2269
rect -22882 2235 -22866 2269
rect -22932 2201 -22866 2235
rect -22932 2167 -22916 2201
rect -22882 2167 -22866 2201
rect -22932 2133 -22866 2167
rect -22932 2099 -22916 2133
rect -22882 2099 -22866 2133
rect -22932 2065 -22866 2099
rect -22932 2031 -22916 2065
rect -22882 2031 -22866 2065
rect -22932 1997 -22866 2031
rect -22932 1963 -22916 1997
rect -22882 1963 -22866 1997
rect -22932 1929 -22866 1963
rect -22932 1895 -22916 1929
rect -22882 1895 -22866 1929
rect -22932 1854 -22866 1895
rect -22836 2813 -22770 2854
rect -22836 2779 -22820 2813
rect -22786 2779 -22770 2813
rect -22836 2745 -22770 2779
rect -22836 2711 -22820 2745
rect -22786 2711 -22770 2745
rect -22836 2677 -22770 2711
rect -22836 2643 -22820 2677
rect -22786 2643 -22770 2677
rect -22836 2609 -22770 2643
rect -22836 2575 -22820 2609
rect -22786 2575 -22770 2609
rect -22836 2541 -22770 2575
rect -22836 2507 -22820 2541
rect -22786 2507 -22770 2541
rect -22836 2473 -22770 2507
rect -22836 2439 -22820 2473
rect -22786 2439 -22770 2473
rect -22836 2405 -22770 2439
rect -22836 2371 -22820 2405
rect -22786 2371 -22770 2405
rect -22836 2337 -22770 2371
rect -22836 2303 -22820 2337
rect -22786 2303 -22770 2337
rect -22836 2269 -22770 2303
rect -22836 2235 -22820 2269
rect -22786 2235 -22770 2269
rect -22836 2201 -22770 2235
rect -22836 2167 -22820 2201
rect -22786 2167 -22770 2201
rect -22836 2133 -22770 2167
rect -22836 2099 -22820 2133
rect -22786 2099 -22770 2133
rect -22836 2065 -22770 2099
rect -22836 2031 -22820 2065
rect -22786 2031 -22770 2065
rect -22836 1997 -22770 2031
rect -22836 1963 -22820 1997
rect -22786 1963 -22770 1997
rect -22836 1929 -22770 1963
rect -22836 1895 -22820 1929
rect -22786 1895 -22770 1929
rect -22836 1854 -22770 1895
rect -22740 2813 -22674 2854
rect -22740 2779 -22724 2813
rect -22690 2779 -22674 2813
rect -22740 2745 -22674 2779
rect -22740 2711 -22724 2745
rect -22690 2711 -22674 2745
rect -22740 2677 -22674 2711
rect -22740 2643 -22724 2677
rect -22690 2643 -22674 2677
rect -22740 2609 -22674 2643
rect -22740 2575 -22724 2609
rect -22690 2575 -22674 2609
rect -22740 2541 -22674 2575
rect -22740 2507 -22724 2541
rect -22690 2507 -22674 2541
rect -22740 2473 -22674 2507
rect -22740 2439 -22724 2473
rect -22690 2439 -22674 2473
rect -22740 2405 -22674 2439
rect -22740 2371 -22724 2405
rect -22690 2371 -22674 2405
rect -22740 2337 -22674 2371
rect -22740 2303 -22724 2337
rect -22690 2303 -22674 2337
rect -22740 2269 -22674 2303
rect -22740 2235 -22724 2269
rect -22690 2235 -22674 2269
rect -22740 2201 -22674 2235
rect -22740 2167 -22724 2201
rect -22690 2167 -22674 2201
rect -22740 2133 -22674 2167
rect -22740 2099 -22724 2133
rect -22690 2099 -22674 2133
rect -22740 2065 -22674 2099
rect -22740 2031 -22724 2065
rect -22690 2031 -22674 2065
rect -22740 1997 -22674 2031
rect -22740 1963 -22724 1997
rect -22690 1963 -22674 1997
rect -22740 1929 -22674 1963
rect -22740 1895 -22724 1929
rect -22690 1895 -22674 1929
rect -22740 1854 -22674 1895
rect -22644 2813 -22578 2854
rect -22644 2779 -22628 2813
rect -22594 2779 -22578 2813
rect -22644 2745 -22578 2779
rect -22644 2711 -22628 2745
rect -22594 2711 -22578 2745
rect -22644 2677 -22578 2711
rect -22644 2643 -22628 2677
rect -22594 2643 -22578 2677
rect -22644 2609 -22578 2643
rect -22644 2575 -22628 2609
rect -22594 2575 -22578 2609
rect -22644 2541 -22578 2575
rect -22644 2507 -22628 2541
rect -22594 2507 -22578 2541
rect -22644 2473 -22578 2507
rect -22644 2439 -22628 2473
rect -22594 2439 -22578 2473
rect -22644 2405 -22578 2439
rect -22644 2371 -22628 2405
rect -22594 2371 -22578 2405
rect -22644 2337 -22578 2371
rect -22644 2303 -22628 2337
rect -22594 2303 -22578 2337
rect -22644 2269 -22578 2303
rect -22644 2235 -22628 2269
rect -22594 2235 -22578 2269
rect -22644 2201 -22578 2235
rect -22644 2167 -22628 2201
rect -22594 2167 -22578 2201
rect -22644 2133 -22578 2167
rect -22644 2099 -22628 2133
rect -22594 2099 -22578 2133
rect -22644 2065 -22578 2099
rect -22644 2031 -22628 2065
rect -22594 2031 -22578 2065
rect -22644 1997 -22578 2031
rect -22644 1963 -22628 1997
rect -22594 1963 -22578 1997
rect -22644 1929 -22578 1963
rect -22644 1895 -22628 1929
rect -22594 1895 -22578 1929
rect -22644 1854 -22578 1895
rect -22548 2813 -22482 2854
rect -22548 2779 -22532 2813
rect -22498 2779 -22482 2813
rect -22548 2745 -22482 2779
rect -22548 2711 -22532 2745
rect -22498 2711 -22482 2745
rect -22548 2677 -22482 2711
rect -22548 2643 -22532 2677
rect -22498 2643 -22482 2677
rect -22548 2609 -22482 2643
rect -22548 2575 -22532 2609
rect -22498 2575 -22482 2609
rect -22548 2541 -22482 2575
rect -22548 2507 -22532 2541
rect -22498 2507 -22482 2541
rect -22548 2473 -22482 2507
rect -22548 2439 -22532 2473
rect -22498 2439 -22482 2473
rect -22548 2405 -22482 2439
rect -22548 2371 -22532 2405
rect -22498 2371 -22482 2405
rect -22548 2337 -22482 2371
rect -22548 2303 -22532 2337
rect -22498 2303 -22482 2337
rect -22548 2269 -22482 2303
rect -22548 2235 -22532 2269
rect -22498 2235 -22482 2269
rect -22548 2201 -22482 2235
rect -22548 2167 -22532 2201
rect -22498 2167 -22482 2201
rect -22548 2133 -22482 2167
rect -22548 2099 -22532 2133
rect -22498 2099 -22482 2133
rect -22548 2065 -22482 2099
rect -22548 2031 -22532 2065
rect -22498 2031 -22482 2065
rect -22548 1997 -22482 2031
rect -22548 1963 -22532 1997
rect -22498 1963 -22482 1997
rect -22548 1929 -22482 1963
rect -22548 1895 -22532 1929
rect -22498 1895 -22482 1929
rect -22548 1854 -22482 1895
rect -22452 2813 -22386 2854
rect -22452 2779 -22436 2813
rect -22402 2779 -22386 2813
rect -22452 2745 -22386 2779
rect -22452 2711 -22436 2745
rect -22402 2711 -22386 2745
rect -22452 2677 -22386 2711
rect -22452 2643 -22436 2677
rect -22402 2643 -22386 2677
rect -22452 2609 -22386 2643
rect -22452 2575 -22436 2609
rect -22402 2575 -22386 2609
rect -22452 2541 -22386 2575
rect -22452 2507 -22436 2541
rect -22402 2507 -22386 2541
rect -22452 2473 -22386 2507
rect -22452 2439 -22436 2473
rect -22402 2439 -22386 2473
rect -22452 2405 -22386 2439
rect -22452 2371 -22436 2405
rect -22402 2371 -22386 2405
rect -22452 2337 -22386 2371
rect -22452 2303 -22436 2337
rect -22402 2303 -22386 2337
rect -22452 2269 -22386 2303
rect -22452 2235 -22436 2269
rect -22402 2235 -22386 2269
rect -22452 2201 -22386 2235
rect -22452 2167 -22436 2201
rect -22402 2167 -22386 2201
rect -22452 2133 -22386 2167
rect -22452 2099 -22436 2133
rect -22402 2099 -22386 2133
rect -22452 2065 -22386 2099
rect -22452 2031 -22436 2065
rect -22402 2031 -22386 2065
rect -22452 1997 -22386 2031
rect -22452 1963 -22436 1997
rect -22402 1963 -22386 1997
rect -22452 1929 -22386 1963
rect -22452 1895 -22436 1929
rect -22402 1895 -22386 1929
rect -22452 1854 -22386 1895
rect -22356 2813 -22290 2854
rect -22356 2779 -22340 2813
rect -22306 2779 -22290 2813
rect -22356 2745 -22290 2779
rect -22356 2711 -22340 2745
rect -22306 2711 -22290 2745
rect -22356 2677 -22290 2711
rect -22356 2643 -22340 2677
rect -22306 2643 -22290 2677
rect -22356 2609 -22290 2643
rect -22356 2575 -22340 2609
rect -22306 2575 -22290 2609
rect -22356 2541 -22290 2575
rect -22356 2507 -22340 2541
rect -22306 2507 -22290 2541
rect -22356 2473 -22290 2507
rect -22356 2439 -22340 2473
rect -22306 2439 -22290 2473
rect -22356 2405 -22290 2439
rect -22356 2371 -22340 2405
rect -22306 2371 -22290 2405
rect -22356 2337 -22290 2371
rect -22356 2303 -22340 2337
rect -22306 2303 -22290 2337
rect -22356 2269 -22290 2303
rect -22356 2235 -22340 2269
rect -22306 2235 -22290 2269
rect -22356 2201 -22290 2235
rect -22356 2167 -22340 2201
rect -22306 2167 -22290 2201
rect -22356 2133 -22290 2167
rect -22356 2099 -22340 2133
rect -22306 2099 -22290 2133
rect -22356 2065 -22290 2099
rect -22356 2031 -22340 2065
rect -22306 2031 -22290 2065
rect -22356 1997 -22290 2031
rect -22356 1963 -22340 1997
rect -22306 1963 -22290 1997
rect -22356 1929 -22290 1963
rect -22356 1895 -22340 1929
rect -22306 1895 -22290 1929
rect -22356 1854 -22290 1895
rect -22260 2813 -22194 2854
rect -22260 2779 -22244 2813
rect -22210 2779 -22194 2813
rect -22260 2745 -22194 2779
rect -22260 2711 -22244 2745
rect -22210 2711 -22194 2745
rect -22260 2677 -22194 2711
rect -22260 2643 -22244 2677
rect -22210 2643 -22194 2677
rect -22260 2609 -22194 2643
rect -22260 2575 -22244 2609
rect -22210 2575 -22194 2609
rect -22260 2541 -22194 2575
rect -22260 2507 -22244 2541
rect -22210 2507 -22194 2541
rect -22260 2473 -22194 2507
rect -22260 2439 -22244 2473
rect -22210 2439 -22194 2473
rect -22260 2405 -22194 2439
rect -22260 2371 -22244 2405
rect -22210 2371 -22194 2405
rect -22260 2337 -22194 2371
rect -22260 2303 -22244 2337
rect -22210 2303 -22194 2337
rect -22260 2269 -22194 2303
rect -22260 2235 -22244 2269
rect -22210 2235 -22194 2269
rect -22260 2201 -22194 2235
rect -22260 2167 -22244 2201
rect -22210 2167 -22194 2201
rect -22260 2133 -22194 2167
rect -22260 2099 -22244 2133
rect -22210 2099 -22194 2133
rect -22260 2065 -22194 2099
rect -22260 2031 -22244 2065
rect -22210 2031 -22194 2065
rect -22260 1997 -22194 2031
rect -22260 1963 -22244 1997
rect -22210 1963 -22194 1997
rect -22260 1929 -22194 1963
rect -22260 1895 -22244 1929
rect -22210 1895 -22194 1929
rect -22260 1854 -22194 1895
rect -22164 2813 -22098 2854
rect -22164 2779 -22148 2813
rect -22114 2779 -22098 2813
rect -22164 2745 -22098 2779
rect -22164 2711 -22148 2745
rect -22114 2711 -22098 2745
rect -22164 2677 -22098 2711
rect -22164 2643 -22148 2677
rect -22114 2643 -22098 2677
rect -22164 2609 -22098 2643
rect -22164 2575 -22148 2609
rect -22114 2575 -22098 2609
rect -22164 2541 -22098 2575
rect -22164 2507 -22148 2541
rect -22114 2507 -22098 2541
rect -22164 2473 -22098 2507
rect -22164 2439 -22148 2473
rect -22114 2439 -22098 2473
rect -22164 2405 -22098 2439
rect -22164 2371 -22148 2405
rect -22114 2371 -22098 2405
rect -22164 2337 -22098 2371
rect -22164 2303 -22148 2337
rect -22114 2303 -22098 2337
rect -22164 2269 -22098 2303
rect -22164 2235 -22148 2269
rect -22114 2235 -22098 2269
rect -22164 2201 -22098 2235
rect -22164 2167 -22148 2201
rect -22114 2167 -22098 2201
rect -22164 2133 -22098 2167
rect -22164 2099 -22148 2133
rect -22114 2099 -22098 2133
rect -22164 2065 -22098 2099
rect -22164 2031 -22148 2065
rect -22114 2031 -22098 2065
rect -22164 1997 -22098 2031
rect -22164 1963 -22148 1997
rect -22114 1963 -22098 1997
rect -22164 1929 -22098 1963
rect -22164 1895 -22148 1929
rect -22114 1895 -22098 1929
rect -22164 1854 -22098 1895
rect -22068 2813 -22002 2854
rect -22068 2779 -22052 2813
rect -22018 2779 -22002 2813
rect -22068 2745 -22002 2779
rect -22068 2711 -22052 2745
rect -22018 2711 -22002 2745
rect -22068 2677 -22002 2711
rect -22068 2643 -22052 2677
rect -22018 2643 -22002 2677
rect -22068 2609 -22002 2643
rect -22068 2575 -22052 2609
rect -22018 2575 -22002 2609
rect -22068 2541 -22002 2575
rect -22068 2507 -22052 2541
rect -22018 2507 -22002 2541
rect -22068 2473 -22002 2507
rect -22068 2439 -22052 2473
rect -22018 2439 -22002 2473
rect -22068 2405 -22002 2439
rect -22068 2371 -22052 2405
rect -22018 2371 -22002 2405
rect -22068 2337 -22002 2371
rect -22068 2303 -22052 2337
rect -22018 2303 -22002 2337
rect -22068 2269 -22002 2303
rect -22068 2235 -22052 2269
rect -22018 2235 -22002 2269
rect -22068 2201 -22002 2235
rect -22068 2167 -22052 2201
rect -22018 2167 -22002 2201
rect -22068 2133 -22002 2167
rect -22068 2099 -22052 2133
rect -22018 2099 -22002 2133
rect -22068 2065 -22002 2099
rect -22068 2031 -22052 2065
rect -22018 2031 -22002 2065
rect -22068 1997 -22002 2031
rect -22068 1963 -22052 1997
rect -22018 1963 -22002 1997
rect -22068 1929 -22002 1963
rect -22068 1895 -22052 1929
rect -22018 1895 -22002 1929
rect -22068 1854 -22002 1895
rect -21972 2813 -21906 2854
rect -21972 2779 -21956 2813
rect -21922 2779 -21906 2813
rect -21972 2745 -21906 2779
rect -21972 2711 -21956 2745
rect -21922 2711 -21906 2745
rect -21972 2677 -21906 2711
rect -21972 2643 -21956 2677
rect -21922 2643 -21906 2677
rect -21972 2609 -21906 2643
rect -21972 2575 -21956 2609
rect -21922 2575 -21906 2609
rect -21972 2541 -21906 2575
rect -21972 2507 -21956 2541
rect -21922 2507 -21906 2541
rect -21972 2473 -21906 2507
rect -21972 2439 -21956 2473
rect -21922 2439 -21906 2473
rect -21972 2405 -21906 2439
rect -21972 2371 -21956 2405
rect -21922 2371 -21906 2405
rect -21972 2337 -21906 2371
rect -21972 2303 -21956 2337
rect -21922 2303 -21906 2337
rect -21972 2269 -21906 2303
rect -21972 2235 -21956 2269
rect -21922 2235 -21906 2269
rect -21972 2201 -21906 2235
rect -21972 2167 -21956 2201
rect -21922 2167 -21906 2201
rect -21972 2133 -21906 2167
rect -21972 2099 -21956 2133
rect -21922 2099 -21906 2133
rect -21972 2065 -21906 2099
rect -21972 2031 -21956 2065
rect -21922 2031 -21906 2065
rect -21972 1997 -21906 2031
rect -21972 1963 -21956 1997
rect -21922 1963 -21906 1997
rect -21972 1929 -21906 1963
rect -21972 1895 -21956 1929
rect -21922 1895 -21906 1929
rect -21972 1854 -21906 1895
rect -21876 2813 -21810 2854
rect -21876 2779 -21860 2813
rect -21826 2779 -21810 2813
rect -21876 2745 -21810 2779
rect -21876 2711 -21860 2745
rect -21826 2711 -21810 2745
rect -21876 2677 -21810 2711
rect -21876 2643 -21860 2677
rect -21826 2643 -21810 2677
rect -21876 2609 -21810 2643
rect -21876 2575 -21860 2609
rect -21826 2575 -21810 2609
rect -21876 2541 -21810 2575
rect -21876 2507 -21860 2541
rect -21826 2507 -21810 2541
rect -21876 2473 -21810 2507
rect -21876 2439 -21860 2473
rect -21826 2439 -21810 2473
rect -21876 2405 -21810 2439
rect -21876 2371 -21860 2405
rect -21826 2371 -21810 2405
rect -21876 2337 -21810 2371
rect -21876 2303 -21860 2337
rect -21826 2303 -21810 2337
rect -21876 2269 -21810 2303
rect -21876 2235 -21860 2269
rect -21826 2235 -21810 2269
rect -21876 2201 -21810 2235
rect -21876 2167 -21860 2201
rect -21826 2167 -21810 2201
rect -21876 2133 -21810 2167
rect -21876 2099 -21860 2133
rect -21826 2099 -21810 2133
rect -21876 2065 -21810 2099
rect -21876 2031 -21860 2065
rect -21826 2031 -21810 2065
rect -21876 1997 -21810 2031
rect -21876 1963 -21860 1997
rect -21826 1963 -21810 1997
rect -21876 1929 -21810 1963
rect -21876 1895 -21860 1929
rect -21826 1895 -21810 1929
rect -21876 1854 -21810 1895
rect -21780 2813 -21714 2854
rect -21780 2779 -21764 2813
rect -21730 2779 -21714 2813
rect -21780 2745 -21714 2779
rect -21780 2711 -21764 2745
rect -21730 2711 -21714 2745
rect -21780 2677 -21714 2711
rect -21780 2643 -21764 2677
rect -21730 2643 -21714 2677
rect -21780 2609 -21714 2643
rect -21780 2575 -21764 2609
rect -21730 2575 -21714 2609
rect -21780 2541 -21714 2575
rect -21780 2507 -21764 2541
rect -21730 2507 -21714 2541
rect -21780 2473 -21714 2507
rect -21780 2439 -21764 2473
rect -21730 2439 -21714 2473
rect -21780 2405 -21714 2439
rect -21780 2371 -21764 2405
rect -21730 2371 -21714 2405
rect -21780 2337 -21714 2371
rect -21780 2303 -21764 2337
rect -21730 2303 -21714 2337
rect -21780 2269 -21714 2303
rect -21780 2235 -21764 2269
rect -21730 2235 -21714 2269
rect -21780 2201 -21714 2235
rect -21780 2167 -21764 2201
rect -21730 2167 -21714 2201
rect -21780 2133 -21714 2167
rect -21780 2099 -21764 2133
rect -21730 2099 -21714 2133
rect -21780 2065 -21714 2099
rect -21780 2031 -21764 2065
rect -21730 2031 -21714 2065
rect -21780 1997 -21714 2031
rect -21780 1963 -21764 1997
rect -21730 1963 -21714 1997
rect -21780 1929 -21714 1963
rect -21780 1895 -21764 1929
rect -21730 1895 -21714 1929
rect -21780 1854 -21714 1895
rect -21684 2813 -21618 2854
rect -21684 2779 -21668 2813
rect -21634 2779 -21618 2813
rect -21684 2745 -21618 2779
rect -21684 2711 -21668 2745
rect -21634 2711 -21618 2745
rect -21684 2677 -21618 2711
rect -21684 2643 -21668 2677
rect -21634 2643 -21618 2677
rect -21684 2609 -21618 2643
rect -21684 2575 -21668 2609
rect -21634 2575 -21618 2609
rect -21684 2541 -21618 2575
rect -21684 2507 -21668 2541
rect -21634 2507 -21618 2541
rect -21684 2473 -21618 2507
rect -21684 2439 -21668 2473
rect -21634 2439 -21618 2473
rect -21684 2405 -21618 2439
rect -21684 2371 -21668 2405
rect -21634 2371 -21618 2405
rect -21684 2337 -21618 2371
rect -21684 2303 -21668 2337
rect -21634 2303 -21618 2337
rect -21684 2269 -21618 2303
rect -21684 2235 -21668 2269
rect -21634 2235 -21618 2269
rect -21684 2201 -21618 2235
rect -21684 2167 -21668 2201
rect -21634 2167 -21618 2201
rect -21684 2133 -21618 2167
rect -21684 2099 -21668 2133
rect -21634 2099 -21618 2133
rect -21684 2065 -21618 2099
rect -21684 2031 -21668 2065
rect -21634 2031 -21618 2065
rect -21684 1997 -21618 2031
rect -21684 1963 -21668 1997
rect -21634 1963 -21618 1997
rect -21684 1929 -21618 1963
rect -21684 1895 -21668 1929
rect -21634 1895 -21618 1929
rect -21684 1854 -21618 1895
rect -21588 2813 -21526 2854
rect -1698 3059 -1636 3093
rect -21588 2779 -21572 2813
rect -21538 2779 -21526 2813
rect -21588 2745 -21526 2779
rect -21588 2711 -21572 2745
rect -21538 2711 -21526 2745
rect -21588 2677 -21526 2711
rect -21588 2643 -21572 2677
rect -21538 2643 -21526 2677
rect -21588 2609 -21526 2643
rect -21588 2575 -21572 2609
rect -21538 2575 -21526 2609
rect -21588 2541 -21526 2575
rect -21588 2507 -21572 2541
rect -21538 2507 -21526 2541
rect -21588 2473 -21526 2507
rect -21588 2439 -21572 2473
rect -21538 2439 -21526 2473
rect -21588 2405 -21526 2439
rect -21588 2371 -21572 2405
rect -21538 2371 -21526 2405
rect -21588 2337 -21526 2371
rect -21588 2303 -21572 2337
rect -21538 2303 -21526 2337
rect -21588 2269 -21526 2303
rect -21588 2235 -21572 2269
rect -21538 2235 -21526 2269
rect -21588 2201 -21526 2235
rect -21588 2167 -21572 2201
rect -21538 2167 -21526 2201
rect -21588 2133 -21526 2167
rect -21588 2099 -21572 2133
rect -21538 2099 -21526 2133
rect -21588 2065 -21526 2099
rect -21588 2031 -21572 2065
rect -21538 2031 -21526 2065
rect -21588 1997 -21526 2031
rect -21588 1963 -21572 1997
rect -21538 1963 -21526 1997
rect -21588 1929 -21526 1963
rect -21588 1895 -21572 1929
rect -21538 1895 -21526 1929
rect -21588 1854 -21526 1895
rect -21356 2805 -21294 2846
rect -21356 2771 -21344 2805
rect -21310 2771 -21294 2805
rect -21356 2737 -21294 2771
rect -21356 2703 -21344 2737
rect -21310 2703 -21294 2737
rect -21356 2669 -21294 2703
rect -21356 2635 -21344 2669
rect -21310 2635 -21294 2669
rect -21356 2601 -21294 2635
rect -21356 2567 -21344 2601
rect -21310 2567 -21294 2601
rect -21356 2533 -21294 2567
rect -21356 2499 -21344 2533
rect -21310 2499 -21294 2533
rect -21356 2465 -21294 2499
rect -21356 2431 -21344 2465
rect -21310 2431 -21294 2465
rect -21356 2397 -21294 2431
rect -21356 2363 -21344 2397
rect -21310 2363 -21294 2397
rect -21356 2329 -21294 2363
rect -21356 2295 -21344 2329
rect -21310 2295 -21294 2329
rect -21356 2261 -21294 2295
rect -21356 2227 -21344 2261
rect -21310 2227 -21294 2261
rect -21356 2193 -21294 2227
rect -21356 2159 -21344 2193
rect -21310 2159 -21294 2193
rect -21356 2125 -21294 2159
rect -21356 2091 -21344 2125
rect -21310 2091 -21294 2125
rect -21356 2057 -21294 2091
rect -21356 2023 -21344 2057
rect -21310 2023 -21294 2057
rect -21356 1989 -21294 2023
rect -21356 1955 -21344 1989
rect -21310 1955 -21294 1989
rect -21356 1921 -21294 1955
rect -21356 1887 -21344 1921
rect -21310 1887 -21294 1921
rect -21356 1846 -21294 1887
rect -21264 2805 -21198 2846
rect -21264 2771 -21248 2805
rect -21214 2771 -21198 2805
rect -21264 2737 -21198 2771
rect -21264 2703 -21248 2737
rect -21214 2703 -21198 2737
rect -21264 2669 -21198 2703
rect -21264 2635 -21248 2669
rect -21214 2635 -21198 2669
rect -21264 2601 -21198 2635
rect -21264 2567 -21248 2601
rect -21214 2567 -21198 2601
rect -21264 2533 -21198 2567
rect -21264 2499 -21248 2533
rect -21214 2499 -21198 2533
rect -21264 2465 -21198 2499
rect -21264 2431 -21248 2465
rect -21214 2431 -21198 2465
rect -21264 2397 -21198 2431
rect -21264 2363 -21248 2397
rect -21214 2363 -21198 2397
rect -21264 2329 -21198 2363
rect -21264 2295 -21248 2329
rect -21214 2295 -21198 2329
rect -21264 2261 -21198 2295
rect -21264 2227 -21248 2261
rect -21214 2227 -21198 2261
rect -21264 2193 -21198 2227
rect -21264 2159 -21248 2193
rect -21214 2159 -21198 2193
rect -21264 2125 -21198 2159
rect -21264 2091 -21248 2125
rect -21214 2091 -21198 2125
rect -21264 2057 -21198 2091
rect -21264 2023 -21248 2057
rect -21214 2023 -21198 2057
rect -21264 1989 -21198 2023
rect -21264 1955 -21248 1989
rect -21214 1955 -21198 1989
rect -21264 1921 -21198 1955
rect -21264 1887 -21248 1921
rect -21214 1887 -21198 1921
rect -21264 1846 -21198 1887
rect -21168 2805 -21102 2846
rect -21168 2771 -21152 2805
rect -21118 2771 -21102 2805
rect -21168 2737 -21102 2771
rect -21168 2703 -21152 2737
rect -21118 2703 -21102 2737
rect -21168 2669 -21102 2703
rect -21168 2635 -21152 2669
rect -21118 2635 -21102 2669
rect -21168 2601 -21102 2635
rect -21168 2567 -21152 2601
rect -21118 2567 -21102 2601
rect -21168 2533 -21102 2567
rect -21168 2499 -21152 2533
rect -21118 2499 -21102 2533
rect -21168 2465 -21102 2499
rect -21168 2431 -21152 2465
rect -21118 2431 -21102 2465
rect -21168 2397 -21102 2431
rect -21168 2363 -21152 2397
rect -21118 2363 -21102 2397
rect -21168 2329 -21102 2363
rect -21168 2295 -21152 2329
rect -21118 2295 -21102 2329
rect -21168 2261 -21102 2295
rect -21168 2227 -21152 2261
rect -21118 2227 -21102 2261
rect -21168 2193 -21102 2227
rect -21168 2159 -21152 2193
rect -21118 2159 -21102 2193
rect -21168 2125 -21102 2159
rect -21168 2091 -21152 2125
rect -21118 2091 -21102 2125
rect -21168 2057 -21102 2091
rect -21168 2023 -21152 2057
rect -21118 2023 -21102 2057
rect -21168 1989 -21102 2023
rect -21168 1955 -21152 1989
rect -21118 1955 -21102 1989
rect -21168 1921 -21102 1955
rect -21168 1887 -21152 1921
rect -21118 1887 -21102 1921
rect -21168 1846 -21102 1887
rect -21072 2805 -21006 2846
rect -21072 2771 -21056 2805
rect -21022 2771 -21006 2805
rect -21072 2737 -21006 2771
rect -21072 2703 -21056 2737
rect -21022 2703 -21006 2737
rect -21072 2669 -21006 2703
rect -21072 2635 -21056 2669
rect -21022 2635 -21006 2669
rect -21072 2601 -21006 2635
rect -21072 2567 -21056 2601
rect -21022 2567 -21006 2601
rect -21072 2533 -21006 2567
rect -21072 2499 -21056 2533
rect -21022 2499 -21006 2533
rect -21072 2465 -21006 2499
rect -21072 2431 -21056 2465
rect -21022 2431 -21006 2465
rect -21072 2397 -21006 2431
rect -21072 2363 -21056 2397
rect -21022 2363 -21006 2397
rect -21072 2329 -21006 2363
rect -21072 2295 -21056 2329
rect -21022 2295 -21006 2329
rect -21072 2261 -21006 2295
rect -21072 2227 -21056 2261
rect -21022 2227 -21006 2261
rect -21072 2193 -21006 2227
rect -21072 2159 -21056 2193
rect -21022 2159 -21006 2193
rect -21072 2125 -21006 2159
rect -21072 2091 -21056 2125
rect -21022 2091 -21006 2125
rect -21072 2057 -21006 2091
rect -21072 2023 -21056 2057
rect -21022 2023 -21006 2057
rect -21072 1989 -21006 2023
rect -21072 1955 -21056 1989
rect -21022 1955 -21006 1989
rect -21072 1921 -21006 1955
rect -21072 1887 -21056 1921
rect -21022 1887 -21006 1921
rect -21072 1846 -21006 1887
rect -20976 2805 -20910 2846
rect -20976 2771 -20960 2805
rect -20926 2771 -20910 2805
rect -20976 2737 -20910 2771
rect -20976 2703 -20960 2737
rect -20926 2703 -20910 2737
rect -20976 2669 -20910 2703
rect -20976 2635 -20960 2669
rect -20926 2635 -20910 2669
rect -20976 2601 -20910 2635
rect -20976 2567 -20960 2601
rect -20926 2567 -20910 2601
rect -20976 2533 -20910 2567
rect -20976 2499 -20960 2533
rect -20926 2499 -20910 2533
rect -20976 2465 -20910 2499
rect -20976 2431 -20960 2465
rect -20926 2431 -20910 2465
rect -20976 2397 -20910 2431
rect -20976 2363 -20960 2397
rect -20926 2363 -20910 2397
rect -20976 2329 -20910 2363
rect -20976 2295 -20960 2329
rect -20926 2295 -20910 2329
rect -20976 2261 -20910 2295
rect -20976 2227 -20960 2261
rect -20926 2227 -20910 2261
rect -20976 2193 -20910 2227
rect -20976 2159 -20960 2193
rect -20926 2159 -20910 2193
rect -20976 2125 -20910 2159
rect -20976 2091 -20960 2125
rect -20926 2091 -20910 2125
rect -20976 2057 -20910 2091
rect -20976 2023 -20960 2057
rect -20926 2023 -20910 2057
rect -20976 1989 -20910 2023
rect -20976 1955 -20960 1989
rect -20926 1955 -20910 1989
rect -20976 1921 -20910 1955
rect -20976 1887 -20960 1921
rect -20926 1887 -20910 1921
rect -20976 1846 -20910 1887
rect -20880 2805 -20814 2846
rect -20880 2771 -20864 2805
rect -20830 2771 -20814 2805
rect -20880 2737 -20814 2771
rect -20880 2703 -20864 2737
rect -20830 2703 -20814 2737
rect -20880 2669 -20814 2703
rect -20880 2635 -20864 2669
rect -20830 2635 -20814 2669
rect -20880 2601 -20814 2635
rect -20880 2567 -20864 2601
rect -20830 2567 -20814 2601
rect -20880 2533 -20814 2567
rect -20880 2499 -20864 2533
rect -20830 2499 -20814 2533
rect -20880 2465 -20814 2499
rect -20880 2431 -20864 2465
rect -20830 2431 -20814 2465
rect -20880 2397 -20814 2431
rect -20880 2363 -20864 2397
rect -20830 2363 -20814 2397
rect -20880 2329 -20814 2363
rect -20880 2295 -20864 2329
rect -20830 2295 -20814 2329
rect -20880 2261 -20814 2295
rect -20880 2227 -20864 2261
rect -20830 2227 -20814 2261
rect -20880 2193 -20814 2227
rect -20880 2159 -20864 2193
rect -20830 2159 -20814 2193
rect -20880 2125 -20814 2159
rect -20880 2091 -20864 2125
rect -20830 2091 -20814 2125
rect -20880 2057 -20814 2091
rect -20880 2023 -20864 2057
rect -20830 2023 -20814 2057
rect -20880 1989 -20814 2023
rect -20880 1955 -20864 1989
rect -20830 1955 -20814 1989
rect -20880 1921 -20814 1955
rect -20880 1887 -20864 1921
rect -20830 1887 -20814 1921
rect -20880 1846 -20814 1887
rect -20784 2805 -20718 2846
rect -20784 2771 -20768 2805
rect -20734 2771 -20718 2805
rect -20784 2737 -20718 2771
rect -20784 2703 -20768 2737
rect -20734 2703 -20718 2737
rect -20784 2669 -20718 2703
rect -20784 2635 -20768 2669
rect -20734 2635 -20718 2669
rect -20784 2601 -20718 2635
rect -20784 2567 -20768 2601
rect -20734 2567 -20718 2601
rect -20784 2533 -20718 2567
rect -20784 2499 -20768 2533
rect -20734 2499 -20718 2533
rect -20784 2465 -20718 2499
rect -20784 2431 -20768 2465
rect -20734 2431 -20718 2465
rect -20784 2397 -20718 2431
rect -20784 2363 -20768 2397
rect -20734 2363 -20718 2397
rect -20784 2329 -20718 2363
rect -20784 2295 -20768 2329
rect -20734 2295 -20718 2329
rect -20784 2261 -20718 2295
rect -20784 2227 -20768 2261
rect -20734 2227 -20718 2261
rect -20784 2193 -20718 2227
rect -20784 2159 -20768 2193
rect -20734 2159 -20718 2193
rect -20784 2125 -20718 2159
rect -20784 2091 -20768 2125
rect -20734 2091 -20718 2125
rect -20784 2057 -20718 2091
rect -20784 2023 -20768 2057
rect -20734 2023 -20718 2057
rect -20784 1989 -20718 2023
rect -20784 1955 -20768 1989
rect -20734 1955 -20718 1989
rect -20784 1921 -20718 1955
rect -20784 1887 -20768 1921
rect -20734 1887 -20718 1921
rect -20784 1846 -20718 1887
rect -20688 2805 -20622 2846
rect -20688 2771 -20672 2805
rect -20638 2771 -20622 2805
rect -20688 2737 -20622 2771
rect -20688 2703 -20672 2737
rect -20638 2703 -20622 2737
rect -20688 2669 -20622 2703
rect -20688 2635 -20672 2669
rect -20638 2635 -20622 2669
rect -20688 2601 -20622 2635
rect -20688 2567 -20672 2601
rect -20638 2567 -20622 2601
rect -20688 2533 -20622 2567
rect -20688 2499 -20672 2533
rect -20638 2499 -20622 2533
rect -20688 2465 -20622 2499
rect -20688 2431 -20672 2465
rect -20638 2431 -20622 2465
rect -20688 2397 -20622 2431
rect -20688 2363 -20672 2397
rect -20638 2363 -20622 2397
rect -20688 2329 -20622 2363
rect -20688 2295 -20672 2329
rect -20638 2295 -20622 2329
rect -20688 2261 -20622 2295
rect -20688 2227 -20672 2261
rect -20638 2227 -20622 2261
rect -20688 2193 -20622 2227
rect -20688 2159 -20672 2193
rect -20638 2159 -20622 2193
rect -20688 2125 -20622 2159
rect -20688 2091 -20672 2125
rect -20638 2091 -20622 2125
rect -20688 2057 -20622 2091
rect -20688 2023 -20672 2057
rect -20638 2023 -20622 2057
rect -20688 1989 -20622 2023
rect -20688 1955 -20672 1989
rect -20638 1955 -20622 1989
rect -20688 1921 -20622 1955
rect -20688 1887 -20672 1921
rect -20638 1887 -20622 1921
rect -20688 1846 -20622 1887
rect -20592 2805 -20526 2846
rect -20592 2771 -20576 2805
rect -20542 2771 -20526 2805
rect -20592 2737 -20526 2771
rect -20592 2703 -20576 2737
rect -20542 2703 -20526 2737
rect -20592 2669 -20526 2703
rect -20592 2635 -20576 2669
rect -20542 2635 -20526 2669
rect -20592 2601 -20526 2635
rect -20592 2567 -20576 2601
rect -20542 2567 -20526 2601
rect -20592 2533 -20526 2567
rect -20592 2499 -20576 2533
rect -20542 2499 -20526 2533
rect -20592 2465 -20526 2499
rect -20592 2431 -20576 2465
rect -20542 2431 -20526 2465
rect -20592 2397 -20526 2431
rect -20592 2363 -20576 2397
rect -20542 2363 -20526 2397
rect -20592 2329 -20526 2363
rect -20592 2295 -20576 2329
rect -20542 2295 -20526 2329
rect -20592 2261 -20526 2295
rect -20592 2227 -20576 2261
rect -20542 2227 -20526 2261
rect -20592 2193 -20526 2227
rect -20592 2159 -20576 2193
rect -20542 2159 -20526 2193
rect -20592 2125 -20526 2159
rect -20592 2091 -20576 2125
rect -20542 2091 -20526 2125
rect -20592 2057 -20526 2091
rect -20592 2023 -20576 2057
rect -20542 2023 -20526 2057
rect -20592 1989 -20526 2023
rect -20592 1955 -20576 1989
rect -20542 1955 -20526 1989
rect -20592 1921 -20526 1955
rect -20592 1887 -20576 1921
rect -20542 1887 -20526 1921
rect -20592 1846 -20526 1887
rect -20496 2805 -20430 2846
rect -20496 2771 -20480 2805
rect -20446 2771 -20430 2805
rect -20496 2737 -20430 2771
rect -20496 2703 -20480 2737
rect -20446 2703 -20430 2737
rect -20496 2669 -20430 2703
rect -20496 2635 -20480 2669
rect -20446 2635 -20430 2669
rect -20496 2601 -20430 2635
rect -20496 2567 -20480 2601
rect -20446 2567 -20430 2601
rect -20496 2533 -20430 2567
rect -20496 2499 -20480 2533
rect -20446 2499 -20430 2533
rect -20496 2465 -20430 2499
rect -20496 2431 -20480 2465
rect -20446 2431 -20430 2465
rect -20496 2397 -20430 2431
rect -20496 2363 -20480 2397
rect -20446 2363 -20430 2397
rect -20496 2329 -20430 2363
rect -20496 2295 -20480 2329
rect -20446 2295 -20430 2329
rect -20496 2261 -20430 2295
rect -20496 2227 -20480 2261
rect -20446 2227 -20430 2261
rect -20496 2193 -20430 2227
rect -20496 2159 -20480 2193
rect -20446 2159 -20430 2193
rect -20496 2125 -20430 2159
rect -20496 2091 -20480 2125
rect -20446 2091 -20430 2125
rect -20496 2057 -20430 2091
rect -20496 2023 -20480 2057
rect -20446 2023 -20430 2057
rect -20496 1989 -20430 2023
rect -20496 1955 -20480 1989
rect -20446 1955 -20430 1989
rect -20496 1921 -20430 1955
rect -20496 1887 -20480 1921
rect -20446 1887 -20430 1921
rect -20496 1846 -20430 1887
rect -20400 2805 -20334 2846
rect -20400 2771 -20384 2805
rect -20350 2771 -20334 2805
rect -20400 2737 -20334 2771
rect -20400 2703 -20384 2737
rect -20350 2703 -20334 2737
rect -20400 2669 -20334 2703
rect -20400 2635 -20384 2669
rect -20350 2635 -20334 2669
rect -20400 2601 -20334 2635
rect -20400 2567 -20384 2601
rect -20350 2567 -20334 2601
rect -20400 2533 -20334 2567
rect -20400 2499 -20384 2533
rect -20350 2499 -20334 2533
rect -20400 2465 -20334 2499
rect -20400 2431 -20384 2465
rect -20350 2431 -20334 2465
rect -20400 2397 -20334 2431
rect -20400 2363 -20384 2397
rect -20350 2363 -20334 2397
rect -20400 2329 -20334 2363
rect -20400 2295 -20384 2329
rect -20350 2295 -20334 2329
rect -20400 2261 -20334 2295
rect -20400 2227 -20384 2261
rect -20350 2227 -20334 2261
rect -20400 2193 -20334 2227
rect -20400 2159 -20384 2193
rect -20350 2159 -20334 2193
rect -20400 2125 -20334 2159
rect -20400 2091 -20384 2125
rect -20350 2091 -20334 2125
rect -20400 2057 -20334 2091
rect -20400 2023 -20384 2057
rect -20350 2023 -20334 2057
rect -20400 1989 -20334 2023
rect -20400 1955 -20384 1989
rect -20350 1955 -20334 1989
rect -20400 1921 -20334 1955
rect -20400 1887 -20384 1921
rect -20350 1887 -20334 1921
rect -20400 1846 -20334 1887
rect -20304 2805 -20238 2846
rect -20304 2771 -20288 2805
rect -20254 2771 -20238 2805
rect -20304 2737 -20238 2771
rect -20304 2703 -20288 2737
rect -20254 2703 -20238 2737
rect -20304 2669 -20238 2703
rect -20304 2635 -20288 2669
rect -20254 2635 -20238 2669
rect -20304 2601 -20238 2635
rect -20304 2567 -20288 2601
rect -20254 2567 -20238 2601
rect -20304 2533 -20238 2567
rect -20304 2499 -20288 2533
rect -20254 2499 -20238 2533
rect -20304 2465 -20238 2499
rect -20304 2431 -20288 2465
rect -20254 2431 -20238 2465
rect -20304 2397 -20238 2431
rect -20304 2363 -20288 2397
rect -20254 2363 -20238 2397
rect -20304 2329 -20238 2363
rect -20304 2295 -20288 2329
rect -20254 2295 -20238 2329
rect -20304 2261 -20238 2295
rect -20304 2227 -20288 2261
rect -20254 2227 -20238 2261
rect -20304 2193 -20238 2227
rect -20304 2159 -20288 2193
rect -20254 2159 -20238 2193
rect -20304 2125 -20238 2159
rect -20304 2091 -20288 2125
rect -20254 2091 -20238 2125
rect -20304 2057 -20238 2091
rect -20304 2023 -20288 2057
rect -20254 2023 -20238 2057
rect -20304 1989 -20238 2023
rect -20304 1955 -20288 1989
rect -20254 1955 -20238 1989
rect -20304 1921 -20238 1955
rect -20304 1887 -20288 1921
rect -20254 1887 -20238 1921
rect -20304 1846 -20238 1887
rect -20208 2805 -20142 2846
rect -20208 2771 -20192 2805
rect -20158 2771 -20142 2805
rect -20208 2737 -20142 2771
rect -20208 2703 -20192 2737
rect -20158 2703 -20142 2737
rect -20208 2669 -20142 2703
rect -20208 2635 -20192 2669
rect -20158 2635 -20142 2669
rect -20208 2601 -20142 2635
rect -20208 2567 -20192 2601
rect -20158 2567 -20142 2601
rect -20208 2533 -20142 2567
rect -20208 2499 -20192 2533
rect -20158 2499 -20142 2533
rect -20208 2465 -20142 2499
rect -20208 2431 -20192 2465
rect -20158 2431 -20142 2465
rect -20208 2397 -20142 2431
rect -20208 2363 -20192 2397
rect -20158 2363 -20142 2397
rect -20208 2329 -20142 2363
rect -20208 2295 -20192 2329
rect -20158 2295 -20142 2329
rect -20208 2261 -20142 2295
rect -20208 2227 -20192 2261
rect -20158 2227 -20142 2261
rect -20208 2193 -20142 2227
rect -20208 2159 -20192 2193
rect -20158 2159 -20142 2193
rect -20208 2125 -20142 2159
rect -20208 2091 -20192 2125
rect -20158 2091 -20142 2125
rect -20208 2057 -20142 2091
rect -20208 2023 -20192 2057
rect -20158 2023 -20142 2057
rect -20208 1989 -20142 2023
rect -20208 1955 -20192 1989
rect -20158 1955 -20142 1989
rect -20208 1921 -20142 1955
rect -20208 1887 -20192 1921
rect -20158 1887 -20142 1921
rect -20208 1846 -20142 1887
rect -20112 2805 -20046 2846
rect -20112 2771 -20096 2805
rect -20062 2771 -20046 2805
rect -20112 2737 -20046 2771
rect -20112 2703 -20096 2737
rect -20062 2703 -20046 2737
rect -20112 2669 -20046 2703
rect -20112 2635 -20096 2669
rect -20062 2635 -20046 2669
rect -20112 2601 -20046 2635
rect -20112 2567 -20096 2601
rect -20062 2567 -20046 2601
rect -20112 2533 -20046 2567
rect -20112 2499 -20096 2533
rect -20062 2499 -20046 2533
rect -20112 2465 -20046 2499
rect -20112 2431 -20096 2465
rect -20062 2431 -20046 2465
rect -20112 2397 -20046 2431
rect -20112 2363 -20096 2397
rect -20062 2363 -20046 2397
rect -20112 2329 -20046 2363
rect -20112 2295 -20096 2329
rect -20062 2295 -20046 2329
rect -20112 2261 -20046 2295
rect -20112 2227 -20096 2261
rect -20062 2227 -20046 2261
rect -20112 2193 -20046 2227
rect -20112 2159 -20096 2193
rect -20062 2159 -20046 2193
rect -20112 2125 -20046 2159
rect -20112 2091 -20096 2125
rect -20062 2091 -20046 2125
rect -20112 2057 -20046 2091
rect -20112 2023 -20096 2057
rect -20062 2023 -20046 2057
rect -20112 1989 -20046 2023
rect -20112 1955 -20096 1989
rect -20062 1955 -20046 1989
rect -20112 1921 -20046 1955
rect -20112 1887 -20096 1921
rect -20062 1887 -20046 1921
rect -20112 1846 -20046 1887
rect -20016 2805 -19950 2846
rect -20016 2771 -20000 2805
rect -19966 2771 -19950 2805
rect -20016 2737 -19950 2771
rect -20016 2703 -20000 2737
rect -19966 2703 -19950 2737
rect -20016 2669 -19950 2703
rect -20016 2635 -20000 2669
rect -19966 2635 -19950 2669
rect -20016 2601 -19950 2635
rect -20016 2567 -20000 2601
rect -19966 2567 -19950 2601
rect -20016 2533 -19950 2567
rect -20016 2499 -20000 2533
rect -19966 2499 -19950 2533
rect -20016 2465 -19950 2499
rect -20016 2431 -20000 2465
rect -19966 2431 -19950 2465
rect -20016 2397 -19950 2431
rect -20016 2363 -20000 2397
rect -19966 2363 -19950 2397
rect -20016 2329 -19950 2363
rect -20016 2295 -20000 2329
rect -19966 2295 -19950 2329
rect -20016 2261 -19950 2295
rect -20016 2227 -20000 2261
rect -19966 2227 -19950 2261
rect -20016 2193 -19950 2227
rect -20016 2159 -20000 2193
rect -19966 2159 -19950 2193
rect -20016 2125 -19950 2159
rect -20016 2091 -20000 2125
rect -19966 2091 -19950 2125
rect -20016 2057 -19950 2091
rect -20016 2023 -20000 2057
rect -19966 2023 -19950 2057
rect -20016 1989 -19950 2023
rect -20016 1955 -20000 1989
rect -19966 1955 -19950 1989
rect -20016 1921 -19950 1955
rect -20016 1887 -20000 1921
rect -19966 1887 -19950 1921
rect -20016 1846 -19950 1887
rect -19920 2805 -19858 2846
rect -19920 2771 -19904 2805
rect -19870 2771 -19858 2805
rect -19920 2737 -19858 2771
rect -19920 2703 -19904 2737
rect -19870 2703 -19858 2737
rect -19920 2669 -19858 2703
rect -19920 2635 -19904 2669
rect -19870 2635 -19858 2669
rect -19920 2601 -19858 2635
rect -19920 2567 -19904 2601
rect -19870 2567 -19858 2601
rect -19920 2533 -19858 2567
rect -19920 2499 -19904 2533
rect -19870 2499 -19858 2533
rect -19920 2465 -19858 2499
rect -19920 2431 -19904 2465
rect -19870 2431 -19858 2465
rect -19920 2397 -19858 2431
rect -19920 2363 -19904 2397
rect -19870 2363 -19858 2397
rect -19920 2329 -19858 2363
rect -19920 2295 -19904 2329
rect -19870 2295 -19858 2329
rect -19920 2261 -19858 2295
rect -19920 2227 -19904 2261
rect -19870 2227 -19858 2261
rect -19920 2193 -19858 2227
rect -19920 2159 -19904 2193
rect -19870 2159 -19858 2193
rect -19920 2125 -19858 2159
rect -19920 2091 -19904 2125
rect -19870 2091 -19858 2125
rect -19920 2057 -19858 2091
rect -19920 2023 -19904 2057
rect -19870 2023 -19858 2057
rect -19920 1989 -19858 2023
rect -19920 1955 -19904 1989
rect -19870 1955 -19858 1989
rect -19920 1921 -19858 1955
rect -19920 1887 -19904 1921
rect -19870 1887 -19858 1921
rect -19920 1846 -19858 1887
rect -19678 2809 -19616 2850
rect -19678 2775 -19666 2809
rect -19632 2775 -19616 2809
rect -19678 2741 -19616 2775
rect -19678 2707 -19666 2741
rect -19632 2707 -19616 2741
rect -19678 2673 -19616 2707
rect -19678 2639 -19666 2673
rect -19632 2639 -19616 2673
rect -19678 2605 -19616 2639
rect -19678 2571 -19666 2605
rect -19632 2571 -19616 2605
rect -19678 2537 -19616 2571
rect -19678 2503 -19666 2537
rect -19632 2503 -19616 2537
rect -19678 2469 -19616 2503
rect -19678 2435 -19666 2469
rect -19632 2435 -19616 2469
rect -19678 2401 -19616 2435
rect -19678 2367 -19666 2401
rect -19632 2367 -19616 2401
rect -19678 2333 -19616 2367
rect -19678 2299 -19666 2333
rect -19632 2299 -19616 2333
rect -19678 2265 -19616 2299
rect -19678 2231 -19666 2265
rect -19632 2231 -19616 2265
rect -19678 2197 -19616 2231
rect -19678 2163 -19666 2197
rect -19632 2163 -19616 2197
rect -19678 2129 -19616 2163
rect -19678 2095 -19666 2129
rect -19632 2095 -19616 2129
rect -19678 2061 -19616 2095
rect -19678 2027 -19666 2061
rect -19632 2027 -19616 2061
rect -19678 1993 -19616 2027
rect -19678 1959 -19666 1993
rect -19632 1959 -19616 1993
rect -19678 1925 -19616 1959
rect -19678 1891 -19666 1925
rect -19632 1891 -19616 1925
rect -19678 1850 -19616 1891
rect -19586 2809 -19520 2850
rect -19586 2775 -19570 2809
rect -19536 2775 -19520 2809
rect -19586 2741 -19520 2775
rect -19586 2707 -19570 2741
rect -19536 2707 -19520 2741
rect -19586 2673 -19520 2707
rect -19586 2639 -19570 2673
rect -19536 2639 -19520 2673
rect -19586 2605 -19520 2639
rect -19586 2571 -19570 2605
rect -19536 2571 -19520 2605
rect -19586 2537 -19520 2571
rect -19586 2503 -19570 2537
rect -19536 2503 -19520 2537
rect -19586 2469 -19520 2503
rect -19586 2435 -19570 2469
rect -19536 2435 -19520 2469
rect -19586 2401 -19520 2435
rect -19586 2367 -19570 2401
rect -19536 2367 -19520 2401
rect -19586 2333 -19520 2367
rect -19586 2299 -19570 2333
rect -19536 2299 -19520 2333
rect -19586 2265 -19520 2299
rect -19586 2231 -19570 2265
rect -19536 2231 -19520 2265
rect -19586 2197 -19520 2231
rect -19586 2163 -19570 2197
rect -19536 2163 -19520 2197
rect -19586 2129 -19520 2163
rect -19586 2095 -19570 2129
rect -19536 2095 -19520 2129
rect -19586 2061 -19520 2095
rect -19586 2027 -19570 2061
rect -19536 2027 -19520 2061
rect -19586 1993 -19520 2027
rect -19586 1959 -19570 1993
rect -19536 1959 -19520 1993
rect -19586 1925 -19520 1959
rect -19586 1891 -19570 1925
rect -19536 1891 -19520 1925
rect -19586 1850 -19520 1891
rect -19490 2809 -19424 2850
rect -19490 2775 -19474 2809
rect -19440 2775 -19424 2809
rect -19490 2741 -19424 2775
rect -19490 2707 -19474 2741
rect -19440 2707 -19424 2741
rect -19490 2673 -19424 2707
rect -19490 2639 -19474 2673
rect -19440 2639 -19424 2673
rect -19490 2605 -19424 2639
rect -19490 2571 -19474 2605
rect -19440 2571 -19424 2605
rect -19490 2537 -19424 2571
rect -19490 2503 -19474 2537
rect -19440 2503 -19424 2537
rect -19490 2469 -19424 2503
rect -19490 2435 -19474 2469
rect -19440 2435 -19424 2469
rect -19490 2401 -19424 2435
rect -19490 2367 -19474 2401
rect -19440 2367 -19424 2401
rect -19490 2333 -19424 2367
rect -19490 2299 -19474 2333
rect -19440 2299 -19424 2333
rect -19490 2265 -19424 2299
rect -19490 2231 -19474 2265
rect -19440 2231 -19424 2265
rect -19490 2197 -19424 2231
rect -19490 2163 -19474 2197
rect -19440 2163 -19424 2197
rect -19490 2129 -19424 2163
rect -19490 2095 -19474 2129
rect -19440 2095 -19424 2129
rect -19490 2061 -19424 2095
rect -19490 2027 -19474 2061
rect -19440 2027 -19424 2061
rect -19490 1993 -19424 2027
rect -19490 1959 -19474 1993
rect -19440 1959 -19424 1993
rect -19490 1925 -19424 1959
rect -19490 1891 -19474 1925
rect -19440 1891 -19424 1925
rect -19490 1850 -19424 1891
rect -19394 2809 -19328 2850
rect -19394 2775 -19378 2809
rect -19344 2775 -19328 2809
rect -19394 2741 -19328 2775
rect -19394 2707 -19378 2741
rect -19344 2707 -19328 2741
rect -19394 2673 -19328 2707
rect -19394 2639 -19378 2673
rect -19344 2639 -19328 2673
rect -19394 2605 -19328 2639
rect -19394 2571 -19378 2605
rect -19344 2571 -19328 2605
rect -19394 2537 -19328 2571
rect -19394 2503 -19378 2537
rect -19344 2503 -19328 2537
rect -19394 2469 -19328 2503
rect -19394 2435 -19378 2469
rect -19344 2435 -19328 2469
rect -19394 2401 -19328 2435
rect -19394 2367 -19378 2401
rect -19344 2367 -19328 2401
rect -19394 2333 -19328 2367
rect -19394 2299 -19378 2333
rect -19344 2299 -19328 2333
rect -19394 2265 -19328 2299
rect -19394 2231 -19378 2265
rect -19344 2231 -19328 2265
rect -19394 2197 -19328 2231
rect -19394 2163 -19378 2197
rect -19344 2163 -19328 2197
rect -19394 2129 -19328 2163
rect -19394 2095 -19378 2129
rect -19344 2095 -19328 2129
rect -19394 2061 -19328 2095
rect -19394 2027 -19378 2061
rect -19344 2027 -19328 2061
rect -19394 1993 -19328 2027
rect -19394 1959 -19378 1993
rect -19344 1959 -19328 1993
rect -19394 1925 -19328 1959
rect -19394 1891 -19378 1925
rect -19344 1891 -19328 1925
rect -19394 1850 -19328 1891
rect -19298 2809 -19232 2850
rect -19298 2775 -19282 2809
rect -19248 2775 -19232 2809
rect -19298 2741 -19232 2775
rect -19298 2707 -19282 2741
rect -19248 2707 -19232 2741
rect -19298 2673 -19232 2707
rect -19298 2639 -19282 2673
rect -19248 2639 -19232 2673
rect -19298 2605 -19232 2639
rect -19298 2571 -19282 2605
rect -19248 2571 -19232 2605
rect -19298 2537 -19232 2571
rect -19298 2503 -19282 2537
rect -19248 2503 -19232 2537
rect -19298 2469 -19232 2503
rect -19298 2435 -19282 2469
rect -19248 2435 -19232 2469
rect -19298 2401 -19232 2435
rect -19298 2367 -19282 2401
rect -19248 2367 -19232 2401
rect -19298 2333 -19232 2367
rect -19298 2299 -19282 2333
rect -19248 2299 -19232 2333
rect -19298 2265 -19232 2299
rect -19298 2231 -19282 2265
rect -19248 2231 -19232 2265
rect -19298 2197 -19232 2231
rect -19298 2163 -19282 2197
rect -19248 2163 -19232 2197
rect -19298 2129 -19232 2163
rect -19298 2095 -19282 2129
rect -19248 2095 -19232 2129
rect -19298 2061 -19232 2095
rect -19298 2027 -19282 2061
rect -19248 2027 -19232 2061
rect -19298 1993 -19232 2027
rect -19298 1959 -19282 1993
rect -19248 1959 -19232 1993
rect -19298 1925 -19232 1959
rect -19298 1891 -19282 1925
rect -19248 1891 -19232 1925
rect -19298 1850 -19232 1891
rect -19202 2809 -19136 2850
rect -19202 2775 -19186 2809
rect -19152 2775 -19136 2809
rect -19202 2741 -19136 2775
rect -19202 2707 -19186 2741
rect -19152 2707 -19136 2741
rect -19202 2673 -19136 2707
rect -19202 2639 -19186 2673
rect -19152 2639 -19136 2673
rect -19202 2605 -19136 2639
rect -19202 2571 -19186 2605
rect -19152 2571 -19136 2605
rect -19202 2537 -19136 2571
rect -19202 2503 -19186 2537
rect -19152 2503 -19136 2537
rect -19202 2469 -19136 2503
rect -19202 2435 -19186 2469
rect -19152 2435 -19136 2469
rect -19202 2401 -19136 2435
rect -19202 2367 -19186 2401
rect -19152 2367 -19136 2401
rect -19202 2333 -19136 2367
rect -19202 2299 -19186 2333
rect -19152 2299 -19136 2333
rect -19202 2265 -19136 2299
rect -19202 2231 -19186 2265
rect -19152 2231 -19136 2265
rect -19202 2197 -19136 2231
rect -19202 2163 -19186 2197
rect -19152 2163 -19136 2197
rect -19202 2129 -19136 2163
rect -19202 2095 -19186 2129
rect -19152 2095 -19136 2129
rect -19202 2061 -19136 2095
rect -19202 2027 -19186 2061
rect -19152 2027 -19136 2061
rect -19202 1993 -19136 2027
rect -19202 1959 -19186 1993
rect -19152 1959 -19136 1993
rect -19202 1925 -19136 1959
rect -19202 1891 -19186 1925
rect -19152 1891 -19136 1925
rect -19202 1850 -19136 1891
rect -19106 2809 -19040 2850
rect -19106 2775 -19090 2809
rect -19056 2775 -19040 2809
rect -19106 2741 -19040 2775
rect -19106 2707 -19090 2741
rect -19056 2707 -19040 2741
rect -19106 2673 -19040 2707
rect -19106 2639 -19090 2673
rect -19056 2639 -19040 2673
rect -19106 2605 -19040 2639
rect -19106 2571 -19090 2605
rect -19056 2571 -19040 2605
rect -19106 2537 -19040 2571
rect -19106 2503 -19090 2537
rect -19056 2503 -19040 2537
rect -19106 2469 -19040 2503
rect -19106 2435 -19090 2469
rect -19056 2435 -19040 2469
rect -19106 2401 -19040 2435
rect -19106 2367 -19090 2401
rect -19056 2367 -19040 2401
rect -19106 2333 -19040 2367
rect -19106 2299 -19090 2333
rect -19056 2299 -19040 2333
rect -19106 2265 -19040 2299
rect -19106 2231 -19090 2265
rect -19056 2231 -19040 2265
rect -19106 2197 -19040 2231
rect -19106 2163 -19090 2197
rect -19056 2163 -19040 2197
rect -19106 2129 -19040 2163
rect -19106 2095 -19090 2129
rect -19056 2095 -19040 2129
rect -19106 2061 -19040 2095
rect -19106 2027 -19090 2061
rect -19056 2027 -19040 2061
rect -19106 1993 -19040 2027
rect -19106 1959 -19090 1993
rect -19056 1959 -19040 1993
rect -19106 1925 -19040 1959
rect -19106 1891 -19090 1925
rect -19056 1891 -19040 1925
rect -19106 1850 -19040 1891
rect -19010 2809 -18944 2850
rect -19010 2775 -18994 2809
rect -18960 2775 -18944 2809
rect -19010 2741 -18944 2775
rect -19010 2707 -18994 2741
rect -18960 2707 -18944 2741
rect -19010 2673 -18944 2707
rect -19010 2639 -18994 2673
rect -18960 2639 -18944 2673
rect -19010 2605 -18944 2639
rect -19010 2571 -18994 2605
rect -18960 2571 -18944 2605
rect -19010 2537 -18944 2571
rect -19010 2503 -18994 2537
rect -18960 2503 -18944 2537
rect -19010 2469 -18944 2503
rect -19010 2435 -18994 2469
rect -18960 2435 -18944 2469
rect -19010 2401 -18944 2435
rect -19010 2367 -18994 2401
rect -18960 2367 -18944 2401
rect -19010 2333 -18944 2367
rect -19010 2299 -18994 2333
rect -18960 2299 -18944 2333
rect -19010 2265 -18944 2299
rect -19010 2231 -18994 2265
rect -18960 2231 -18944 2265
rect -19010 2197 -18944 2231
rect -19010 2163 -18994 2197
rect -18960 2163 -18944 2197
rect -19010 2129 -18944 2163
rect -19010 2095 -18994 2129
rect -18960 2095 -18944 2129
rect -19010 2061 -18944 2095
rect -19010 2027 -18994 2061
rect -18960 2027 -18944 2061
rect -19010 1993 -18944 2027
rect -19010 1959 -18994 1993
rect -18960 1959 -18944 1993
rect -19010 1925 -18944 1959
rect -19010 1891 -18994 1925
rect -18960 1891 -18944 1925
rect -19010 1850 -18944 1891
rect -18914 2809 -18848 2850
rect -18914 2775 -18898 2809
rect -18864 2775 -18848 2809
rect -18914 2741 -18848 2775
rect -18914 2707 -18898 2741
rect -18864 2707 -18848 2741
rect -18914 2673 -18848 2707
rect -18914 2639 -18898 2673
rect -18864 2639 -18848 2673
rect -18914 2605 -18848 2639
rect -18914 2571 -18898 2605
rect -18864 2571 -18848 2605
rect -18914 2537 -18848 2571
rect -18914 2503 -18898 2537
rect -18864 2503 -18848 2537
rect -18914 2469 -18848 2503
rect -18914 2435 -18898 2469
rect -18864 2435 -18848 2469
rect -18914 2401 -18848 2435
rect -18914 2367 -18898 2401
rect -18864 2367 -18848 2401
rect -18914 2333 -18848 2367
rect -18914 2299 -18898 2333
rect -18864 2299 -18848 2333
rect -18914 2265 -18848 2299
rect -18914 2231 -18898 2265
rect -18864 2231 -18848 2265
rect -18914 2197 -18848 2231
rect -18914 2163 -18898 2197
rect -18864 2163 -18848 2197
rect -18914 2129 -18848 2163
rect -18914 2095 -18898 2129
rect -18864 2095 -18848 2129
rect -18914 2061 -18848 2095
rect -18914 2027 -18898 2061
rect -18864 2027 -18848 2061
rect -18914 1993 -18848 2027
rect -18914 1959 -18898 1993
rect -18864 1959 -18848 1993
rect -18914 1925 -18848 1959
rect -18914 1891 -18898 1925
rect -18864 1891 -18848 1925
rect -18914 1850 -18848 1891
rect -18818 2809 -18752 2850
rect -18818 2775 -18802 2809
rect -18768 2775 -18752 2809
rect -18818 2741 -18752 2775
rect -18818 2707 -18802 2741
rect -18768 2707 -18752 2741
rect -18818 2673 -18752 2707
rect -18818 2639 -18802 2673
rect -18768 2639 -18752 2673
rect -18818 2605 -18752 2639
rect -18818 2571 -18802 2605
rect -18768 2571 -18752 2605
rect -18818 2537 -18752 2571
rect -18818 2503 -18802 2537
rect -18768 2503 -18752 2537
rect -18818 2469 -18752 2503
rect -18818 2435 -18802 2469
rect -18768 2435 -18752 2469
rect -18818 2401 -18752 2435
rect -18818 2367 -18802 2401
rect -18768 2367 -18752 2401
rect -18818 2333 -18752 2367
rect -18818 2299 -18802 2333
rect -18768 2299 -18752 2333
rect -18818 2265 -18752 2299
rect -18818 2231 -18802 2265
rect -18768 2231 -18752 2265
rect -18818 2197 -18752 2231
rect -18818 2163 -18802 2197
rect -18768 2163 -18752 2197
rect -18818 2129 -18752 2163
rect -18818 2095 -18802 2129
rect -18768 2095 -18752 2129
rect -18818 2061 -18752 2095
rect -18818 2027 -18802 2061
rect -18768 2027 -18752 2061
rect -18818 1993 -18752 2027
rect -18818 1959 -18802 1993
rect -18768 1959 -18752 1993
rect -18818 1925 -18752 1959
rect -18818 1891 -18802 1925
rect -18768 1891 -18752 1925
rect -18818 1850 -18752 1891
rect -18722 2809 -18660 2850
rect -18722 2775 -18706 2809
rect -18672 2775 -18660 2809
rect -18722 2741 -18660 2775
rect -18722 2707 -18706 2741
rect -18672 2707 -18660 2741
rect -18722 2673 -18660 2707
rect -18722 2639 -18706 2673
rect -18672 2639 -18660 2673
rect -18722 2605 -18660 2639
rect -18722 2571 -18706 2605
rect -18672 2571 -18660 2605
rect -18722 2537 -18660 2571
rect -18722 2503 -18706 2537
rect -18672 2503 -18660 2537
rect -18722 2469 -18660 2503
rect -18722 2435 -18706 2469
rect -18672 2435 -18660 2469
rect -18722 2401 -18660 2435
rect -18722 2367 -18706 2401
rect -18672 2367 -18660 2401
rect -18722 2333 -18660 2367
rect -18722 2299 -18706 2333
rect -18672 2299 -18660 2333
rect -18722 2265 -18660 2299
rect -18722 2231 -18706 2265
rect -18672 2231 -18660 2265
rect -18722 2197 -18660 2231
rect -18722 2163 -18706 2197
rect -18672 2163 -18660 2197
rect -18722 2129 -18660 2163
rect -18722 2095 -18706 2129
rect -18672 2095 -18660 2129
rect -18722 2061 -18660 2095
rect -18722 2027 -18706 2061
rect -18672 2027 -18660 2061
rect -18722 1993 -18660 2027
rect -18722 1959 -18706 1993
rect -18672 1959 -18660 1993
rect -18722 1925 -18660 1959
rect -18722 1891 -18706 1925
rect -18672 1891 -18660 1925
rect -18722 1850 -18660 1891
rect -18506 2819 -18444 2860
rect -18506 2785 -18494 2819
rect -18460 2785 -18444 2819
rect -18506 2751 -18444 2785
rect -18506 2717 -18494 2751
rect -18460 2717 -18444 2751
rect -18506 2683 -18444 2717
rect -18506 2649 -18494 2683
rect -18460 2649 -18444 2683
rect -18506 2615 -18444 2649
rect -18506 2581 -18494 2615
rect -18460 2581 -18444 2615
rect -18506 2547 -18444 2581
rect -18506 2513 -18494 2547
rect -18460 2513 -18444 2547
rect -18506 2479 -18444 2513
rect -18506 2445 -18494 2479
rect -18460 2445 -18444 2479
rect -18506 2411 -18444 2445
rect -18506 2377 -18494 2411
rect -18460 2377 -18444 2411
rect -18506 2343 -18444 2377
rect -18506 2309 -18494 2343
rect -18460 2309 -18444 2343
rect -18506 2275 -18444 2309
rect -18506 2241 -18494 2275
rect -18460 2241 -18444 2275
rect -18506 2207 -18444 2241
rect -18506 2173 -18494 2207
rect -18460 2173 -18444 2207
rect -18506 2139 -18444 2173
rect -18506 2105 -18494 2139
rect -18460 2105 -18444 2139
rect -18506 2071 -18444 2105
rect -18506 2037 -18494 2071
rect -18460 2037 -18444 2071
rect -18506 2003 -18444 2037
rect -18506 1969 -18494 2003
rect -18460 1969 -18444 2003
rect -18506 1935 -18444 1969
rect -18506 1901 -18494 1935
rect -18460 1901 -18444 1935
rect -18506 1860 -18444 1901
rect -18414 2819 -18348 2860
rect -18414 2785 -18398 2819
rect -18364 2785 -18348 2819
rect -18414 2751 -18348 2785
rect -18414 2717 -18398 2751
rect -18364 2717 -18348 2751
rect -18414 2683 -18348 2717
rect -18414 2649 -18398 2683
rect -18364 2649 -18348 2683
rect -18414 2615 -18348 2649
rect -18414 2581 -18398 2615
rect -18364 2581 -18348 2615
rect -18414 2547 -18348 2581
rect -18414 2513 -18398 2547
rect -18364 2513 -18348 2547
rect -18414 2479 -18348 2513
rect -18414 2445 -18398 2479
rect -18364 2445 -18348 2479
rect -18414 2411 -18348 2445
rect -18414 2377 -18398 2411
rect -18364 2377 -18348 2411
rect -18414 2343 -18348 2377
rect -18414 2309 -18398 2343
rect -18364 2309 -18348 2343
rect -18414 2275 -18348 2309
rect -18414 2241 -18398 2275
rect -18364 2241 -18348 2275
rect -18414 2207 -18348 2241
rect -18414 2173 -18398 2207
rect -18364 2173 -18348 2207
rect -18414 2139 -18348 2173
rect -18414 2105 -18398 2139
rect -18364 2105 -18348 2139
rect -18414 2071 -18348 2105
rect -18414 2037 -18398 2071
rect -18364 2037 -18348 2071
rect -18414 2003 -18348 2037
rect -18414 1969 -18398 2003
rect -18364 1969 -18348 2003
rect -18414 1935 -18348 1969
rect -18414 1901 -18398 1935
rect -18364 1901 -18348 1935
rect -18414 1860 -18348 1901
rect -18318 2819 -18252 2860
rect -18318 2785 -18302 2819
rect -18268 2785 -18252 2819
rect -18318 2751 -18252 2785
rect -18318 2717 -18302 2751
rect -18268 2717 -18252 2751
rect -18318 2683 -18252 2717
rect -18318 2649 -18302 2683
rect -18268 2649 -18252 2683
rect -18318 2615 -18252 2649
rect -18318 2581 -18302 2615
rect -18268 2581 -18252 2615
rect -18318 2547 -18252 2581
rect -18318 2513 -18302 2547
rect -18268 2513 -18252 2547
rect -18318 2479 -18252 2513
rect -18318 2445 -18302 2479
rect -18268 2445 -18252 2479
rect -18318 2411 -18252 2445
rect -18318 2377 -18302 2411
rect -18268 2377 -18252 2411
rect -18318 2343 -18252 2377
rect -18318 2309 -18302 2343
rect -18268 2309 -18252 2343
rect -18318 2275 -18252 2309
rect -18318 2241 -18302 2275
rect -18268 2241 -18252 2275
rect -18318 2207 -18252 2241
rect -18318 2173 -18302 2207
rect -18268 2173 -18252 2207
rect -18318 2139 -18252 2173
rect -18318 2105 -18302 2139
rect -18268 2105 -18252 2139
rect -18318 2071 -18252 2105
rect -18318 2037 -18302 2071
rect -18268 2037 -18252 2071
rect -18318 2003 -18252 2037
rect -18318 1969 -18302 2003
rect -18268 1969 -18252 2003
rect -18318 1935 -18252 1969
rect -18318 1901 -18302 1935
rect -18268 1901 -18252 1935
rect -18318 1860 -18252 1901
rect -18222 2819 -18156 2860
rect -18222 2785 -18206 2819
rect -18172 2785 -18156 2819
rect -18222 2751 -18156 2785
rect -18222 2717 -18206 2751
rect -18172 2717 -18156 2751
rect -18222 2683 -18156 2717
rect -18222 2649 -18206 2683
rect -18172 2649 -18156 2683
rect -18222 2615 -18156 2649
rect -18222 2581 -18206 2615
rect -18172 2581 -18156 2615
rect -18222 2547 -18156 2581
rect -18222 2513 -18206 2547
rect -18172 2513 -18156 2547
rect -18222 2479 -18156 2513
rect -18222 2445 -18206 2479
rect -18172 2445 -18156 2479
rect -18222 2411 -18156 2445
rect -18222 2377 -18206 2411
rect -18172 2377 -18156 2411
rect -18222 2343 -18156 2377
rect -18222 2309 -18206 2343
rect -18172 2309 -18156 2343
rect -18222 2275 -18156 2309
rect -18222 2241 -18206 2275
rect -18172 2241 -18156 2275
rect -18222 2207 -18156 2241
rect -18222 2173 -18206 2207
rect -18172 2173 -18156 2207
rect -18222 2139 -18156 2173
rect -18222 2105 -18206 2139
rect -18172 2105 -18156 2139
rect -18222 2071 -18156 2105
rect -18222 2037 -18206 2071
rect -18172 2037 -18156 2071
rect -18222 2003 -18156 2037
rect -18222 1969 -18206 2003
rect -18172 1969 -18156 2003
rect -18222 1935 -18156 1969
rect -18222 1901 -18206 1935
rect -18172 1901 -18156 1935
rect -18222 1860 -18156 1901
rect -18126 2819 -18060 2860
rect -18126 2785 -18110 2819
rect -18076 2785 -18060 2819
rect -18126 2751 -18060 2785
rect -18126 2717 -18110 2751
rect -18076 2717 -18060 2751
rect -18126 2683 -18060 2717
rect -18126 2649 -18110 2683
rect -18076 2649 -18060 2683
rect -18126 2615 -18060 2649
rect -18126 2581 -18110 2615
rect -18076 2581 -18060 2615
rect -18126 2547 -18060 2581
rect -18126 2513 -18110 2547
rect -18076 2513 -18060 2547
rect -18126 2479 -18060 2513
rect -18126 2445 -18110 2479
rect -18076 2445 -18060 2479
rect -18126 2411 -18060 2445
rect -18126 2377 -18110 2411
rect -18076 2377 -18060 2411
rect -18126 2343 -18060 2377
rect -18126 2309 -18110 2343
rect -18076 2309 -18060 2343
rect -18126 2275 -18060 2309
rect -18126 2241 -18110 2275
rect -18076 2241 -18060 2275
rect -18126 2207 -18060 2241
rect -18126 2173 -18110 2207
rect -18076 2173 -18060 2207
rect -18126 2139 -18060 2173
rect -18126 2105 -18110 2139
rect -18076 2105 -18060 2139
rect -18126 2071 -18060 2105
rect -18126 2037 -18110 2071
rect -18076 2037 -18060 2071
rect -18126 2003 -18060 2037
rect -18126 1969 -18110 2003
rect -18076 1969 -18060 2003
rect -18126 1935 -18060 1969
rect -18126 1901 -18110 1935
rect -18076 1901 -18060 1935
rect -18126 1860 -18060 1901
rect -18030 2819 -17968 2860
rect -18030 2785 -18014 2819
rect -17980 2785 -17968 2819
rect -18030 2751 -17968 2785
rect -18030 2717 -18014 2751
rect -17980 2717 -17968 2751
rect -18030 2683 -17968 2717
rect -18030 2649 -18014 2683
rect -17980 2649 -17968 2683
rect -18030 2615 -17968 2649
rect -18030 2581 -18014 2615
rect -17980 2581 -17968 2615
rect -18030 2547 -17968 2581
rect -18030 2513 -18014 2547
rect -17980 2513 -17968 2547
rect -18030 2479 -17968 2513
rect -18030 2445 -18014 2479
rect -17980 2445 -17968 2479
rect -18030 2411 -17968 2445
rect -18030 2377 -18014 2411
rect -17980 2377 -17968 2411
rect -18030 2343 -17968 2377
rect -18030 2309 -18014 2343
rect -17980 2309 -17968 2343
rect -18030 2275 -17968 2309
rect -18030 2241 -18014 2275
rect -17980 2241 -17968 2275
rect -18030 2207 -17968 2241
rect -18030 2173 -18014 2207
rect -17980 2173 -17968 2207
rect -18030 2139 -17968 2173
rect -18030 2105 -18014 2139
rect -17980 2105 -17968 2139
rect -18030 2071 -17968 2105
rect -18030 2037 -18014 2071
rect -17980 2037 -17968 2071
rect -18030 2003 -17968 2037
rect -18030 1969 -18014 2003
rect -17980 1969 -17968 2003
rect -18030 1935 -17968 1969
rect -18030 1901 -18014 1935
rect -17980 1901 -17968 1935
rect -18030 1860 -17968 1901
rect -16674 2825 -16612 2866
rect -16674 2791 -16662 2825
rect -16628 2791 -16612 2825
rect -16674 2757 -16612 2791
rect -16674 2723 -16662 2757
rect -16628 2723 -16612 2757
rect -16674 2689 -16612 2723
rect -16674 2655 -16662 2689
rect -16628 2655 -16612 2689
rect -16674 2621 -16612 2655
rect -16674 2587 -16662 2621
rect -16628 2587 -16612 2621
rect -16674 2553 -16612 2587
rect -16674 2519 -16662 2553
rect -16628 2519 -16612 2553
rect -16674 2485 -16612 2519
rect -16674 2451 -16662 2485
rect -16628 2451 -16612 2485
rect -16674 2417 -16612 2451
rect -16674 2383 -16662 2417
rect -16628 2383 -16612 2417
rect -16674 2349 -16612 2383
rect -16674 2315 -16662 2349
rect -16628 2315 -16612 2349
rect -16674 2281 -16612 2315
rect -16674 2247 -16662 2281
rect -16628 2247 -16612 2281
rect -16674 2213 -16612 2247
rect -16674 2179 -16662 2213
rect -16628 2179 -16612 2213
rect -16674 2145 -16612 2179
rect -16674 2111 -16662 2145
rect -16628 2111 -16612 2145
rect -16674 2077 -16612 2111
rect -16674 2043 -16662 2077
rect -16628 2043 -16612 2077
rect -16674 2009 -16612 2043
rect -16674 1975 -16662 2009
rect -16628 1975 -16612 2009
rect -16674 1941 -16612 1975
rect -16674 1907 -16662 1941
rect -16628 1907 -16612 1941
rect -16674 1866 -16612 1907
rect -16582 2825 -16516 2866
rect -16582 2791 -16566 2825
rect -16532 2791 -16516 2825
rect -16582 2757 -16516 2791
rect -16582 2723 -16566 2757
rect -16532 2723 -16516 2757
rect -16582 2689 -16516 2723
rect -16582 2655 -16566 2689
rect -16532 2655 -16516 2689
rect -16582 2621 -16516 2655
rect -16582 2587 -16566 2621
rect -16532 2587 -16516 2621
rect -16582 2553 -16516 2587
rect -16582 2519 -16566 2553
rect -16532 2519 -16516 2553
rect -16582 2485 -16516 2519
rect -16582 2451 -16566 2485
rect -16532 2451 -16516 2485
rect -16582 2417 -16516 2451
rect -16582 2383 -16566 2417
rect -16532 2383 -16516 2417
rect -16582 2349 -16516 2383
rect -16582 2315 -16566 2349
rect -16532 2315 -16516 2349
rect -16582 2281 -16516 2315
rect -16582 2247 -16566 2281
rect -16532 2247 -16516 2281
rect -16582 2213 -16516 2247
rect -16582 2179 -16566 2213
rect -16532 2179 -16516 2213
rect -16582 2145 -16516 2179
rect -16582 2111 -16566 2145
rect -16532 2111 -16516 2145
rect -16582 2077 -16516 2111
rect -16582 2043 -16566 2077
rect -16532 2043 -16516 2077
rect -16582 2009 -16516 2043
rect -16582 1975 -16566 2009
rect -16532 1975 -16516 2009
rect -16582 1941 -16516 1975
rect -16582 1907 -16566 1941
rect -16532 1907 -16516 1941
rect -16582 1866 -16516 1907
rect -16486 2825 -16420 2866
rect -16486 2791 -16470 2825
rect -16436 2791 -16420 2825
rect -16486 2757 -16420 2791
rect -16486 2723 -16470 2757
rect -16436 2723 -16420 2757
rect -16486 2689 -16420 2723
rect -16486 2655 -16470 2689
rect -16436 2655 -16420 2689
rect -16486 2621 -16420 2655
rect -16486 2587 -16470 2621
rect -16436 2587 -16420 2621
rect -16486 2553 -16420 2587
rect -16486 2519 -16470 2553
rect -16436 2519 -16420 2553
rect -16486 2485 -16420 2519
rect -16486 2451 -16470 2485
rect -16436 2451 -16420 2485
rect -16486 2417 -16420 2451
rect -16486 2383 -16470 2417
rect -16436 2383 -16420 2417
rect -16486 2349 -16420 2383
rect -16486 2315 -16470 2349
rect -16436 2315 -16420 2349
rect -16486 2281 -16420 2315
rect -16486 2247 -16470 2281
rect -16436 2247 -16420 2281
rect -16486 2213 -16420 2247
rect -16486 2179 -16470 2213
rect -16436 2179 -16420 2213
rect -16486 2145 -16420 2179
rect -16486 2111 -16470 2145
rect -16436 2111 -16420 2145
rect -16486 2077 -16420 2111
rect -16486 2043 -16470 2077
rect -16436 2043 -16420 2077
rect -16486 2009 -16420 2043
rect -16486 1975 -16470 2009
rect -16436 1975 -16420 2009
rect -16486 1941 -16420 1975
rect -16486 1907 -16470 1941
rect -16436 1907 -16420 1941
rect -16486 1866 -16420 1907
rect -16390 2825 -16324 2866
rect -16390 2791 -16374 2825
rect -16340 2791 -16324 2825
rect -16390 2757 -16324 2791
rect -16390 2723 -16374 2757
rect -16340 2723 -16324 2757
rect -16390 2689 -16324 2723
rect -16390 2655 -16374 2689
rect -16340 2655 -16324 2689
rect -16390 2621 -16324 2655
rect -16390 2587 -16374 2621
rect -16340 2587 -16324 2621
rect -16390 2553 -16324 2587
rect -16390 2519 -16374 2553
rect -16340 2519 -16324 2553
rect -16390 2485 -16324 2519
rect -16390 2451 -16374 2485
rect -16340 2451 -16324 2485
rect -16390 2417 -16324 2451
rect -16390 2383 -16374 2417
rect -16340 2383 -16324 2417
rect -16390 2349 -16324 2383
rect -16390 2315 -16374 2349
rect -16340 2315 -16324 2349
rect -16390 2281 -16324 2315
rect -16390 2247 -16374 2281
rect -16340 2247 -16324 2281
rect -16390 2213 -16324 2247
rect -16390 2179 -16374 2213
rect -16340 2179 -16324 2213
rect -16390 2145 -16324 2179
rect -16390 2111 -16374 2145
rect -16340 2111 -16324 2145
rect -16390 2077 -16324 2111
rect -16390 2043 -16374 2077
rect -16340 2043 -16324 2077
rect -16390 2009 -16324 2043
rect -16390 1975 -16374 2009
rect -16340 1975 -16324 2009
rect -16390 1941 -16324 1975
rect -16390 1907 -16374 1941
rect -16340 1907 -16324 1941
rect -16390 1866 -16324 1907
rect -16294 2825 -16228 2866
rect -16294 2791 -16278 2825
rect -16244 2791 -16228 2825
rect -16294 2757 -16228 2791
rect -16294 2723 -16278 2757
rect -16244 2723 -16228 2757
rect -16294 2689 -16228 2723
rect -16294 2655 -16278 2689
rect -16244 2655 -16228 2689
rect -16294 2621 -16228 2655
rect -16294 2587 -16278 2621
rect -16244 2587 -16228 2621
rect -16294 2553 -16228 2587
rect -16294 2519 -16278 2553
rect -16244 2519 -16228 2553
rect -16294 2485 -16228 2519
rect -16294 2451 -16278 2485
rect -16244 2451 -16228 2485
rect -16294 2417 -16228 2451
rect -16294 2383 -16278 2417
rect -16244 2383 -16228 2417
rect -16294 2349 -16228 2383
rect -16294 2315 -16278 2349
rect -16244 2315 -16228 2349
rect -16294 2281 -16228 2315
rect -16294 2247 -16278 2281
rect -16244 2247 -16228 2281
rect -16294 2213 -16228 2247
rect -16294 2179 -16278 2213
rect -16244 2179 -16228 2213
rect -16294 2145 -16228 2179
rect -16294 2111 -16278 2145
rect -16244 2111 -16228 2145
rect -16294 2077 -16228 2111
rect -16294 2043 -16278 2077
rect -16244 2043 -16228 2077
rect -16294 2009 -16228 2043
rect -16294 1975 -16278 2009
rect -16244 1975 -16228 2009
rect -16294 1941 -16228 1975
rect -16294 1907 -16278 1941
rect -16244 1907 -16228 1941
rect -16294 1866 -16228 1907
rect -16198 2825 -16132 2866
rect -16198 2791 -16182 2825
rect -16148 2791 -16132 2825
rect -16198 2757 -16132 2791
rect -16198 2723 -16182 2757
rect -16148 2723 -16132 2757
rect -16198 2689 -16132 2723
rect -16198 2655 -16182 2689
rect -16148 2655 -16132 2689
rect -16198 2621 -16132 2655
rect -16198 2587 -16182 2621
rect -16148 2587 -16132 2621
rect -16198 2553 -16132 2587
rect -16198 2519 -16182 2553
rect -16148 2519 -16132 2553
rect -16198 2485 -16132 2519
rect -16198 2451 -16182 2485
rect -16148 2451 -16132 2485
rect -16198 2417 -16132 2451
rect -16198 2383 -16182 2417
rect -16148 2383 -16132 2417
rect -16198 2349 -16132 2383
rect -16198 2315 -16182 2349
rect -16148 2315 -16132 2349
rect -16198 2281 -16132 2315
rect -16198 2247 -16182 2281
rect -16148 2247 -16132 2281
rect -16198 2213 -16132 2247
rect -16198 2179 -16182 2213
rect -16148 2179 -16132 2213
rect -16198 2145 -16132 2179
rect -16198 2111 -16182 2145
rect -16148 2111 -16132 2145
rect -16198 2077 -16132 2111
rect -16198 2043 -16182 2077
rect -16148 2043 -16132 2077
rect -16198 2009 -16132 2043
rect -16198 1975 -16182 2009
rect -16148 1975 -16132 2009
rect -16198 1941 -16132 1975
rect -16198 1907 -16182 1941
rect -16148 1907 -16132 1941
rect -16198 1866 -16132 1907
rect -16102 2825 -16036 2866
rect -16102 2791 -16086 2825
rect -16052 2791 -16036 2825
rect -16102 2757 -16036 2791
rect -16102 2723 -16086 2757
rect -16052 2723 -16036 2757
rect -16102 2689 -16036 2723
rect -16102 2655 -16086 2689
rect -16052 2655 -16036 2689
rect -16102 2621 -16036 2655
rect -16102 2587 -16086 2621
rect -16052 2587 -16036 2621
rect -16102 2553 -16036 2587
rect -16102 2519 -16086 2553
rect -16052 2519 -16036 2553
rect -16102 2485 -16036 2519
rect -16102 2451 -16086 2485
rect -16052 2451 -16036 2485
rect -16102 2417 -16036 2451
rect -16102 2383 -16086 2417
rect -16052 2383 -16036 2417
rect -16102 2349 -16036 2383
rect -16102 2315 -16086 2349
rect -16052 2315 -16036 2349
rect -16102 2281 -16036 2315
rect -16102 2247 -16086 2281
rect -16052 2247 -16036 2281
rect -16102 2213 -16036 2247
rect -16102 2179 -16086 2213
rect -16052 2179 -16036 2213
rect -16102 2145 -16036 2179
rect -16102 2111 -16086 2145
rect -16052 2111 -16036 2145
rect -16102 2077 -16036 2111
rect -16102 2043 -16086 2077
rect -16052 2043 -16036 2077
rect -16102 2009 -16036 2043
rect -16102 1975 -16086 2009
rect -16052 1975 -16036 2009
rect -16102 1941 -16036 1975
rect -16102 1907 -16086 1941
rect -16052 1907 -16036 1941
rect -16102 1866 -16036 1907
rect -16006 2825 -15940 2866
rect -16006 2791 -15990 2825
rect -15956 2791 -15940 2825
rect -16006 2757 -15940 2791
rect -16006 2723 -15990 2757
rect -15956 2723 -15940 2757
rect -16006 2689 -15940 2723
rect -16006 2655 -15990 2689
rect -15956 2655 -15940 2689
rect -16006 2621 -15940 2655
rect -16006 2587 -15990 2621
rect -15956 2587 -15940 2621
rect -16006 2553 -15940 2587
rect -16006 2519 -15990 2553
rect -15956 2519 -15940 2553
rect -16006 2485 -15940 2519
rect -16006 2451 -15990 2485
rect -15956 2451 -15940 2485
rect -16006 2417 -15940 2451
rect -16006 2383 -15990 2417
rect -15956 2383 -15940 2417
rect -16006 2349 -15940 2383
rect -16006 2315 -15990 2349
rect -15956 2315 -15940 2349
rect -16006 2281 -15940 2315
rect -16006 2247 -15990 2281
rect -15956 2247 -15940 2281
rect -16006 2213 -15940 2247
rect -16006 2179 -15990 2213
rect -15956 2179 -15940 2213
rect -16006 2145 -15940 2179
rect -16006 2111 -15990 2145
rect -15956 2111 -15940 2145
rect -16006 2077 -15940 2111
rect -16006 2043 -15990 2077
rect -15956 2043 -15940 2077
rect -16006 2009 -15940 2043
rect -16006 1975 -15990 2009
rect -15956 1975 -15940 2009
rect -16006 1941 -15940 1975
rect -16006 1907 -15990 1941
rect -15956 1907 -15940 1941
rect -16006 1866 -15940 1907
rect -15910 2825 -15844 2866
rect -15910 2791 -15894 2825
rect -15860 2791 -15844 2825
rect -15910 2757 -15844 2791
rect -15910 2723 -15894 2757
rect -15860 2723 -15844 2757
rect -15910 2689 -15844 2723
rect -15910 2655 -15894 2689
rect -15860 2655 -15844 2689
rect -15910 2621 -15844 2655
rect -15910 2587 -15894 2621
rect -15860 2587 -15844 2621
rect -15910 2553 -15844 2587
rect -15910 2519 -15894 2553
rect -15860 2519 -15844 2553
rect -15910 2485 -15844 2519
rect -15910 2451 -15894 2485
rect -15860 2451 -15844 2485
rect -15910 2417 -15844 2451
rect -15910 2383 -15894 2417
rect -15860 2383 -15844 2417
rect -15910 2349 -15844 2383
rect -15910 2315 -15894 2349
rect -15860 2315 -15844 2349
rect -15910 2281 -15844 2315
rect -15910 2247 -15894 2281
rect -15860 2247 -15844 2281
rect -15910 2213 -15844 2247
rect -15910 2179 -15894 2213
rect -15860 2179 -15844 2213
rect -15910 2145 -15844 2179
rect -15910 2111 -15894 2145
rect -15860 2111 -15844 2145
rect -15910 2077 -15844 2111
rect -15910 2043 -15894 2077
rect -15860 2043 -15844 2077
rect -15910 2009 -15844 2043
rect -15910 1975 -15894 2009
rect -15860 1975 -15844 2009
rect -15910 1941 -15844 1975
rect -15910 1907 -15894 1941
rect -15860 1907 -15844 1941
rect -15910 1866 -15844 1907
rect -15814 2825 -15748 2866
rect -15814 2791 -15798 2825
rect -15764 2791 -15748 2825
rect -15814 2757 -15748 2791
rect -15814 2723 -15798 2757
rect -15764 2723 -15748 2757
rect -15814 2689 -15748 2723
rect -15814 2655 -15798 2689
rect -15764 2655 -15748 2689
rect -15814 2621 -15748 2655
rect -15814 2587 -15798 2621
rect -15764 2587 -15748 2621
rect -15814 2553 -15748 2587
rect -15814 2519 -15798 2553
rect -15764 2519 -15748 2553
rect -15814 2485 -15748 2519
rect -15814 2451 -15798 2485
rect -15764 2451 -15748 2485
rect -15814 2417 -15748 2451
rect -15814 2383 -15798 2417
rect -15764 2383 -15748 2417
rect -15814 2349 -15748 2383
rect -15814 2315 -15798 2349
rect -15764 2315 -15748 2349
rect -15814 2281 -15748 2315
rect -15814 2247 -15798 2281
rect -15764 2247 -15748 2281
rect -15814 2213 -15748 2247
rect -15814 2179 -15798 2213
rect -15764 2179 -15748 2213
rect -15814 2145 -15748 2179
rect -15814 2111 -15798 2145
rect -15764 2111 -15748 2145
rect -15814 2077 -15748 2111
rect -15814 2043 -15798 2077
rect -15764 2043 -15748 2077
rect -15814 2009 -15748 2043
rect -15814 1975 -15798 2009
rect -15764 1975 -15748 2009
rect -15814 1941 -15748 1975
rect -15814 1907 -15798 1941
rect -15764 1907 -15748 1941
rect -15814 1866 -15748 1907
rect -15718 2825 -15652 2866
rect -15718 2791 -15702 2825
rect -15668 2791 -15652 2825
rect -15718 2757 -15652 2791
rect -15718 2723 -15702 2757
rect -15668 2723 -15652 2757
rect -15718 2689 -15652 2723
rect -15718 2655 -15702 2689
rect -15668 2655 -15652 2689
rect -15718 2621 -15652 2655
rect -15718 2587 -15702 2621
rect -15668 2587 -15652 2621
rect -15718 2553 -15652 2587
rect -15718 2519 -15702 2553
rect -15668 2519 -15652 2553
rect -15718 2485 -15652 2519
rect -15718 2451 -15702 2485
rect -15668 2451 -15652 2485
rect -15718 2417 -15652 2451
rect -15718 2383 -15702 2417
rect -15668 2383 -15652 2417
rect -15718 2349 -15652 2383
rect -15718 2315 -15702 2349
rect -15668 2315 -15652 2349
rect -15718 2281 -15652 2315
rect -15718 2247 -15702 2281
rect -15668 2247 -15652 2281
rect -15718 2213 -15652 2247
rect -15718 2179 -15702 2213
rect -15668 2179 -15652 2213
rect -15718 2145 -15652 2179
rect -15718 2111 -15702 2145
rect -15668 2111 -15652 2145
rect -15718 2077 -15652 2111
rect -15718 2043 -15702 2077
rect -15668 2043 -15652 2077
rect -15718 2009 -15652 2043
rect -15718 1975 -15702 2009
rect -15668 1975 -15652 2009
rect -15718 1941 -15652 1975
rect -15718 1907 -15702 1941
rect -15668 1907 -15652 1941
rect -15718 1866 -15652 1907
rect -15622 2825 -15556 2866
rect -15622 2791 -15606 2825
rect -15572 2791 -15556 2825
rect -15622 2757 -15556 2791
rect -15622 2723 -15606 2757
rect -15572 2723 -15556 2757
rect -15622 2689 -15556 2723
rect -15622 2655 -15606 2689
rect -15572 2655 -15556 2689
rect -15622 2621 -15556 2655
rect -15622 2587 -15606 2621
rect -15572 2587 -15556 2621
rect -15622 2553 -15556 2587
rect -15622 2519 -15606 2553
rect -15572 2519 -15556 2553
rect -15622 2485 -15556 2519
rect -15622 2451 -15606 2485
rect -15572 2451 -15556 2485
rect -15622 2417 -15556 2451
rect -15622 2383 -15606 2417
rect -15572 2383 -15556 2417
rect -15622 2349 -15556 2383
rect -15622 2315 -15606 2349
rect -15572 2315 -15556 2349
rect -15622 2281 -15556 2315
rect -15622 2247 -15606 2281
rect -15572 2247 -15556 2281
rect -15622 2213 -15556 2247
rect -15622 2179 -15606 2213
rect -15572 2179 -15556 2213
rect -15622 2145 -15556 2179
rect -15622 2111 -15606 2145
rect -15572 2111 -15556 2145
rect -15622 2077 -15556 2111
rect -15622 2043 -15606 2077
rect -15572 2043 -15556 2077
rect -15622 2009 -15556 2043
rect -15622 1975 -15606 2009
rect -15572 1975 -15556 2009
rect -15622 1941 -15556 1975
rect -15622 1907 -15606 1941
rect -15572 1907 -15556 1941
rect -15622 1866 -15556 1907
rect -15526 2825 -15460 2866
rect -15526 2791 -15510 2825
rect -15476 2791 -15460 2825
rect -15526 2757 -15460 2791
rect -15526 2723 -15510 2757
rect -15476 2723 -15460 2757
rect -15526 2689 -15460 2723
rect -15526 2655 -15510 2689
rect -15476 2655 -15460 2689
rect -15526 2621 -15460 2655
rect -15526 2587 -15510 2621
rect -15476 2587 -15460 2621
rect -15526 2553 -15460 2587
rect -15526 2519 -15510 2553
rect -15476 2519 -15460 2553
rect -15526 2485 -15460 2519
rect -15526 2451 -15510 2485
rect -15476 2451 -15460 2485
rect -15526 2417 -15460 2451
rect -15526 2383 -15510 2417
rect -15476 2383 -15460 2417
rect -15526 2349 -15460 2383
rect -15526 2315 -15510 2349
rect -15476 2315 -15460 2349
rect -15526 2281 -15460 2315
rect -15526 2247 -15510 2281
rect -15476 2247 -15460 2281
rect -15526 2213 -15460 2247
rect -15526 2179 -15510 2213
rect -15476 2179 -15460 2213
rect -15526 2145 -15460 2179
rect -15526 2111 -15510 2145
rect -15476 2111 -15460 2145
rect -15526 2077 -15460 2111
rect -15526 2043 -15510 2077
rect -15476 2043 -15460 2077
rect -15526 2009 -15460 2043
rect -15526 1975 -15510 2009
rect -15476 1975 -15460 2009
rect -15526 1941 -15460 1975
rect -15526 1907 -15510 1941
rect -15476 1907 -15460 1941
rect -15526 1866 -15460 1907
rect -15430 2825 -15364 2866
rect -15430 2791 -15414 2825
rect -15380 2791 -15364 2825
rect -15430 2757 -15364 2791
rect -15430 2723 -15414 2757
rect -15380 2723 -15364 2757
rect -15430 2689 -15364 2723
rect -15430 2655 -15414 2689
rect -15380 2655 -15364 2689
rect -15430 2621 -15364 2655
rect -15430 2587 -15414 2621
rect -15380 2587 -15364 2621
rect -15430 2553 -15364 2587
rect -15430 2519 -15414 2553
rect -15380 2519 -15364 2553
rect -15430 2485 -15364 2519
rect -15430 2451 -15414 2485
rect -15380 2451 -15364 2485
rect -15430 2417 -15364 2451
rect -15430 2383 -15414 2417
rect -15380 2383 -15364 2417
rect -15430 2349 -15364 2383
rect -15430 2315 -15414 2349
rect -15380 2315 -15364 2349
rect -15430 2281 -15364 2315
rect -15430 2247 -15414 2281
rect -15380 2247 -15364 2281
rect -15430 2213 -15364 2247
rect -15430 2179 -15414 2213
rect -15380 2179 -15364 2213
rect -15430 2145 -15364 2179
rect -15430 2111 -15414 2145
rect -15380 2111 -15364 2145
rect -15430 2077 -15364 2111
rect -15430 2043 -15414 2077
rect -15380 2043 -15364 2077
rect -15430 2009 -15364 2043
rect -15430 1975 -15414 2009
rect -15380 1975 -15364 2009
rect -15430 1941 -15364 1975
rect -15430 1907 -15414 1941
rect -15380 1907 -15364 1941
rect -15430 1866 -15364 1907
rect -15334 2825 -15268 2866
rect -15334 2791 -15318 2825
rect -15284 2791 -15268 2825
rect -15334 2757 -15268 2791
rect -15334 2723 -15318 2757
rect -15284 2723 -15268 2757
rect -15334 2689 -15268 2723
rect -15334 2655 -15318 2689
rect -15284 2655 -15268 2689
rect -15334 2621 -15268 2655
rect -15334 2587 -15318 2621
rect -15284 2587 -15268 2621
rect -15334 2553 -15268 2587
rect -15334 2519 -15318 2553
rect -15284 2519 -15268 2553
rect -15334 2485 -15268 2519
rect -15334 2451 -15318 2485
rect -15284 2451 -15268 2485
rect -15334 2417 -15268 2451
rect -15334 2383 -15318 2417
rect -15284 2383 -15268 2417
rect -15334 2349 -15268 2383
rect -15334 2315 -15318 2349
rect -15284 2315 -15268 2349
rect -15334 2281 -15268 2315
rect -15334 2247 -15318 2281
rect -15284 2247 -15268 2281
rect -15334 2213 -15268 2247
rect -15334 2179 -15318 2213
rect -15284 2179 -15268 2213
rect -15334 2145 -15268 2179
rect -15334 2111 -15318 2145
rect -15284 2111 -15268 2145
rect -15334 2077 -15268 2111
rect -15334 2043 -15318 2077
rect -15284 2043 -15268 2077
rect -15334 2009 -15268 2043
rect -15334 1975 -15318 2009
rect -15284 1975 -15268 2009
rect -15334 1941 -15268 1975
rect -15334 1907 -15318 1941
rect -15284 1907 -15268 1941
rect -15334 1866 -15268 1907
rect -15238 2825 -15172 2866
rect -15238 2791 -15222 2825
rect -15188 2791 -15172 2825
rect -15238 2757 -15172 2791
rect -15238 2723 -15222 2757
rect -15188 2723 -15172 2757
rect -15238 2689 -15172 2723
rect -15238 2655 -15222 2689
rect -15188 2655 -15172 2689
rect -15238 2621 -15172 2655
rect -15238 2587 -15222 2621
rect -15188 2587 -15172 2621
rect -15238 2553 -15172 2587
rect -15238 2519 -15222 2553
rect -15188 2519 -15172 2553
rect -15238 2485 -15172 2519
rect -15238 2451 -15222 2485
rect -15188 2451 -15172 2485
rect -15238 2417 -15172 2451
rect -15238 2383 -15222 2417
rect -15188 2383 -15172 2417
rect -15238 2349 -15172 2383
rect -15238 2315 -15222 2349
rect -15188 2315 -15172 2349
rect -15238 2281 -15172 2315
rect -15238 2247 -15222 2281
rect -15188 2247 -15172 2281
rect -15238 2213 -15172 2247
rect -15238 2179 -15222 2213
rect -15188 2179 -15172 2213
rect -15238 2145 -15172 2179
rect -15238 2111 -15222 2145
rect -15188 2111 -15172 2145
rect -15238 2077 -15172 2111
rect -15238 2043 -15222 2077
rect -15188 2043 -15172 2077
rect -15238 2009 -15172 2043
rect -15238 1975 -15222 2009
rect -15188 1975 -15172 2009
rect -15238 1941 -15172 1975
rect -15238 1907 -15222 1941
rect -15188 1907 -15172 1941
rect -15238 1866 -15172 1907
rect -15142 2825 -15076 2866
rect -15142 2791 -15126 2825
rect -15092 2791 -15076 2825
rect -15142 2757 -15076 2791
rect -15142 2723 -15126 2757
rect -15092 2723 -15076 2757
rect -15142 2689 -15076 2723
rect -15142 2655 -15126 2689
rect -15092 2655 -15076 2689
rect -15142 2621 -15076 2655
rect -15142 2587 -15126 2621
rect -15092 2587 -15076 2621
rect -15142 2553 -15076 2587
rect -15142 2519 -15126 2553
rect -15092 2519 -15076 2553
rect -15142 2485 -15076 2519
rect -15142 2451 -15126 2485
rect -15092 2451 -15076 2485
rect -15142 2417 -15076 2451
rect -15142 2383 -15126 2417
rect -15092 2383 -15076 2417
rect -15142 2349 -15076 2383
rect -15142 2315 -15126 2349
rect -15092 2315 -15076 2349
rect -15142 2281 -15076 2315
rect -15142 2247 -15126 2281
rect -15092 2247 -15076 2281
rect -15142 2213 -15076 2247
rect -15142 2179 -15126 2213
rect -15092 2179 -15076 2213
rect -15142 2145 -15076 2179
rect -15142 2111 -15126 2145
rect -15092 2111 -15076 2145
rect -15142 2077 -15076 2111
rect -15142 2043 -15126 2077
rect -15092 2043 -15076 2077
rect -15142 2009 -15076 2043
rect -15142 1975 -15126 2009
rect -15092 1975 -15076 2009
rect -15142 1941 -15076 1975
rect -15142 1907 -15126 1941
rect -15092 1907 -15076 1941
rect -15142 1866 -15076 1907
rect -15046 2825 -14980 2866
rect -15046 2791 -15030 2825
rect -14996 2791 -14980 2825
rect -15046 2757 -14980 2791
rect -15046 2723 -15030 2757
rect -14996 2723 -14980 2757
rect -15046 2689 -14980 2723
rect -15046 2655 -15030 2689
rect -14996 2655 -14980 2689
rect -15046 2621 -14980 2655
rect -15046 2587 -15030 2621
rect -14996 2587 -14980 2621
rect -15046 2553 -14980 2587
rect -15046 2519 -15030 2553
rect -14996 2519 -14980 2553
rect -15046 2485 -14980 2519
rect -15046 2451 -15030 2485
rect -14996 2451 -14980 2485
rect -15046 2417 -14980 2451
rect -15046 2383 -15030 2417
rect -14996 2383 -14980 2417
rect -15046 2349 -14980 2383
rect -15046 2315 -15030 2349
rect -14996 2315 -14980 2349
rect -15046 2281 -14980 2315
rect -15046 2247 -15030 2281
rect -14996 2247 -14980 2281
rect -15046 2213 -14980 2247
rect -15046 2179 -15030 2213
rect -14996 2179 -14980 2213
rect -15046 2145 -14980 2179
rect -15046 2111 -15030 2145
rect -14996 2111 -14980 2145
rect -15046 2077 -14980 2111
rect -15046 2043 -15030 2077
rect -14996 2043 -14980 2077
rect -15046 2009 -14980 2043
rect -15046 1975 -15030 2009
rect -14996 1975 -14980 2009
rect -15046 1941 -14980 1975
rect -15046 1907 -15030 1941
rect -14996 1907 -14980 1941
rect -15046 1866 -14980 1907
rect -14950 2825 -14884 2866
rect -14950 2791 -14934 2825
rect -14900 2791 -14884 2825
rect -14950 2757 -14884 2791
rect -14950 2723 -14934 2757
rect -14900 2723 -14884 2757
rect -14950 2689 -14884 2723
rect -14950 2655 -14934 2689
rect -14900 2655 -14884 2689
rect -14950 2621 -14884 2655
rect -14950 2587 -14934 2621
rect -14900 2587 -14884 2621
rect -14950 2553 -14884 2587
rect -14950 2519 -14934 2553
rect -14900 2519 -14884 2553
rect -14950 2485 -14884 2519
rect -14950 2451 -14934 2485
rect -14900 2451 -14884 2485
rect -14950 2417 -14884 2451
rect -14950 2383 -14934 2417
rect -14900 2383 -14884 2417
rect -14950 2349 -14884 2383
rect -14950 2315 -14934 2349
rect -14900 2315 -14884 2349
rect -14950 2281 -14884 2315
rect -14950 2247 -14934 2281
rect -14900 2247 -14884 2281
rect -14950 2213 -14884 2247
rect -14950 2179 -14934 2213
rect -14900 2179 -14884 2213
rect -14950 2145 -14884 2179
rect -14950 2111 -14934 2145
rect -14900 2111 -14884 2145
rect -14950 2077 -14884 2111
rect -14950 2043 -14934 2077
rect -14900 2043 -14884 2077
rect -14950 2009 -14884 2043
rect -14950 1975 -14934 2009
rect -14900 1975 -14884 2009
rect -14950 1941 -14884 1975
rect -14950 1907 -14934 1941
rect -14900 1907 -14884 1941
rect -14950 1866 -14884 1907
rect -14854 2825 -14788 2866
rect -14854 2791 -14838 2825
rect -14804 2791 -14788 2825
rect -14854 2757 -14788 2791
rect -14854 2723 -14838 2757
rect -14804 2723 -14788 2757
rect -14854 2689 -14788 2723
rect -14854 2655 -14838 2689
rect -14804 2655 -14788 2689
rect -14854 2621 -14788 2655
rect -14854 2587 -14838 2621
rect -14804 2587 -14788 2621
rect -14854 2553 -14788 2587
rect -14854 2519 -14838 2553
rect -14804 2519 -14788 2553
rect -14854 2485 -14788 2519
rect -14854 2451 -14838 2485
rect -14804 2451 -14788 2485
rect -14854 2417 -14788 2451
rect -14854 2383 -14838 2417
rect -14804 2383 -14788 2417
rect -14854 2349 -14788 2383
rect -14854 2315 -14838 2349
rect -14804 2315 -14788 2349
rect -14854 2281 -14788 2315
rect -14854 2247 -14838 2281
rect -14804 2247 -14788 2281
rect -14854 2213 -14788 2247
rect -14854 2179 -14838 2213
rect -14804 2179 -14788 2213
rect -14854 2145 -14788 2179
rect -14854 2111 -14838 2145
rect -14804 2111 -14788 2145
rect -14854 2077 -14788 2111
rect -14854 2043 -14838 2077
rect -14804 2043 -14788 2077
rect -14854 2009 -14788 2043
rect -14854 1975 -14838 2009
rect -14804 1975 -14788 2009
rect -14854 1941 -14788 1975
rect -14854 1907 -14838 1941
rect -14804 1907 -14788 1941
rect -14854 1866 -14788 1907
rect -14758 2825 -14696 2866
rect -1698 3025 -1686 3059
rect -1652 3025 -1636 3059
rect -1698 2991 -1636 3025
rect -1698 2957 -1686 2991
rect -1652 2957 -1636 2991
rect -1698 2923 -1636 2957
rect -14758 2791 -14742 2825
rect -14708 2791 -14696 2825
rect -14758 2757 -14696 2791
rect -14758 2723 -14742 2757
rect -14708 2723 -14696 2757
rect -14758 2689 -14696 2723
rect -14758 2655 -14742 2689
rect -14708 2655 -14696 2689
rect -14758 2621 -14696 2655
rect -14758 2587 -14742 2621
rect -14708 2587 -14696 2621
rect -14758 2553 -14696 2587
rect -14758 2519 -14742 2553
rect -14708 2519 -14696 2553
rect -14758 2485 -14696 2519
rect -14758 2451 -14742 2485
rect -14708 2451 -14696 2485
rect -14758 2417 -14696 2451
rect -14758 2383 -14742 2417
rect -14708 2383 -14696 2417
rect -14758 2349 -14696 2383
rect -14758 2315 -14742 2349
rect -14708 2315 -14696 2349
rect -14758 2281 -14696 2315
rect -14758 2247 -14742 2281
rect -14708 2247 -14696 2281
rect -14758 2213 -14696 2247
rect -14758 2179 -14742 2213
rect -14708 2179 -14696 2213
rect -14758 2145 -14696 2179
rect -14758 2111 -14742 2145
rect -14708 2111 -14696 2145
rect -14758 2077 -14696 2111
rect -14758 2043 -14742 2077
rect -14708 2043 -14696 2077
rect -14758 2009 -14696 2043
rect -14758 1975 -14742 2009
rect -14708 1975 -14696 2009
rect -14758 1941 -14696 1975
rect -14758 1907 -14742 1941
rect -14708 1907 -14696 1941
rect -14758 1866 -14696 1907
rect -14526 2817 -14464 2858
rect -14526 2783 -14514 2817
rect -14480 2783 -14464 2817
rect -14526 2749 -14464 2783
rect -14526 2715 -14514 2749
rect -14480 2715 -14464 2749
rect -14526 2681 -14464 2715
rect -14526 2647 -14514 2681
rect -14480 2647 -14464 2681
rect -14526 2613 -14464 2647
rect -14526 2579 -14514 2613
rect -14480 2579 -14464 2613
rect -14526 2545 -14464 2579
rect -14526 2511 -14514 2545
rect -14480 2511 -14464 2545
rect -14526 2477 -14464 2511
rect -14526 2443 -14514 2477
rect -14480 2443 -14464 2477
rect -14526 2409 -14464 2443
rect -14526 2375 -14514 2409
rect -14480 2375 -14464 2409
rect -14526 2341 -14464 2375
rect -14526 2307 -14514 2341
rect -14480 2307 -14464 2341
rect -14526 2273 -14464 2307
rect -14526 2239 -14514 2273
rect -14480 2239 -14464 2273
rect -14526 2205 -14464 2239
rect -14526 2171 -14514 2205
rect -14480 2171 -14464 2205
rect -14526 2137 -14464 2171
rect -14526 2103 -14514 2137
rect -14480 2103 -14464 2137
rect -14526 2069 -14464 2103
rect -14526 2035 -14514 2069
rect -14480 2035 -14464 2069
rect -14526 2001 -14464 2035
rect -14526 1967 -14514 2001
rect -14480 1967 -14464 2001
rect -14526 1933 -14464 1967
rect -14526 1899 -14514 1933
rect -14480 1899 -14464 1933
rect -14526 1858 -14464 1899
rect -14434 2817 -14368 2858
rect -14434 2783 -14418 2817
rect -14384 2783 -14368 2817
rect -14434 2749 -14368 2783
rect -14434 2715 -14418 2749
rect -14384 2715 -14368 2749
rect -14434 2681 -14368 2715
rect -14434 2647 -14418 2681
rect -14384 2647 -14368 2681
rect -14434 2613 -14368 2647
rect -14434 2579 -14418 2613
rect -14384 2579 -14368 2613
rect -14434 2545 -14368 2579
rect -14434 2511 -14418 2545
rect -14384 2511 -14368 2545
rect -14434 2477 -14368 2511
rect -14434 2443 -14418 2477
rect -14384 2443 -14368 2477
rect -14434 2409 -14368 2443
rect -14434 2375 -14418 2409
rect -14384 2375 -14368 2409
rect -14434 2341 -14368 2375
rect -14434 2307 -14418 2341
rect -14384 2307 -14368 2341
rect -14434 2273 -14368 2307
rect -14434 2239 -14418 2273
rect -14384 2239 -14368 2273
rect -14434 2205 -14368 2239
rect -14434 2171 -14418 2205
rect -14384 2171 -14368 2205
rect -14434 2137 -14368 2171
rect -14434 2103 -14418 2137
rect -14384 2103 -14368 2137
rect -14434 2069 -14368 2103
rect -14434 2035 -14418 2069
rect -14384 2035 -14368 2069
rect -14434 2001 -14368 2035
rect -14434 1967 -14418 2001
rect -14384 1967 -14368 2001
rect -14434 1933 -14368 1967
rect -14434 1899 -14418 1933
rect -14384 1899 -14368 1933
rect -14434 1858 -14368 1899
rect -14338 2817 -14272 2858
rect -14338 2783 -14322 2817
rect -14288 2783 -14272 2817
rect -14338 2749 -14272 2783
rect -14338 2715 -14322 2749
rect -14288 2715 -14272 2749
rect -14338 2681 -14272 2715
rect -14338 2647 -14322 2681
rect -14288 2647 -14272 2681
rect -14338 2613 -14272 2647
rect -14338 2579 -14322 2613
rect -14288 2579 -14272 2613
rect -14338 2545 -14272 2579
rect -14338 2511 -14322 2545
rect -14288 2511 -14272 2545
rect -14338 2477 -14272 2511
rect -14338 2443 -14322 2477
rect -14288 2443 -14272 2477
rect -14338 2409 -14272 2443
rect -14338 2375 -14322 2409
rect -14288 2375 -14272 2409
rect -14338 2341 -14272 2375
rect -14338 2307 -14322 2341
rect -14288 2307 -14272 2341
rect -14338 2273 -14272 2307
rect -14338 2239 -14322 2273
rect -14288 2239 -14272 2273
rect -14338 2205 -14272 2239
rect -14338 2171 -14322 2205
rect -14288 2171 -14272 2205
rect -14338 2137 -14272 2171
rect -14338 2103 -14322 2137
rect -14288 2103 -14272 2137
rect -14338 2069 -14272 2103
rect -14338 2035 -14322 2069
rect -14288 2035 -14272 2069
rect -14338 2001 -14272 2035
rect -14338 1967 -14322 2001
rect -14288 1967 -14272 2001
rect -14338 1933 -14272 1967
rect -14338 1899 -14322 1933
rect -14288 1899 -14272 1933
rect -14338 1858 -14272 1899
rect -14242 2817 -14176 2858
rect -14242 2783 -14226 2817
rect -14192 2783 -14176 2817
rect -14242 2749 -14176 2783
rect -14242 2715 -14226 2749
rect -14192 2715 -14176 2749
rect -14242 2681 -14176 2715
rect -14242 2647 -14226 2681
rect -14192 2647 -14176 2681
rect -14242 2613 -14176 2647
rect -14242 2579 -14226 2613
rect -14192 2579 -14176 2613
rect -14242 2545 -14176 2579
rect -14242 2511 -14226 2545
rect -14192 2511 -14176 2545
rect -14242 2477 -14176 2511
rect -14242 2443 -14226 2477
rect -14192 2443 -14176 2477
rect -14242 2409 -14176 2443
rect -14242 2375 -14226 2409
rect -14192 2375 -14176 2409
rect -14242 2341 -14176 2375
rect -14242 2307 -14226 2341
rect -14192 2307 -14176 2341
rect -14242 2273 -14176 2307
rect -14242 2239 -14226 2273
rect -14192 2239 -14176 2273
rect -14242 2205 -14176 2239
rect -14242 2171 -14226 2205
rect -14192 2171 -14176 2205
rect -14242 2137 -14176 2171
rect -14242 2103 -14226 2137
rect -14192 2103 -14176 2137
rect -14242 2069 -14176 2103
rect -14242 2035 -14226 2069
rect -14192 2035 -14176 2069
rect -14242 2001 -14176 2035
rect -14242 1967 -14226 2001
rect -14192 1967 -14176 2001
rect -14242 1933 -14176 1967
rect -14242 1899 -14226 1933
rect -14192 1899 -14176 1933
rect -14242 1858 -14176 1899
rect -14146 2817 -14080 2858
rect -14146 2783 -14130 2817
rect -14096 2783 -14080 2817
rect -14146 2749 -14080 2783
rect -14146 2715 -14130 2749
rect -14096 2715 -14080 2749
rect -14146 2681 -14080 2715
rect -14146 2647 -14130 2681
rect -14096 2647 -14080 2681
rect -14146 2613 -14080 2647
rect -14146 2579 -14130 2613
rect -14096 2579 -14080 2613
rect -14146 2545 -14080 2579
rect -14146 2511 -14130 2545
rect -14096 2511 -14080 2545
rect -14146 2477 -14080 2511
rect -14146 2443 -14130 2477
rect -14096 2443 -14080 2477
rect -14146 2409 -14080 2443
rect -14146 2375 -14130 2409
rect -14096 2375 -14080 2409
rect -14146 2341 -14080 2375
rect -14146 2307 -14130 2341
rect -14096 2307 -14080 2341
rect -14146 2273 -14080 2307
rect -14146 2239 -14130 2273
rect -14096 2239 -14080 2273
rect -14146 2205 -14080 2239
rect -14146 2171 -14130 2205
rect -14096 2171 -14080 2205
rect -14146 2137 -14080 2171
rect -14146 2103 -14130 2137
rect -14096 2103 -14080 2137
rect -14146 2069 -14080 2103
rect -14146 2035 -14130 2069
rect -14096 2035 -14080 2069
rect -14146 2001 -14080 2035
rect -14146 1967 -14130 2001
rect -14096 1967 -14080 2001
rect -14146 1933 -14080 1967
rect -14146 1899 -14130 1933
rect -14096 1899 -14080 1933
rect -14146 1858 -14080 1899
rect -14050 2817 -13984 2858
rect -14050 2783 -14034 2817
rect -14000 2783 -13984 2817
rect -14050 2749 -13984 2783
rect -14050 2715 -14034 2749
rect -14000 2715 -13984 2749
rect -14050 2681 -13984 2715
rect -14050 2647 -14034 2681
rect -14000 2647 -13984 2681
rect -14050 2613 -13984 2647
rect -14050 2579 -14034 2613
rect -14000 2579 -13984 2613
rect -14050 2545 -13984 2579
rect -14050 2511 -14034 2545
rect -14000 2511 -13984 2545
rect -14050 2477 -13984 2511
rect -14050 2443 -14034 2477
rect -14000 2443 -13984 2477
rect -14050 2409 -13984 2443
rect -14050 2375 -14034 2409
rect -14000 2375 -13984 2409
rect -14050 2341 -13984 2375
rect -14050 2307 -14034 2341
rect -14000 2307 -13984 2341
rect -14050 2273 -13984 2307
rect -14050 2239 -14034 2273
rect -14000 2239 -13984 2273
rect -14050 2205 -13984 2239
rect -14050 2171 -14034 2205
rect -14000 2171 -13984 2205
rect -14050 2137 -13984 2171
rect -14050 2103 -14034 2137
rect -14000 2103 -13984 2137
rect -14050 2069 -13984 2103
rect -14050 2035 -14034 2069
rect -14000 2035 -13984 2069
rect -14050 2001 -13984 2035
rect -14050 1967 -14034 2001
rect -14000 1967 -13984 2001
rect -14050 1933 -13984 1967
rect -14050 1899 -14034 1933
rect -14000 1899 -13984 1933
rect -14050 1858 -13984 1899
rect -13954 2817 -13888 2858
rect -13954 2783 -13938 2817
rect -13904 2783 -13888 2817
rect -13954 2749 -13888 2783
rect -13954 2715 -13938 2749
rect -13904 2715 -13888 2749
rect -13954 2681 -13888 2715
rect -13954 2647 -13938 2681
rect -13904 2647 -13888 2681
rect -13954 2613 -13888 2647
rect -13954 2579 -13938 2613
rect -13904 2579 -13888 2613
rect -13954 2545 -13888 2579
rect -13954 2511 -13938 2545
rect -13904 2511 -13888 2545
rect -13954 2477 -13888 2511
rect -13954 2443 -13938 2477
rect -13904 2443 -13888 2477
rect -13954 2409 -13888 2443
rect -13954 2375 -13938 2409
rect -13904 2375 -13888 2409
rect -13954 2341 -13888 2375
rect -13954 2307 -13938 2341
rect -13904 2307 -13888 2341
rect -13954 2273 -13888 2307
rect -13954 2239 -13938 2273
rect -13904 2239 -13888 2273
rect -13954 2205 -13888 2239
rect -13954 2171 -13938 2205
rect -13904 2171 -13888 2205
rect -13954 2137 -13888 2171
rect -13954 2103 -13938 2137
rect -13904 2103 -13888 2137
rect -13954 2069 -13888 2103
rect -13954 2035 -13938 2069
rect -13904 2035 -13888 2069
rect -13954 2001 -13888 2035
rect -13954 1967 -13938 2001
rect -13904 1967 -13888 2001
rect -13954 1933 -13888 1967
rect -13954 1899 -13938 1933
rect -13904 1899 -13888 1933
rect -13954 1858 -13888 1899
rect -13858 2817 -13792 2858
rect -13858 2783 -13842 2817
rect -13808 2783 -13792 2817
rect -13858 2749 -13792 2783
rect -13858 2715 -13842 2749
rect -13808 2715 -13792 2749
rect -13858 2681 -13792 2715
rect -13858 2647 -13842 2681
rect -13808 2647 -13792 2681
rect -13858 2613 -13792 2647
rect -13858 2579 -13842 2613
rect -13808 2579 -13792 2613
rect -13858 2545 -13792 2579
rect -13858 2511 -13842 2545
rect -13808 2511 -13792 2545
rect -13858 2477 -13792 2511
rect -13858 2443 -13842 2477
rect -13808 2443 -13792 2477
rect -13858 2409 -13792 2443
rect -13858 2375 -13842 2409
rect -13808 2375 -13792 2409
rect -13858 2341 -13792 2375
rect -13858 2307 -13842 2341
rect -13808 2307 -13792 2341
rect -13858 2273 -13792 2307
rect -13858 2239 -13842 2273
rect -13808 2239 -13792 2273
rect -13858 2205 -13792 2239
rect -13858 2171 -13842 2205
rect -13808 2171 -13792 2205
rect -13858 2137 -13792 2171
rect -13858 2103 -13842 2137
rect -13808 2103 -13792 2137
rect -13858 2069 -13792 2103
rect -13858 2035 -13842 2069
rect -13808 2035 -13792 2069
rect -13858 2001 -13792 2035
rect -13858 1967 -13842 2001
rect -13808 1967 -13792 2001
rect -13858 1933 -13792 1967
rect -13858 1899 -13842 1933
rect -13808 1899 -13792 1933
rect -13858 1858 -13792 1899
rect -13762 2817 -13696 2858
rect -13762 2783 -13746 2817
rect -13712 2783 -13696 2817
rect -13762 2749 -13696 2783
rect -13762 2715 -13746 2749
rect -13712 2715 -13696 2749
rect -13762 2681 -13696 2715
rect -13762 2647 -13746 2681
rect -13712 2647 -13696 2681
rect -13762 2613 -13696 2647
rect -13762 2579 -13746 2613
rect -13712 2579 -13696 2613
rect -13762 2545 -13696 2579
rect -13762 2511 -13746 2545
rect -13712 2511 -13696 2545
rect -13762 2477 -13696 2511
rect -13762 2443 -13746 2477
rect -13712 2443 -13696 2477
rect -13762 2409 -13696 2443
rect -13762 2375 -13746 2409
rect -13712 2375 -13696 2409
rect -13762 2341 -13696 2375
rect -13762 2307 -13746 2341
rect -13712 2307 -13696 2341
rect -13762 2273 -13696 2307
rect -13762 2239 -13746 2273
rect -13712 2239 -13696 2273
rect -13762 2205 -13696 2239
rect -13762 2171 -13746 2205
rect -13712 2171 -13696 2205
rect -13762 2137 -13696 2171
rect -13762 2103 -13746 2137
rect -13712 2103 -13696 2137
rect -13762 2069 -13696 2103
rect -13762 2035 -13746 2069
rect -13712 2035 -13696 2069
rect -13762 2001 -13696 2035
rect -13762 1967 -13746 2001
rect -13712 1967 -13696 2001
rect -13762 1933 -13696 1967
rect -13762 1899 -13746 1933
rect -13712 1899 -13696 1933
rect -13762 1858 -13696 1899
rect -13666 2817 -13600 2858
rect -13666 2783 -13650 2817
rect -13616 2783 -13600 2817
rect -13666 2749 -13600 2783
rect -13666 2715 -13650 2749
rect -13616 2715 -13600 2749
rect -13666 2681 -13600 2715
rect -13666 2647 -13650 2681
rect -13616 2647 -13600 2681
rect -13666 2613 -13600 2647
rect -13666 2579 -13650 2613
rect -13616 2579 -13600 2613
rect -13666 2545 -13600 2579
rect -13666 2511 -13650 2545
rect -13616 2511 -13600 2545
rect -13666 2477 -13600 2511
rect -13666 2443 -13650 2477
rect -13616 2443 -13600 2477
rect -13666 2409 -13600 2443
rect -13666 2375 -13650 2409
rect -13616 2375 -13600 2409
rect -13666 2341 -13600 2375
rect -13666 2307 -13650 2341
rect -13616 2307 -13600 2341
rect -13666 2273 -13600 2307
rect -13666 2239 -13650 2273
rect -13616 2239 -13600 2273
rect -13666 2205 -13600 2239
rect -13666 2171 -13650 2205
rect -13616 2171 -13600 2205
rect -13666 2137 -13600 2171
rect -13666 2103 -13650 2137
rect -13616 2103 -13600 2137
rect -13666 2069 -13600 2103
rect -13666 2035 -13650 2069
rect -13616 2035 -13600 2069
rect -13666 2001 -13600 2035
rect -13666 1967 -13650 2001
rect -13616 1967 -13600 2001
rect -13666 1933 -13600 1967
rect -13666 1899 -13650 1933
rect -13616 1899 -13600 1933
rect -13666 1858 -13600 1899
rect -13570 2817 -13504 2858
rect -13570 2783 -13554 2817
rect -13520 2783 -13504 2817
rect -13570 2749 -13504 2783
rect -13570 2715 -13554 2749
rect -13520 2715 -13504 2749
rect -13570 2681 -13504 2715
rect -13570 2647 -13554 2681
rect -13520 2647 -13504 2681
rect -13570 2613 -13504 2647
rect -13570 2579 -13554 2613
rect -13520 2579 -13504 2613
rect -13570 2545 -13504 2579
rect -13570 2511 -13554 2545
rect -13520 2511 -13504 2545
rect -13570 2477 -13504 2511
rect -13570 2443 -13554 2477
rect -13520 2443 -13504 2477
rect -13570 2409 -13504 2443
rect -13570 2375 -13554 2409
rect -13520 2375 -13504 2409
rect -13570 2341 -13504 2375
rect -13570 2307 -13554 2341
rect -13520 2307 -13504 2341
rect -13570 2273 -13504 2307
rect -13570 2239 -13554 2273
rect -13520 2239 -13504 2273
rect -13570 2205 -13504 2239
rect -13570 2171 -13554 2205
rect -13520 2171 -13504 2205
rect -13570 2137 -13504 2171
rect -13570 2103 -13554 2137
rect -13520 2103 -13504 2137
rect -13570 2069 -13504 2103
rect -13570 2035 -13554 2069
rect -13520 2035 -13504 2069
rect -13570 2001 -13504 2035
rect -13570 1967 -13554 2001
rect -13520 1967 -13504 2001
rect -13570 1933 -13504 1967
rect -13570 1899 -13554 1933
rect -13520 1899 -13504 1933
rect -13570 1858 -13504 1899
rect -13474 2817 -13408 2858
rect -13474 2783 -13458 2817
rect -13424 2783 -13408 2817
rect -13474 2749 -13408 2783
rect -13474 2715 -13458 2749
rect -13424 2715 -13408 2749
rect -13474 2681 -13408 2715
rect -13474 2647 -13458 2681
rect -13424 2647 -13408 2681
rect -13474 2613 -13408 2647
rect -13474 2579 -13458 2613
rect -13424 2579 -13408 2613
rect -13474 2545 -13408 2579
rect -13474 2511 -13458 2545
rect -13424 2511 -13408 2545
rect -13474 2477 -13408 2511
rect -13474 2443 -13458 2477
rect -13424 2443 -13408 2477
rect -13474 2409 -13408 2443
rect -13474 2375 -13458 2409
rect -13424 2375 -13408 2409
rect -13474 2341 -13408 2375
rect -13474 2307 -13458 2341
rect -13424 2307 -13408 2341
rect -13474 2273 -13408 2307
rect -13474 2239 -13458 2273
rect -13424 2239 -13408 2273
rect -13474 2205 -13408 2239
rect -13474 2171 -13458 2205
rect -13424 2171 -13408 2205
rect -13474 2137 -13408 2171
rect -13474 2103 -13458 2137
rect -13424 2103 -13408 2137
rect -13474 2069 -13408 2103
rect -13474 2035 -13458 2069
rect -13424 2035 -13408 2069
rect -13474 2001 -13408 2035
rect -13474 1967 -13458 2001
rect -13424 1967 -13408 2001
rect -13474 1933 -13408 1967
rect -13474 1899 -13458 1933
rect -13424 1899 -13408 1933
rect -13474 1858 -13408 1899
rect -13378 2817 -13312 2858
rect -13378 2783 -13362 2817
rect -13328 2783 -13312 2817
rect -13378 2749 -13312 2783
rect -13378 2715 -13362 2749
rect -13328 2715 -13312 2749
rect -13378 2681 -13312 2715
rect -13378 2647 -13362 2681
rect -13328 2647 -13312 2681
rect -13378 2613 -13312 2647
rect -13378 2579 -13362 2613
rect -13328 2579 -13312 2613
rect -13378 2545 -13312 2579
rect -13378 2511 -13362 2545
rect -13328 2511 -13312 2545
rect -13378 2477 -13312 2511
rect -13378 2443 -13362 2477
rect -13328 2443 -13312 2477
rect -13378 2409 -13312 2443
rect -13378 2375 -13362 2409
rect -13328 2375 -13312 2409
rect -13378 2341 -13312 2375
rect -13378 2307 -13362 2341
rect -13328 2307 -13312 2341
rect -13378 2273 -13312 2307
rect -13378 2239 -13362 2273
rect -13328 2239 -13312 2273
rect -13378 2205 -13312 2239
rect -13378 2171 -13362 2205
rect -13328 2171 -13312 2205
rect -13378 2137 -13312 2171
rect -13378 2103 -13362 2137
rect -13328 2103 -13312 2137
rect -13378 2069 -13312 2103
rect -13378 2035 -13362 2069
rect -13328 2035 -13312 2069
rect -13378 2001 -13312 2035
rect -13378 1967 -13362 2001
rect -13328 1967 -13312 2001
rect -13378 1933 -13312 1967
rect -13378 1899 -13362 1933
rect -13328 1899 -13312 1933
rect -13378 1858 -13312 1899
rect -13282 2817 -13216 2858
rect -13282 2783 -13266 2817
rect -13232 2783 -13216 2817
rect -13282 2749 -13216 2783
rect -13282 2715 -13266 2749
rect -13232 2715 -13216 2749
rect -13282 2681 -13216 2715
rect -13282 2647 -13266 2681
rect -13232 2647 -13216 2681
rect -13282 2613 -13216 2647
rect -13282 2579 -13266 2613
rect -13232 2579 -13216 2613
rect -13282 2545 -13216 2579
rect -13282 2511 -13266 2545
rect -13232 2511 -13216 2545
rect -13282 2477 -13216 2511
rect -13282 2443 -13266 2477
rect -13232 2443 -13216 2477
rect -13282 2409 -13216 2443
rect -13282 2375 -13266 2409
rect -13232 2375 -13216 2409
rect -13282 2341 -13216 2375
rect -13282 2307 -13266 2341
rect -13232 2307 -13216 2341
rect -13282 2273 -13216 2307
rect -13282 2239 -13266 2273
rect -13232 2239 -13216 2273
rect -13282 2205 -13216 2239
rect -13282 2171 -13266 2205
rect -13232 2171 -13216 2205
rect -13282 2137 -13216 2171
rect -13282 2103 -13266 2137
rect -13232 2103 -13216 2137
rect -13282 2069 -13216 2103
rect -13282 2035 -13266 2069
rect -13232 2035 -13216 2069
rect -13282 2001 -13216 2035
rect -13282 1967 -13266 2001
rect -13232 1967 -13216 2001
rect -13282 1933 -13216 1967
rect -13282 1899 -13266 1933
rect -13232 1899 -13216 1933
rect -13282 1858 -13216 1899
rect -13186 2817 -13120 2858
rect -13186 2783 -13170 2817
rect -13136 2783 -13120 2817
rect -13186 2749 -13120 2783
rect -13186 2715 -13170 2749
rect -13136 2715 -13120 2749
rect -13186 2681 -13120 2715
rect -13186 2647 -13170 2681
rect -13136 2647 -13120 2681
rect -13186 2613 -13120 2647
rect -13186 2579 -13170 2613
rect -13136 2579 -13120 2613
rect -13186 2545 -13120 2579
rect -13186 2511 -13170 2545
rect -13136 2511 -13120 2545
rect -13186 2477 -13120 2511
rect -13186 2443 -13170 2477
rect -13136 2443 -13120 2477
rect -13186 2409 -13120 2443
rect -13186 2375 -13170 2409
rect -13136 2375 -13120 2409
rect -13186 2341 -13120 2375
rect -13186 2307 -13170 2341
rect -13136 2307 -13120 2341
rect -13186 2273 -13120 2307
rect -13186 2239 -13170 2273
rect -13136 2239 -13120 2273
rect -13186 2205 -13120 2239
rect -13186 2171 -13170 2205
rect -13136 2171 -13120 2205
rect -13186 2137 -13120 2171
rect -13186 2103 -13170 2137
rect -13136 2103 -13120 2137
rect -13186 2069 -13120 2103
rect -13186 2035 -13170 2069
rect -13136 2035 -13120 2069
rect -13186 2001 -13120 2035
rect -13186 1967 -13170 2001
rect -13136 1967 -13120 2001
rect -13186 1933 -13120 1967
rect -13186 1899 -13170 1933
rect -13136 1899 -13120 1933
rect -13186 1858 -13120 1899
rect -13090 2817 -13028 2858
rect -13090 2783 -13074 2817
rect -13040 2783 -13028 2817
rect -13090 2749 -13028 2783
rect -13090 2715 -13074 2749
rect -13040 2715 -13028 2749
rect -13090 2681 -13028 2715
rect -13090 2647 -13074 2681
rect -13040 2647 -13028 2681
rect -13090 2613 -13028 2647
rect -13090 2579 -13074 2613
rect -13040 2579 -13028 2613
rect -13090 2545 -13028 2579
rect -13090 2511 -13074 2545
rect -13040 2511 -13028 2545
rect -13090 2477 -13028 2511
rect -13090 2443 -13074 2477
rect -13040 2443 -13028 2477
rect -13090 2409 -13028 2443
rect -13090 2375 -13074 2409
rect -13040 2375 -13028 2409
rect -13090 2341 -13028 2375
rect -13090 2307 -13074 2341
rect -13040 2307 -13028 2341
rect -13090 2273 -13028 2307
rect -13090 2239 -13074 2273
rect -13040 2239 -13028 2273
rect -13090 2205 -13028 2239
rect -13090 2171 -13074 2205
rect -13040 2171 -13028 2205
rect -13090 2137 -13028 2171
rect -13090 2103 -13074 2137
rect -13040 2103 -13028 2137
rect -13090 2069 -13028 2103
rect -13090 2035 -13074 2069
rect -13040 2035 -13028 2069
rect -13090 2001 -13028 2035
rect -13090 1967 -13074 2001
rect -13040 1967 -13028 2001
rect -13090 1933 -13028 1967
rect -13090 1899 -13074 1933
rect -13040 1899 -13028 1933
rect -13090 1858 -13028 1899
rect -12848 2821 -12786 2862
rect -12848 2787 -12836 2821
rect -12802 2787 -12786 2821
rect -12848 2753 -12786 2787
rect -12848 2719 -12836 2753
rect -12802 2719 -12786 2753
rect -12848 2685 -12786 2719
rect -12848 2651 -12836 2685
rect -12802 2651 -12786 2685
rect -12848 2617 -12786 2651
rect -12848 2583 -12836 2617
rect -12802 2583 -12786 2617
rect -12848 2549 -12786 2583
rect -12848 2515 -12836 2549
rect -12802 2515 -12786 2549
rect -12848 2481 -12786 2515
rect -12848 2447 -12836 2481
rect -12802 2447 -12786 2481
rect -12848 2413 -12786 2447
rect -12848 2379 -12836 2413
rect -12802 2379 -12786 2413
rect -12848 2345 -12786 2379
rect -12848 2311 -12836 2345
rect -12802 2311 -12786 2345
rect -12848 2277 -12786 2311
rect -12848 2243 -12836 2277
rect -12802 2243 -12786 2277
rect -12848 2209 -12786 2243
rect -12848 2175 -12836 2209
rect -12802 2175 -12786 2209
rect -12848 2141 -12786 2175
rect -12848 2107 -12836 2141
rect -12802 2107 -12786 2141
rect -12848 2073 -12786 2107
rect -12848 2039 -12836 2073
rect -12802 2039 -12786 2073
rect -12848 2005 -12786 2039
rect -12848 1971 -12836 2005
rect -12802 1971 -12786 2005
rect -12848 1937 -12786 1971
rect -12848 1903 -12836 1937
rect -12802 1903 -12786 1937
rect -12848 1862 -12786 1903
rect -12756 2821 -12690 2862
rect -12756 2787 -12740 2821
rect -12706 2787 -12690 2821
rect -12756 2753 -12690 2787
rect -12756 2719 -12740 2753
rect -12706 2719 -12690 2753
rect -12756 2685 -12690 2719
rect -12756 2651 -12740 2685
rect -12706 2651 -12690 2685
rect -12756 2617 -12690 2651
rect -12756 2583 -12740 2617
rect -12706 2583 -12690 2617
rect -12756 2549 -12690 2583
rect -12756 2515 -12740 2549
rect -12706 2515 -12690 2549
rect -12756 2481 -12690 2515
rect -12756 2447 -12740 2481
rect -12706 2447 -12690 2481
rect -12756 2413 -12690 2447
rect -12756 2379 -12740 2413
rect -12706 2379 -12690 2413
rect -12756 2345 -12690 2379
rect -12756 2311 -12740 2345
rect -12706 2311 -12690 2345
rect -12756 2277 -12690 2311
rect -12756 2243 -12740 2277
rect -12706 2243 -12690 2277
rect -12756 2209 -12690 2243
rect -12756 2175 -12740 2209
rect -12706 2175 -12690 2209
rect -12756 2141 -12690 2175
rect -12756 2107 -12740 2141
rect -12706 2107 -12690 2141
rect -12756 2073 -12690 2107
rect -12756 2039 -12740 2073
rect -12706 2039 -12690 2073
rect -12756 2005 -12690 2039
rect -12756 1971 -12740 2005
rect -12706 1971 -12690 2005
rect -12756 1937 -12690 1971
rect -12756 1903 -12740 1937
rect -12706 1903 -12690 1937
rect -12756 1862 -12690 1903
rect -12660 2821 -12594 2862
rect -12660 2787 -12644 2821
rect -12610 2787 -12594 2821
rect -12660 2753 -12594 2787
rect -12660 2719 -12644 2753
rect -12610 2719 -12594 2753
rect -12660 2685 -12594 2719
rect -12660 2651 -12644 2685
rect -12610 2651 -12594 2685
rect -12660 2617 -12594 2651
rect -12660 2583 -12644 2617
rect -12610 2583 -12594 2617
rect -12660 2549 -12594 2583
rect -12660 2515 -12644 2549
rect -12610 2515 -12594 2549
rect -12660 2481 -12594 2515
rect -12660 2447 -12644 2481
rect -12610 2447 -12594 2481
rect -12660 2413 -12594 2447
rect -12660 2379 -12644 2413
rect -12610 2379 -12594 2413
rect -12660 2345 -12594 2379
rect -12660 2311 -12644 2345
rect -12610 2311 -12594 2345
rect -12660 2277 -12594 2311
rect -12660 2243 -12644 2277
rect -12610 2243 -12594 2277
rect -12660 2209 -12594 2243
rect -12660 2175 -12644 2209
rect -12610 2175 -12594 2209
rect -12660 2141 -12594 2175
rect -12660 2107 -12644 2141
rect -12610 2107 -12594 2141
rect -12660 2073 -12594 2107
rect -12660 2039 -12644 2073
rect -12610 2039 -12594 2073
rect -12660 2005 -12594 2039
rect -12660 1971 -12644 2005
rect -12610 1971 -12594 2005
rect -12660 1937 -12594 1971
rect -12660 1903 -12644 1937
rect -12610 1903 -12594 1937
rect -12660 1862 -12594 1903
rect -12564 2821 -12498 2862
rect -12564 2787 -12548 2821
rect -12514 2787 -12498 2821
rect -12564 2753 -12498 2787
rect -12564 2719 -12548 2753
rect -12514 2719 -12498 2753
rect -12564 2685 -12498 2719
rect -12564 2651 -12548 2685
rect -12514 2651 -12498 2685
rect -12564 2617 -12498 2651
rect -12564 2583 -12548 2617
rect -12514 2583 -12498 2617
rect -12564 2549 -12498 2583
rect -12564 2515 -12548 2549
rect -12514 2515 -12498 2549
rect -12564 2481 -12498 2515
rect -12564 2447 -12548 2481
rect -12514 2447 -12498 2481
rect -12564 2413 -12498 2447
rect -12564 2379 -12548 2413
rect -12514 2379 -12498 2413
rect -12564 2345 -12498 2379
rect -12564 2311 -12548 2345
rect -12514 2311 -12498 2345
rect -12564 2277 -12498 2311
rect -12564 2243 -12548 2277
rect -12514 2243 -12498 2277
rect -12564 2209 -12498 2243
rect -12564 2175 -12548 2209
rect -12514 2175 -12498 2209
rect -12564 2141 -12498 2175
rect -12564 2107 -12548 2141
rect -12514 2107 -12498 2141
rect -12564 2073 -12498 2107
rect -12564 2039 -12548 2073
rect -12514 2039 -12498 2073
rect -12564 2005 -12498 2039
rect -12564 1971 -12548 2005
rect -12514 1971 -12498 2005
rect -12564 1937 -12498 1971
rect -12564 1903 -12548 1937
rect -12514 1903 -12498 1937
rect -12564 1862 -12498 1903
rect -12468 2821 -12402 2862
rect -12468 2787 -12452 2821
rect -12418 2787 -12402 2821
rect -12468 2753 -12402 2787
rect -12468 2719 -12452 2753
rect -12418 2719 -12402 2753
rect -12468 2685 -12402 2719
rect -12468 2651 -12452 2685
rect -12418 2651 -12402 2685
rect -12468 2617 -12402 2651
rect -12468 2583 -12452 2617
rect -12418 2583 -12402 2617
rect -12468 2549 -12402 2583
rect -12468 2515 -12452 2549
rect -12418 2515 -12402 2549
rect -12468 2481 -12402 2515
rect -12468 2447 -12452 2481
rect -12418 2447 -12402 2481
rect -12468 2413 -12402 2447
rect -12468 2379 -12452 2413
rect -12418 2379 -12402 2413
rect -12468 2345 -12402 2379
rect -12468 2311 -12452 2345
rect -12418 2311 -12402 2345
rect -12468 2277 -12402 2311
rect -12468 2243 -12452 2277
rect -12418 2243 -12402 2277
rect -12468 2209 -12402 2243
rect -12468 2175 -12452 2209
rect -12418 2175 -12402 2209
rect -12468 2141 -12402 2175
rect -12468 2107 -12452 2141
rect -12418 2107 -12402 2141
rect -12468 2073 -12402 2107
rect -12468 2039 -12452 2073
rect -12418 2039 -12402 2073
rect -12468 2005 -12402 2039
rect -12468 1971 -12452 2005
rect -12418 1971 -12402 2005
rect -12468 1937 -12402 1971
rect -12468 1903 -12452 1937
rect -12418 1903 -12402 1937
rect -12468 1862 -12402 1903
rect -12372 2821 -12306 2862
rect -12372 2787 -12356 2821
rect -12322 2787 -12306 2821
rect -12372 2753 -12306 2787
rect -12372 2719 -12356 2753
rect -12322 2719 -12306 2753
rect -12372 2685 -12306 2719
rect -12372 2651 -12356 2685
rect -12322 2651 -12306 2685
rect -12372 2617 -12306 2651
rect -12372 2583 -12356 2617
rect -12322 2583 -12306 2617
rect -12372 2549 -12306 2583
rect -12372 2515 -12356 2549
rect -12322 2515 -12306 2549
rect -12372 2481 -12306 2515
rect -12372 2447 -12356 2481
rect -12322 2447 -12306 2481
rect -12372 2413 -12306 2447
rect -12372 2379 -12356 2413
rect -12322 2379 -12306 2413
rect -12372 2345 -12306 2379
rect -12372 2311 -12356 2345
rect -12322 2311 -12306 2345
rect -12372 2277 -12306 2311
rect -12372 2243 -12356 2277
rect -12322 2243 -12306 2277
rect -12372 2209 -12306 2243
rect -12372 2175 -12356 2209
rect -12322 2175 -12306 2209
rect -12372 2141 -12306 2175
rect -12372 2107 -12356 2141
rect -12322 2107 -12306 2141
rect -12372 2073 -12306 2107
rect -12372 2039 -12356 2073
rect -12322 2039 -12306 2073
rect -12372 2005 -12306 2039
rect -12372 1971 -12356 2005
rect -12322 1971 -12306 2005
rect -12372 1937 -12306 1971
rect -12372 1903 -12356 1937
rect -12322 1903 -12306 1937
rect -12372 1862 -12306 1903
rect -12276 2821 -12210 2862
rect -12276 2787 -12260 2821
rect -12226 2787 -12210 2821
rect -12276 2753 -12210 2787
rect -12276 2719 -12260 2753
rect -12226 2719 -12210 2753
rect -12276 2685 -12210 2719
rect -12276 2651 -12260 2685
rect -12226 2651 -12210 2685
rect -12276 2617 -12210 2651
rect -12276 2583 -12260 2617
rect -12226 2583 -12210 2617
rect -12276 2549 -12210 2583
rect -12276 2515 -12260 2549
rect -12226 2515 -12210 2549
rect -12276 2481 -12210 2515
rect -12276 2447 -12260 2481
rect -12226 2447 -12210 2481
rect -12276 2413 -12210 2447
rect -12276 2379 -12260 2413
rect -12226 2379 -12210 2413
rect -12276 2345 -12210 2379
rect -12276 2311 -12260 2345
rect -12226 2311 -12210 2345
rect -12276 2277 -12210 2311
rect -12276 2243 -12260 2277
rect -12226 2243 -12210 2277
rect -12276 2209 -12210 2243
rect -12276 2175 -12260 2209
rect -12226 2175 -12210 2209
rect -12276 2141 -12210 2175
rect -12276 2107 -12260 2141
rect -12226 2107 -12210 2141
rect -12276 2073 -12210 2107
rect -12276 2039 -12260 2073
rect -12226 2039 -12210 2073
rect -12276 2005 -12210 2039
rect -12276 1971 -12260 2005
rect -12226 1971 -12210 2005
rect -12276 1937 -12210 1971
rect -12276 1903 -12260 1937
rect -12226 1903 -12210 1937
rect -12276 1862 -12210 1903
rect -12180 2821 -12114 2862
rect -12180 2787 -12164 2821
rect -12130 2787 -12114 2821
rect -12180 2753 -12114 2787
rect -12180 2719 -12164 2753
rect -12130 2719 -12114 2753
rect -12180 2685 -12114 2719
rect -12180 2651 -12164 2685
rect -12130 2651 -12114 2685
rect -12180 2617 -12114 2651
rect -12180 2583 -12164 2617
rect -12130 2583 -12114 2617
rect -12180 2549 -12114 2583
rect -12180 2515 -12164 2549
rect -12130 2515 -12114 2549
rect -12180 2481 -12114 2515
rect -12180 2447 -12164 2481
rect -12130 2447 -12114 2481
rect -12180 2413 -12114 2447
rect -12180 2379 -12164 2413
rect -12130 2379 -12114 2413
rect -12180 2345 -12114 2379
rect -12180 2311 -12164 2345
rect -12130 2311 -12114 2345
rect -12180 2277 -12114 2311
rect -12180 2243 -12164 2277
rect -12130 2243 -12114 2277
rect -12180 2209 -12114 2243
rect -12180 2175 -12164 2209
rect -12130 2175 -12114 2209
rect -12180 2141 -12114 2175
rect -12180 2107 -12164 2141
rect -12130 2107 -12114 2141
rect -12180 2073 -12114 2107
rect -12180 2039 -12164 2073
rect -12130 2039 -12114 2073
rect -12180 2005 -12114 2039
rect -12180 1971 -12164 2005
rect -12130 1971 -12114 2005
rect -12180 1937 -12114 1971
rect -12180 1903 -12164 1937
rect -12130 1903 -12114 1937
rect -12180 1862 -12114 1903
rect -12084 2821 -12018 2862
rect -12084 2787 -12068 2821
rect -12034 2787 -12018 2821
rect -12084 2753 -12018 2787
rect -12084 2719 -12068 2753
rect -12034 2719 -12018 2753
rect -12084 2685 -12018 2719
rect -12084 2651 -12068 2685
rect -12034 2651 -12018 2685
rect -12084 2617 -12018 2651
rect -12084 2583 -12068 2617
rect -12034 2583 -12018 2617
rect -12084 2549 -12018 2583
rect -12084 2515 -12068 2549
rect -12034 2515 -12018 2549
rect -12084 2481 -12018 2515
rect -12084 2447 -12068 2481
rect -12034 2447 -12018 2481
rect -12084 2413 -12018 2447
rect -12084 2379 -12068 2413
rect -12034 2379 -12018 2413
rect -12084 2345 -12018 2379
rect -12084 2311 -12068 2345
rect -12034 2311 -12018 2345
rect -12084 2277 -12018 2311
rect -12084 2243 -12068 2277
rect -12034 2243 -12018 2277
rect -12084 2209 -12018 2243
rect -12084 2175 -12068 2209
rect -12034 2175 -12018 2209
rect -12084 2141 -12018 2175
rect -12084 2107 -12068 2141
rect -12034 2107 -12018 2141
rect -12084 2073 -12018 2107
rect -12084 2039 -12068 2073
rect -12034 2039 -12018 2073
rect -12084 2005 -12018 2039
rect -12084 1971 -12068 2005
rect -12034 1971 -12018 2005
rect -12084 1937 -12018 1971
rect -12084 1903 -12068 1937
rect -12034 1903 -12018 1937
rect -12084 1862 -12018 1903
rect -11988 2821 -11922 2862
rect -11988 2787 -11972 2821
rect -11938 2787 -11922 2821
rect -11988 2753 -11922 2787
rect -11988 2719 -11972 2753
rect -11938 2719 -11922 2753
rect -11988 2685 -11922 2719
rect -11988 2651 -11972 2685
rect -11938 2651 -11922 2685
rect -11988 2617 -11922 2651
rect -11988 2583 -11972 2617
rect -11938 2583 -11922 2617
rect -11988 2549 -11922 2583
rect -11988 2515 -11972 2549
rect -11938 2515 -11922 2549
rect -11988 2481 -11922 2515
rect -11988 2447 -11972 2481
rect -11938 2447 -11922 2481
rect -11988 2413 -11922 2447
rect -11988 2379 -11972 2413
rect -11938 2379 -11922 2413
rect -11988 2345 -11922 2379
rect -11988 2311 -11972 2345
rect -11938 2311 -11922 2345
rect -11988 2277 -11922 2311
rect -11988 2243 -11972 2277
rect -11938 2243 -11922 2277
rect -11988 2209 -11922 2243
rect -11988 2175 -11972 2209
rect -11938 2175 -11922 2209
rect -11988 2141 -11922 2175
rect -11988 2107 -11972 2141
rect -11938 2107 -11922 2141
rect -11988 2073 -11922 2107
rect -11988 2039 -11972 2073
rect -11938 2039 -11922 2073
rect -11988 2005 -11922 2039
rect -11988 1971 -11972 2005
rect -11938 1971 -11922 2005
rect -11988 1937 -11922 1971
rect -11988 1903 -11972 1937
rect -11938 1903 -11922 1937
rect -11988 1862 -11922 1903
rect -11892 2821 -11830 2862
rect -11892 2787 -11876 2821
rect -11842 2787 -11830 2821
rect -11892 2753 -11830 2787
rect -11892 2719 -11876 2753
rect -11842 2719 -11830 2753
rect -11892 2685 -11830 2719
rect -11892 2651 -11876 2685
rect -11842 2651 -11830 2685
rect -11892 2617 -11830 2651
rect -11892 2583 -11876 2617
rect -11842 2583 -11830 2617
rect -11892 2549 -11830 2583
rect -11892 2515 -11876 2549
rect -11842 2515 -11830 2549
rect -11892 2481 -11830 2515
rect -11892 2447 -11876 2481
rect -11842 2447 -11830 2481
rect -11892 2413 -11830 2447
rect -11892 2379 -11876 2413
rect -11842 2379 -11830 2413
rect -11892 2345 -11830 2379
rect -11892 2311 -11876 2345
rect -11842 2311 -11830 2345
rect -11892 2277 -11830 2311
rect -11892 2243 -11876 2277
rect -11842 2243 -11830 2277
rect -11892 2209 -11830 2243
rect -11892 2175 -11876 2209
rect -11842 2175 -11830 2209
rect -11892 2141 -11830 2175
rect -11892 2107 -11876 2141
rect -11842 2107 -11830 2141
rect -11892 2073 -11830 2107
rect -11892 2039 -11876 2073
rect -11842 2039 -11830 2073
rect -11892 2005 -11830 2039
rect -11892 1971 -11876 2005
rect -11842 1971 -11830 2005
rect -11892 1937 -11830 1971
rect -11892 1903 -11876 1937
rect -11842 1903 -11830 1937
rect -11892 1862 -11830 1903
rect -11676 2831 -11614 2872
rect -11676 2797 -11664 2831
rect -11630 2797 -11614 2831
rect -11676 2763 -11614 2797
rect -11676 2729 -11664 2763
rect -11630 2729 -11614 2763
rect -11676 2695 -11614 2729
rect -11676 2661 -11664 2695
rect -11630 2661 -11614 2695
rect -11676 2627 -11614 2661
rect -11676 2593 -11664 2627
rect -11630 2593 -11614 2627
rect -11676 2559 -11614 2593
rect -11676 2525 -11664 2559
rect -11630 2525 -11614 2559
rect -11676 2491 -11614 2525
rect -11676 2457 -11664 2491
rect -11630 2457 -11614 2491
rect -11676 2423 -11614 2457
rect -11676 2389 -11664 2423
rect -11630 2389 -11614 2423
rect -11676 2355 -11614 2389
rect -11676 2321 -11664 2355
rect -11630 2321 -11614 2355
rect -11676 2287 -11614 2321
rect -11676 2253 -11664 2287
rect -11630 2253 -11614 2287
rect -11676 2219 -11614 2253
rect -11676 2185 -11664 2219
rect -11630 2185 -11614 2219
rect -11676 2151 -11614 2185
rect -11676 2117 -11664 2151
rect -11630 2117 -11614 2151
rect -11676 2083 -11614 2117
rect -11676 2049 -11664 2083
rect -11630 2049 -11614 2083
rect -11676 2015 -11614 2049
rect -11676 1981 -11664 2015
rect -11630 1981 -11614 2015
rect -11676 1947 -11614 1981
rect -11676 1913 -11664 1947
rect -11630 1913 -11614 1947
rect -11676 1872 -11614 1913
rect -11584 2831 -11518 2872
rect -11584 2797 -11568 2831
rect -11534 2797 -11518 2831
rect -11584 2763 -11518 2797
rect -11584 2729 -11568 2763
rect -11534 2729 -11518 2763
rect -11584 2695 -11518 2729
rect -11584 2661 -11568 2695
rect -11534 2661 -11518 2695
rect -11584 2627 -11518 2661
rect -11584 2593 -11568 2627
rect -11534 2593 -11518 2627
rect -11584 2559 -11518 2593
rect -11584 2525 -11568 2559
rect -11534 2525 -11518 2559
rect -11584 2491 -11518 2525
rect -11584 2457 -11568 2491
rect -11534 2457 -11518 2491
rect -11584 2423 -11518 2457
rect -11584 2389 -11568 2423
rect -11534 2389 -11518 2423
rect -11584 2355 -11518 2389
rect -11584 2321 -11568 2355
rect -11534 2321 -11518 2355
rect -11584 2287 -11518 2321
rect -11584 2253 -11568 2287
rect -11534 2253 -11518 2287
rect -11584 2219 -11518 2253
rect -11584 2185 -11568 2219
rect -11534 2185 -11518 2219
rect -11584 2151 -11518 2185
rect -11584 2117 -11568 2151
rect -11534 2117 -11518 2151
rect -11584 2083 -11518 2117
rect -11584 2049 -11568 2083
rect -11534 2049 -11518 2083
rect -11584 2015 -11518 2049
rect -11584 1981 -11568 2015
rect -11534 1981 -11518 2015
rect -11584 1947 -11518 1981
rect -11584 1913 -11568 1947
rect -11534 1913 -11518 1947
rect -11584 1872 -11518 1913
rect -11488 2831 -11422 2872
rect -11488 2797 -11472 2831
rect -11438 2797 -11422 2831
rect -11488 2763 -11422 2797
rect -11488 2729 -11472 2763
rect -11438 2729 -11422 2763
rect -11488 2695 -11422 2729
rect -11488 2661 -11472 2695
rect -11438 2661 -11422 2695
rect -11488 2627 -11422 2661
rect -11488 2593 -11472 2627
rect -11438 2593 -11422 2627
rect -11488 2559 -11422 2593
rect -11488 2525 -11472 2559
rect -11438 2525 -11422 2559
rect -11488 2491 -11422 2525
rect -11488 2457 -11472 2491
rect -11438 2457 -11422 2491
rect -11488 2423 -11422 2457
rect -11488 2389 -11472 2423
rect -11438 2389 -11422 2423
rect -11488 2355 -11422 2389
rect -11488 2321 -11472 2355
rect -11438 2321 -11422 2355
rect -11488 2287 -11422 2321
rect -11488 2253 -11472 2287
rect -11438 2253 -11422 2287
rect -11488 2219 -11422 2253
rect -11488 2185 -11472 2219
rect -11438 2185 -11422 2219
rect -11488 2151 -11422 2185
rect -11488 2117 -11472 2151
rect -11438 2117 -11422 2151
rect -11488 2083 -11422 2117
rect -11488 2049 -11472 2083
rect -11438 2049 -11422 2083
rect -11488 2015 -11422 2049
rect -11488 1981 -11472 2015
rect -11438 1981 -11422 2015
rect -11488 1947 -11422 1981
rect -11488 1913 -11472 1947
rect -11438 1913 -11422 1947
rect -11488 1872 -11422 1913
rect -11392 2831 -11326 2872
rect -11392 2797 -11376 2831
rect -11342 2797 -11326 2831
rect -11392 2763 -11326 2797
rect -11392 2729 -11376 2763
rect -11342 2729 -11326 2763
rect -11392 2695 -11326 2729
rect -11392 2661 -11376 2695
rect -11342 2661 -11326 2695
rect -11392 2627 -11326 2661
rect -11392 2593 -11376 2627
rect -11342 2593 -11326 2627
rect -11392 2559 -11326 2593
rect -11392 2525 -11376 2559
rect -11342 2525 -11326 2559
rect -11392 2491 -11326 2525
rect -11392 2457 -11376 2491
rect -11342 2457 -11326 2491
rect -11392 2423 -11326 2457
rect -11392 2389 -11376 2423
rect -11342 2389 -11326 2423
rect -11392 2355 -11326 2389
rect -11392 2321 -11376 2355
rect -11342 2321 -11326 2355
rect -11392 2287 -11326 2321
rect -11392 2253 -11376 2287
rect -11342 2253 -11326 2287
rect -11392 2219 -11326 2253
rect -11392 2185 -11376 2219
rect -11342 2185 -11326 2219
rect -11392 2151 -11326 2185
rect -11392 2117 -11376 2151
rect -11342 2117 -11326 2151
rect -11392 2083 -11326 2117
rect -11392 2049 -11376 2083
rect -11342 2049 -11326 2083
rect -11392 2015 -11326 2049
rect -11392 1981 -11376 2015
rect -11342 1981 -11326 2015
rect -11392 1947 -11326 1981
rect -11392 1913 -11376 1947
rect -11342 1913 -11326 1947
rect -11392 1872 -11326 1913
rect -11296 2831 -11230 2872
rect -11296 2797 -11280 2831
rect -11246 2797 -11230 2831
rect -11296 2763 -11230 2797
rect -11296 2729 -11280 2763
rect -11246 2729 -11230 2763
rect -11296 2695 -11230 2729
rect -11296 2661 -11280 2695
rect -11246 2661 -11230 2695
rect -11296 2627 -11230 2661
rect -11296 2593 -11280 2627
rect -11246 2593 -11230 2627
rect -11296 2559 -11230 2593
rect -11296 2525 -11280 2559
rect -11246 2525 -11230 2559
rect -11296 2491 -11230 2525
rect -11296 2457 -11280 2491
rect -11246 2457 -11230 2491
rect -11296 2423 -11230 2457
rect -11296 2389 -11280 2423
rect -11246 2389 -11230 2423
rect -11296 2355 -11230 2389
rect -11296 2321 -11280 2355
rect -11246 2321 -11230 2355
rect -11296 2287 -11230 2321
rect -11296 2253 -11280 2287
rect -11246 2253 -11230 2287
rect -11296 2219 -11230 2253
rect -11296 2185 -11280 2219
rect -11246 2185 -11230 2219
rect -11296 2151 -11230 2185
rect -11296 2117 -11280 2151
rect -11246 2117 -11230 2151
rect -11296 2083 -11230 2117
rect -11296 2049 -11280 2083
rect -11246 2049 -11230 2083
rect -11296 2015 -11230 2049
rect -11296 1981 -11280 2015
rect -11246 1981 -11230 2015
rect -11296 1947 -11230 1981
rect -11296 1913 -11280 1947
rect -11246 1913 -11230 1947
rect -11296 1872 -11230 1913
rect -11200 2831 -11138 2872
rect -11200 2797 -11184 2831
rect -11150 2797 -11138 2831
rect -11200 2763 -11138 2797
rect -11200 2729 -11184 2763
rect -11150 2729 -11138 2763
rect -11200 2695 -11138 2729
rect -11200 2661 -11184 2695
rect -11150 2661 -11138 2695
rect -11200 2627 -11138 2661
rect -11200 2593 -11184 2627
rect -11150 2593 -11138 2627
rect -11200 2559 -11138 2593
rect -11200 2525 -11184 2559
rect -11150 2525 -11138 2559
rect -11200 2491 -11138 2525
rect -11200 2457 -11184 2491
rect -11150 2457 -11138 2491
rect -11200 2423 -11138 2457
rect -11200 2389 -11184 2423
rect -11150 2389 -11138 2423
rect -11200 2355 -11138 2389
rect -11200 2321 -11184 2355
rect -11150 2321 -11138 2355
rect -11200 2287 -11138 2321
rect -11200 2253 -11184 2287
rect -11150 2253 -11138 2287
rect -11200 2219 -11138 2253
rect -11200 2185 -11184 2219
rect -11150 2185 -11138 2219
rect -11200 2151 -11138 2185
rect -11200 2117 -11184 2151
rect -11150 2117 -11138 2151
rect -11200 2083 -11138 2117
rect -11200 2049 -11184 2083
rect -11150 2049 -11138 2083
rect -11200 2015 -11138 2049
rect -11200 1981 -11184 2015
rect -11150 1981 -11138 2015
rect -11200 1947 -11138 1981
rect -11200 1913 -11184 1947
rect -11150 1913 -11138 1947
rect -11200 1872 -11138 1913
rect -10208 2823 -10146 2864
rect -10208 2789 -10196 2823
rect -10162 2789 -10146 2823
rect -10208 2755 -10146 2789
rect -10208 2721 -10196 2755
rect -10162 2721 -10146 2755
rect -10208 2687 -10146 2721
rect -10208 2653 -10196 2687
rect -10162 2653 -10146 2687
rect -10208 2619 -10146 2653
rect -10208 2585 -10196 2619
rect -10162 2585 -10146 2619
rect -10208 2551 -10146 2585
rect -10208 2517 -10196 2551
rect -10162 2517 -10146 2551
rect -10208 2483 -10146 2517
rect -10208 2449 -10196 2483
rect -10162 2449 -10146 2483
rect -10208 2415 -10146 2449
rect -10208 2381 -10196 2415
rect -10162 2381 -10146 2415
rect -10208 2347 -10146 2381
rect -10208 2313 -10196 2347
rect -10162 2313 -10146 2347
rect -10208 2279 -10146 2313
rect -10208 2245 -10196 2279
rect -10162 2245 -10146 2279
rect -10208 2211 -10146 2245
rect -10208 2177 -10196 2211
rect -10162 2177 -10146 2211
rect -10208 2143 -10146 2177
rect -10208 2109 -10196 2143
rect -10162 2109 -10146 2143
rect -10208 2075 -10146 2109
rect -10208 2041 -10196 2075
rect -10162 2041 -10146 2075
rect -10208 2007 -10146 2041
rect -10208 1973 -10196 2007
rect -10162 1973 -10146 2007
rect -10208 1939 -10146 1973
rect -10208 1905 -10196 1939
rect -10162 1905 -10146 1939
rect -10208 1864 -10146 1905
rect -10116 2823 -10050 2864
rect -10116 2789 -10100 2823
rect -10066 2789 -10050 2823
rect -10116 2755 -10050 2789
rect -10116 2721 -10100 2755
rect -10066 2721 -10050 2755
rect -10116 2687 -10050 2721
rect -10116 2653 -10100 2687
rect -10066 2653 -10050 2687
rect -10116 2619 -10050 2653
rect -10116 2585 -10100 2619
rect -10066 2585 -10050 2619
rect -10116 2551 -10050 2585
rect -10116 2517 -10100 2551
rect -10066 2517 -10050 2551
rect -10116 2483 -10050 2517
rect -10116 2449 -10100 2483
rect -10066 2449 -10050 2483
rect -10116 2415 -10050 2449
rect -10116 2381 -10100 2415
rect -10066 2381 -10050 2415
rect -10116 2347 -10050 2381
rect -10116 2313 -10100 2347
rect -10066 2313 -10050 2347
rect -10116 2279 -10050 2313
rect -10116 2245 -10100 2279
rect -10066 2245 -10050 2279
rect -10116 2211 -10050 2245
rect -10116 2177 -10100 2211
rect -10066 2177 -10050 2211
rect -10116 2143 -10050 2177
rect -10116 2109 -10100 2143
rect -10066 2109 -10050 2143
rect -10116 2075 -10050 2109
rect -10116 2041 -10100 2075
rect -10066 2041 -10050 2075
rect -10116 2007 -10050 2041
rect -10116 1973 -10100 2007
rect -10066 1973 -10050 2007
rect -10116 1939 -10050 1973
rect -10116 1905 -10100 1939
rect -10066 1905 -10050 1939
rect -10116 1864 -10050 1905
rect -10020 2823 -9954 2864
rect -10020 2789 -10004 2823
rect -9970 2789 -9954 2823
rect -10020 2755 -9954 2789
rect -10020 2721 -10004 2755
rect -9970 2721 -9954 2755
rect -10020 2687 -9954 2721
rect -10020 2653 -10004 2687
rect -9970 2653 -9954 2687
rect -10020 2619 -9954 2653
rect -10020 2585 -10004 2619
rect -9970 2585 -9954 2619
rect -10020 2551 -9954 2585
rect -10020 2517 -10004 2551
rect -9970 2517 -9954 2551
rect -10020 2483 -9954 2517
rect -10020 2449 -10004 2483
rect -9970 2449 -9954 2483
rect -10020 2415 -9954 2449
rect -10020 2381 -10004 2415
rect -9970 2381 -9954 2415
rect -10020 2347 -9954 2381
rect -10020 2313 -10004 2347
rect -9970 2313 -9954 2347
rect -10020 2279 -9954 2313
rect -10020 2245 -10004 2279
rect -9970 2245 -9954 2279
rect -10020 2211 -9954 2245
rect -10020 2177 -10004 2211
rect -9970 2177 -9954 2211
rect -10020 2143 -9954 2177
rect -10020 2109 -10004 2143
rect -9970 2109 -9954 2143
rect -10020 2075 -9954 2109
rect -10020 2041 -10004 2075
rect -9970 2041 -9954 2075
rect -10020 2007 -9954 2041
rect -10020 1973 -10004 2007
rect -9970 1973 -9954 2007
rect -10020 1939 -9954 1973
rect -10020 1905 -10004 1939
rect -9970 1905 -9954 1939
rect -10020 1864 -9954 1905
rect -9924 2823 -9858 2864
rect -9924 2789 -9908 2823
rect -9874 2789 -9858 2823
rect -9924 2755 -9858 2789
rect -9924 2721 -9908 2755
rect -9874 2721 -9858 2755
rect -9924 2687 -9858 2721
rect -9924 2653 -9908 2687
rect -9874 2653 -9858 2687
rect -9924 2619 -9858 2653
rect -9924 2585 -9908 2619
rect -9874 2585 -9858 2619
rect -9924 2551 -9858 2585
rect -9924 2517 -9908 2551
rect -9874 2517 -9858 2551
rect -9924 2483 -9858 2517
rect -9924 2449 -9908 2483
rect -9874 2449 -9858 2483
rect -9924 2415 -9858 2449
rect -9924 2381 -9908 2415
rect -9874 2381 -9858 2415
rect -9924 2347 -9858 2381
rect -9924 2313 -9908 2347
rect -9874 2313 -9858 2347
rect -9924 2279 -9858 2313
rect -9924 2245 -9908 2279
rect -9874 2245 -9858 2279
rect -9924 2211 -9858 2245
rect -9924 2177 -9908 2211
rect -9874 2177 -9858 2211
rect -9924 2143 -9858 2177
rect -9924 2109 -9908 2143
rect -9874 2109 -9858 2143
rect -9924 2075 -9858 2109
rect -9924 2041 -9908 2075
rect -9874 2041 -9858 2075
rect -9924 2007 -9858 2041
rect -9924 1973 -9908 2007
rect -9874 1973 -9858 2007
rect -9924 1939 -9858 1973
rect -9924 1905 -9908 1939
rect -9874 1905 -9858 1939
rect -9924 1864 -9858 1905
rect -9828 2823 -9762 2864
rect -9828 2789 -9812 2823
rect -9778 2789 -9762 2823
rect -9828 2755 -9762 2789
rect -9828 2721 -9812 2755
rect -9778 2721 -9762 2755
rect -9828 2687 -9762 2721
rect -9828 2653 -9812 2687
rect -9778 2653 -9762 2687
rect -9828 2619 -9762 2653
rect -9828 2585 -9812 2619
rect -9778 2585 -9762 2619
rect -9828 2551 -9762 2585
rect -9828 2517 -9812 2551
rect -9778 2517 -9762 2551
rect -9828 2483 -9762 2517
rect -9828 2449 -9812 2483
rect -9778 2449 -9762 2483
rect -9828 2415 -9762 2449
rect -9828 2381 -9812 2415
rect -9778 2381 -9762 2415
rect -9828 2347 -9762 2381
rect -9828 2313 -9812 2347
rect -9778 2313 -9762 2347
rect -9828 2279 -9762 2313
rect -9828 2245 -9812 2279
rect -9778 2245 -9762 2279
rect -9828 2211 -9762 2245
rect -9828 2177 -9812 2211
rect -9778 2177 -9762 2211
rect -9828 2143 -9762 2177
rect -9828 2109 -9812 2143
rect -9778 2109 -9762 2143
rect -9828 2075 -9762 2109
rect -9828 2041 -9812 2075
rect -9778 2041 -9762 2075
rect -9828 2007 -9762 2041
rect -9828 1973 -9812 2007
rect -9778 1973 -9762 2007
rect -9828 1939 -9762 1973
rect -9828 1905 -9812 1939
rect -9778 1905 -9762 1939
rect -9828 1864 -9762 1905
rect -9732 2823 -9666 2864
rect -9732 2789 -9716 2823
rect -9682 2789 -9666 2823
rect -9732 2755 -9666 2789
rect -9732 2721 -9716 2755
rect -9682 2721 -9666 2755
rect -9732 2687 -9666 2721
rect -9732 2653 -9716 2687
rect -9682 2653 -9666 2687
rect -9732 2619 -9666 2653
rect -9732 2585 -9716 2619
rect -9682 2585 -9666 2619
rect -9732 2551 -9666 2585
rect -9732 2517 -9716 2551
rect -9682 2517 -9666 2551
rect -9732 2483 -9666 2517
rect -9732 2449 -9716 2483
rect -9682 2449 -9666 2483
rect -9732 2415 -9666 2449
rect -9732 2381 -9716 2415
rect -9682 2381 -9666 2415
rect -9732 2347 -9666 2381
rect -9732 2313 -9716 2347
rect -9682 2313 -9666 2347
rect -9732 2279 -9666 2313
rect -9732 2245 -9716 2279
rect -9682 2245 -9666 2279
rect -9732 2211 -9666 2245
rect -9732 2177 -9716 2211
rect -9682 2177 -9666 2211
rect -9732 2143 -9666 2177
rect -9732 2109 -9716 2143
rect -9682 2109 -9666 2143
rect -9732 2075 -9666 2109
rect -9732 2041 -9716 2075
rect -9682 2041 -9666 2075
rect -9732 2007 -9666 2041
rect -9732 1973 -9716 2007
rect -9682 1973 -9666 2007
rect -9732 1939 -9666 1973
rect -9732 1905 -9716 1939
rect -9682 1905 -9666 1939
rect -9732 1864 -9666 1905
rect -9636 2823 -9570 2864
rect -9636 2789 -9620 2823
rect -9586 2789 -9570 2823
rect -9636 2755 -9570 2789
rect -9636 2721 -9620 2755
rect -9586 2721 -9570 2755
rect -9636 2687 -9570 2721
rect -9636 2653 -9620 2687
rect -9586 2653 -9570 2687
rect -9636 2619 -9570 2653
rect -9636 2585 -9620 2619
rect -9586 2585 -9570 2619
rect -9636 2551 -9570 2585
rect -9636 2517 -9620 2551
rect -9586 2517 -9570 2551
rect -9636 2483 -9570 2517
rect -9636 2449 -9620 2483
rect -9586 2449 -9570 2483
rect -9636 2415 -9570 2449
rect -9636 2381 -9620 2415
rect -9586 2381 -9570 2415
rect -9636 2347 -9570 2381
rect -9636 2313 -9620 2347
rect -9586 2313 -9570 2347
rect -9636 2279 -9570 2313
rect -9636 2245 -9620 2279
rect -9586 2245 -9570 2279
rect -9636 2211 -9570 2245
rect -9636 2177 -9620 2211
rect -9586 2177 -9570 2211
rect -9636 2143 -9570 2177
rect -9636 2109 -9620 2143
rect -9586 2109 -9570 2143
rect -9636 2075 -9570 2109
rect -9636 2041 -9620 2075
rect -9586 2041 -9570 2075
rect -9636 2007 -9570 2041
rect -9636 1973 -9620 2007
rect -9586 1973 -9570 2007
rect -9636 1939 -9570 1973
rect -9636 1905 -9620 1939
rect -9586 1905 -9570 1939
rect -9636 1864 -9570 1905
rect -9540 2823 -9474 2864
rect -9540 2789 -9524 2823
rect -9490 2789 -9474 2823
rect -9540 2755 -9474 2789
rect -9540 2721 -9524 2755
rect -9490 2721 -9474 2755
rect -9540 2687 -9474 2721
rect -9540 2653 -9524 2687
rect -9490 2653 -9474 2687
rect -9540 2619 -9474 2653
rect -9540 2585 -9524 2619
rect -9490 2585 -9474 2619
rect -9540 2551 -9474 2585
rect -9540 2517 -9524 2551
rect -9490 2517 -9474 2551
rect -9540 2483 -9474 2517
rect -9540 2449 -9524 2483
rect -9490 2449 -9474 2483
rect -9540 2415 -9474 2449
rect -9540 2381 -9524 2415
rect -9490 2381 -9474 2415
rect -9540 2347 -9474 2381
rect -9540 2313 -9524 2347
rect -9490 2313 -9474 2347
rect -9540 2279 -9474 2313
rect -9540 2245 -9524 2279
rect -9490 2245 -9474 2279
rect -9540 2211 -9474 2245
rect -9540 2177 -9524 2211
rect -9490 2177 -9474 2211
rect -9540 2143 -9474 2177
rect -9540 2109 -9524 2143
rect -9490 2109 -9474 2143
rect -9540 2075 -9474 2109
rect -9540 2041 -9524 2075
rect -9490 2041 -9474 2075
rect -9540 2007 -9474 2041
rect -9540 1973 -9524 2007
rect -9490 1973 -9474 2007
rect -9540 1939 -9474 1973
rect -9540 1905 -9524 1939
rect -9490 1905 -9474 1939
rect -9540 1864 -9474 1905
rect -9444 2823 -9378 2864
rect -9444 2789 -9428 2823
rect -9394 2789 -9378 2823
rect -9444 2755 -9378 2789
rect -9444 2721 -9428 2755
rect -9394 2721 -9378 2755
rect -9444 2687 -9378 2721
rect -9444 2653 -9428 2687
rect -9394 2653 -9378 2687
rect -9444 2619 -9378 2653
rect -9444 2585 -9428 2619
rect -9394 2585 -9378 2619
rect -9444 2551 -9378 2585
rect -9444 2517 -9428 2551
rect -9394 2517 -9378 2551
rect -9444 2483 -9378 2517
rect -9444 2449 -9428 2483
rect -9394 2449 -9378 2483
rect -9444 2415 -9378 2449
rect -9444 2381 -9428 2415
rect -9394 2381 -9378 2415
rect -9444 2347 -9378 2381
rect -9444 2313 -9428 2347
rect -9394 2313 -9378 2347
rect -9444 2279 -9378 2313
rect -9444 2245 -9428 2279
rect -9394 2245 -9378 2279
rect -9444 2211 -9378 2245
rect -9444 2177 -9428 2211
rect -9394 2177 -9378 2211
rect -9444 2143 -9378 2177
rect -9444 2109 -9428 2143
rect -9394 2109 -9378 2143
rect -9444 2075 -9378 2109
rect -9444 2041 -9428 2075
rect -9394 2041 -9378 2075
rect -9444 2007 -9378 2041
rect -9444 1973 -9428 2007
rect -9394 1973 -9378 2007
rect -9444 1939 -9378 1973
rect -9444 1905 -9428 1939
rect -9394 1905 -9378 1939
rect -9444 1864 -9378 1905
rect -9348 2823 -9282 2864
rect -9348 2789 -9332 2823
rect -9298 2789 -9282 2823
rect -9348 2755 -9282 2789
rect -9348 2721 -9332 2755
rect -9298 2721 -9282 2755
rect -9348 2687 -9282 2721
rect -9348 2653 -9332 2687
rect -9298 2653 -9282 2687
rect -9348 2619 -9282 2653
rect -9348 2585 -9332 2619
rect -9298 2585 -9282 2619
rect -9348 2551 -9282 2585
rect -9348 2517 -9332 2551
rect -9298 2517 -9282 2551
rect -9348 2483 -9282 2517
rect -9348 2449 -9332 2483
rect -9298 2449 -9282 2483
rect -9348 2415 -9282 2449
rect -9348 2381 -9332 2415
rect -9298 2381 -9282 2415
rect -9348 2347 -9282 2381
rect -9348 2313 -9332 2347
rect -9298 2313 -9282 2347
rect -9348 2279 -9282 2313
rect -9348 2245 -9332 2279
rect -9298 2245 -9282 2279
rect -9348 2211 -9282 2245
rect -9348 2177 -9332 2211
rect -9298 2177 -9282 2211
rect -9348 2143 -9282 2177
rect -9348 2109 -9332 2143
rect -9298 2109 -9282 2143
rect -9348 2075 -9282 2109
rect -9348 2041 -9332 2075
rect -9298 2041 -9282 2075
rect -9348 2007 -9282 2041
rect -9348 1973 -9332 2007
rect -9298 1973 -9282 2007
rect -9348 1939 -9282 1973
rect -9348 1905 -9332 1939
rect -9298 1905 -9282 1939
rect -9348 1864 -9282 1905
rect -9252 2823 -9186 2864
rect -9252 2789 -9236 2823
rect -9202 2789 -9186 2823
rect -9252 2755 -9186 2789
rect -9252 2721 -9236 2755
rect -9202 2721 -9186 2755
rect -9252 2687 -9186 2721
rect -9252 2653 -9236 2687
rect -9202 2653 -9186 2687
rect -9252 2619 -9186 2653
rect -9252 2585 -9236 2619
rect -9202 2585 -9186 2619
rect -9252 2551 -9186 2585
rect -9252 2517 -9236 2551
rect -9202 2517 -9186 2551
rect -9252 2483 -9186 2517
rect -9252 2449 -9236 2483
rect -9202 2449 -9186 2483
rect -9252 2415 -9186 2449
rect -9252 2381 -9236 2415
rect -9202 2381 -9186 2415
rect -9252 2347 -9186 2381
rect -9252 2313 -9236 2347
rect -9202 2313 -9186 2347
rect -9252 2279 -9186 2313
rect -9252 2245 -9236 2279
rect -9202 2245 -9186 2279
rect -9252 2211 -9186 2245
rect -9252 2177 -9236 2211
rect -9202 2177 -9186 2211
rect -9252 2143 -9186 2177
rect -9252 2109 -9236 2143
rect -9202 2109 -9186 2143
rect -9252 2075 -9186 2109
rect -9252 2041 -9236 2075
rect -9202 2041 -9186 2075
rect -9252 2007 -9186 2041
rect -9252 1973 -9236 2007
rect -9202 1973 -9186 2007
rect -9252 1939 -9186 1973
rect -9252 1905 -9236 1939
rect -9202 1905 -9186 1939
rect -9252 1864 -9186 1905
rect -9156 2823 -9090 2864
rect -9156 2789 -9140 2823
rect -9106 2789 -9090 2823
rect -9156 2755 -9090 2789
rect -9156 2721 -9140 2755
rect -9106 2721 -9090 2755
rect -9156 2687 -9090 2721
rect -9156 2653 -9140 2687
rect -9106 2653 -9090 2687
rect -9156 2619 -9090 2653
rect -9156 2585 -9140 2619
rect -9106 2585 -9090 2619
rect -9156 2551 -9090 2585
rect -9156 2517 -9140 2551
rect -9106 2517 -9090 2551
rect -9156 2483 -9090 2517
rect -9156 2449 -9140 2483
rect -9106 2449 -9090 2483
rect -9156 2415 -9090 2449
rect -9156 2381 -9140 2415
rect -9106 2381 -9090 2415
rect -9156 2347 -9090 2381
rect -9156 2313 -9140 2347
rect -9106 2313 -9090 2347
rect -9156 2279 -9090 2313
rect -9156 2245 -9140 2279
rect -9106 2245 -9090 2279
rect -9156 2211 -9090 2245
rect -9156 2177 -9140 2211
rect -9106 2177 -9090 2211
rect -9156 2143 -9090 2177
rect -9156 2109 -9140 2143
rect -9106 2109 -9090 2143
rect -9156 2075 -9090 2109
rect -9156 2041 -9140 2075
rect -9106 2041 -9090 2075
rect -9156 2007 -9090 2041
rect -9156 1973 -9140 2007
rect -9106 1973 -9090 2007
rect -9156 1939 -9090 1973
rect -9156 1905 -9140 1939
rect -9106 1905 -9090 1939
rect -9156 1864 -9090 1905
rect -9060 2823 -8994 2864
rect -9060 2789 -9044 2823
rect -9010 2789 -8994 2823
rect -9060 2755 -8994 2789
rect -9060 2721 -9044 2755
rect -9010 2721 -8994 2755
rect -9060 2687 -8994 2721
rect -9060 2653 -9044 2687
rect -9010 2653 -8994 2687
rect -9060 2619 -8994 2653
rect -9060 2585 -9044 2619
rect -9010 2585 -8994 2619
rect -9060 2551 -8994 2585
rect -9060 2517 -9044 2551
rect -9010 2517 -8994 2551
rect -9060 2483 -8994 2517
rect -9060 2449 -9044 2483
rect -9010 2449 -8994 2483
rect -9060 2415 -8994 2449
rect -9060 2381 -9044 2415
rect -9010 2381 -8994 2415
rect -9060 2347 -8994 2381
rect -9060 2313 -9044 2347
rect -9010 2313 -8994 2347
rect -9060 2279 -8994 2313
rect -9060 2245 -9044 2279
rect -9010 2245 -8994 2279
rect -9060 2211 -8994 2245
rect -9060 2177 -9044 2211
rect -9010 2177 -8994 2211
rect -9060 2143 -8994 2177
rect -9060 2109 -9044 2143
rect -9010 2109 -8994 2143
rect -9060 2075 -8994 2109
rect -9060 2041 -9044 2075
rect -9010 2041 -8994 2075
rect -9060 2007 -8994 2041
rect -9060 1973 -9044 2007
rect -9010 1973 -8994 2007
rect -9060 1939 -8994 1973
rect -9060 1905 -9044 1939
rect -9010 1905 -8994 1939
rect -9060 1864 -8994 1905
rect -8964 2823 -8898 2864
rect -8964 2789 -8948 2823
rect -8914 2789 -8898 2823
rect -8964 2755 -8898 2789
rect -8964 2721 -8948 2755
rect -8914 2721 -8898 2755
rect -8964 2687 -8898 2721
rect -8964 2653 -8948 2687
rect -8914 2653 -8898 2687
rect -8964 2619 -8898 2653
rect -8964 2585 -8948 2619
rect -8914 2585 -8898 2619
rect -8964 2551 -8898 2585
rect -8964 2517 -8948 2551
rect -8914 2517 -8898 2551
rect -8964 2483 -8898 2517
rect -8964 2449 -8948 2483
rect -8914 2449 -8898 2483
rect -8964 2415 -8898 2449
rect -8964 2381 -8948 2415
rect -8914 2381 -8898 2415
rect -8964 2347 -8898 2381
rect -8964 2313 -8948 2347
rect -8914 2313 -8898 2347
rect -8964 2279 -8898 2313
rect -8964 2245 -8948 2279
rect -8914 2245 -8898 2279
rect -8964 2211 -8898 2245
rect -8964 2177 -8948 2211
rect -8914 2177 -8898 2211
rect -8964 2143 -8898 2177
rect -8964 2109 -8948 2143
rect -8914 2109 -8898 2143
rect -8964 2075 -8898 2109
rect -8964 2041 -8948 2075
rect -8914 2041 -8898 2075
rect -8964 2007 -8898 2041
rect -8964 1973 -8948 2007
rect -8914 1973 -8898 2007
rect -8964 1939 -8898 1973
rect -8964 1905 -8948 1939
rect -8914 1905 -8898 1939
rect -8964 1864 -8898 1905
rect -8868 2823 -8802 2864
rect -8868 2789 -8852 2823
rect -8818 2789 -8802 2823
rect -8868 2755 -8802 2789
rect -8868 2721 -8852 2755
rect -8818 2721 -8802 2755
rect -8868 2687 -8802 2721
rect -8868 2653 -8852 2687
rect -8818 2653 -8802 2687
rect -8868 2619 -8802 2653
rect -8868 2585 -8852 2619
rect -8818 2585 -8802 2619
rect -8868 2551 -8802 2585
rect -8868 2517 -8852 2551
rect -8818 2517 -8802 2551
rect -8868 2483 -8802 2517
rect -8868 2449 -8852 2483
rect -8818 2449 -8802 2483
rect -8868 2415 -8802 2449
rect -8868 2381 -8852 2415
rect -8818 2381 -8802 2415
rect -8868 2347 -8802 2381
rect -8868 2313 -8852 2347
rect -8818 2313 -8802 2347
rect -8868 2279 -8802 2313
rect -8868 2245 -8852 2279
rect -8818 2245 -8802 2279
rect -8868 2211 -8802 2245
rect -8868 2177 -8852 2211
rect -8818 2177 -8802 2211
rect -8868 2143 -8802 2177
rect -8868 2109 -8852 2143
rect -8818 2109 -8802 2143
rect -8868 2075 -8802 2109
rect -8868 2041 -8852 2075
rect -8818 2041 -8802 2075
rect -8868 2007 -8802 2041
rect -8868 1973 -8852 2007
rect -8818 1973 -8802 2007
rect -8868 1939 -8802 1973
rect -8868 1905 -8852 1939
rect -8818 1905 -8802 1939
rect -8868 1864 -8802 1905
rect -8772 2823 -8706 2864
rect -8772 2789 -8756 2823
rect -8722 2789 -8706 2823
rect -8772 2755 -8706 2789
rect -8772 2721 -8756 2755
rect -8722 2721 -8706 2755
rect -8772 2687 -8706 2721
rect -8772 2653 -8756 2687
rect -8722 2653 -8706 2687
rect -8772 2619 -8706 2653
rect -8772 2585 -8756 2619
rect -8722 2585 -8706 2619
rect -8772 2551 -8706 2585
rect -8772 2517 -8756 2551
rect -8722 2517 -8706 2551
rect -8772 2483 -8706 2517
rect -8772 2449 -8756 2483
rect -8722 2449 -8706 2483
rect -8772 2415 -8706 2449
rect -8772 2381 -8756 2415
rect -8722 2381 -8706 2415
rect -8772 2347 -8706 2381
rect -8772 2313 -8756 2347
rect -8722 2313 -8706 2347
rect -8772 2279 -8706 2313
rect -8772 2245 -8756 2279
rect -8722 2245 -8706 2279
rect -8772 2211 -8706 2245
rect -8772 2177 -8756 2211
rect -8722 2177 -8706 2211
rect -8772 2143 -8706 2177
rect -8772 2109 -8756 2143
rect -8722 2109 -8706 2143
rect -8772 2075 -8706 2109
rect -8772 2041 -8756 2075
rect -8722 2041 -8706 2075
rect -8772 2007 -8706 2041
rect -8772 1973 -8756 2007
rect -8722 1973 -8706 2007
rect -8772 1939 -8706 1973
rect -8772 1905 -8756 1939
rect -8722 1905 -8706 1939
rect -8772 1864 -8706 1905
rect -8676 2823 -8610 2864
rect -8676 2789 -8660 2823
rect -8626 2789 -8610 2823
rect -8676 2755 -8610 2789
rect -8676 2721 -8660 2755
rect -8626 2721 -8610 2755
rect -8676 2687 -8610 2721
rect -8676 2653 -8660 2687
rect -8626 2653 -8610 2687
rect -8676 2619 -8610 2653
rect -8676 2585 -8660 2619
rect -8626 2585 -8610 2619
rect -8676 2551 -8610 2585
rect -8676 2517 -8660 2551
rect -8626 2517 -8610 2551
rect -8676 2483 -8610 2517
rect -8676 2449 -8660 2483
rect -8626 2449 -8610 2483
rect -8676 2415 -8610 2449
rect -8676 2381 -8660 2415
rect -8626 2381 -8610 2415
rect -8676 2347 -8610 2381
rect -8676 2313 -8660 2347
rect -8626 2313 -8610 2347
rect -8676 2279 -8610 2313
rect -8676 2245 -8660 2279
rect -8626 2245 -8610 2279
rect -8676 2211 -8610 2245
rect -8676 2177 -8660 2211
rect -8626 2177 -8610 2211
rect -8676 2143 -8610 2177
rect -8676 2109 -8660 2143
rect -8626 2109 -8610 2143
rect -8676 2075 -8610 2109
rect -8676 2041 -8660 2075
rect -8626 2041 -8610 2075
rect -8676 2007 -8610 2041
rect -8676 1973 -8660 2007
rect -8626 1973 -8610 2007
rect -8676 1939 -8610 1973
rect -8676 1905 -8660 1939
rect -8626 1905 -8610 1939
rect -8676 1864 -8610 1905
rect -8580 2823 -8514 2864
rect -8580 2789 -8564 2823
rect -8530 2789 -8514 2823
rect -8580 2755 -8514 2789
rect -8580 2721 -8564 2755
rect -8530 2721 -8514 2755
rect -8580 2687 -8514 2721
rect -8580 2653 -8564 2687
rect -8530 2653 -8514 2687
rect -8580 2619 -8514 2653
rect -8580 2585 -8564 2619
rect -8530 2585 -8514 2619
rect -8580 2551 -8514 2585
rect -8580 2517 -8564 2551
rect -8530 2517 -8514 2551
rect -8580 2483 -8514 2517
rect -8580 2449 -8564 2483
rect -8530 2449 -8514 2483
rect -8580 2415 -8514 2449
rect -8580 2381 -8564 2415
rect -8530 2381 -8514 2415
rect -8580 2347 -8514 2381
rect -8580 2313 -8564 2347
rect -8530 2313 -8514 2347
rect -8580 2279 -8514 2313
rect -8580 2245 -8564 2279
rect -8530 2245 -8514 2279
rect -8580 2211 -8514 2245
rect -8580 2177 -8564 2211
rect -8530 2177 -8514 2211
rect -8580 2143 -8514 2177
rect -8580 2109 -8564 2143
rect -8530 2109 -8514 2143
rect -8580 2075 -8514 2109
rect -8580 2041 -8564 2075
rect -8530 2041 -8514 2075
rect -8580 2007 -8514 2041
rect -8580 1973 -8564 2007
rect -8530 1973 -8514 2007
rect -8580 1939 -8514 1973
rect -8580 1905 -8564 1939
rect -8530 1905 -8514 1939
rect -8580 1864 -8514 1905
rect -8484 2823 -8418 2864
rect -8484 2789 -8468 2823
rect -8434 2789 -8418 2823
rect -8484 2755 -8418 2789
rect -8484 2721 -8468 2755
rect -8434 2721 -8418 2755
rect -8484 2687 -8418 2721
rect -8484 2653 -8468 2687
rect -8434 2653 -8418 2687
rect -8484 2619 -8418 2653
rect -8484 2585 -8468 2619
rect -8434 2585 -8418 2619
rect -8484 2551 -8418 2585
rect -8484 2517 -8468 2551
rect -8434 2517 -8418 2551
rect -8484 2483 -8418 2517
rect -8484 2449 -8468 2483
rect -8434 2449 -8418 2483
rect -8484 2415 -8418 2449
rect -8484 2381 -8468 2415
rect -8434 2381 -8418 2415
rect -8484 2347 -8418 2381
rect -8484 2313 -8468 2347
rect -8434 2313 -8418 2347
rect -8484 2279 -8418 2313
rect -8484 2245 -8468 2279
rect -8434 2245 -8418 2279
rect -8484 2211 -8418 2245
rect -8484 2177 -8468 2211
rect -8434 2177 -8418 2211
rect -8484 2143 -8418 2177
rect -8484 2109 -8468 2143
rect -8434 2109 -8418 2143
rect -8484 2075 -8418 2109
rect -8484 2041 -8468 2075
rect -8434 2041 -8418 2075
rect -8484 2007 -8418 2041
rect -8484 1973 -8468 2007
rect -8434 1973 -8418 2007
rect -8484 1939 -8418 1973
rect -8484 1905 -8468 1939
rect -8434 1905 -8418 1939
rect -8484 1864 -8418 1905
rect -8388 2823 -8322 2864
rect -8388 2789 -8372 2823
rect -8338 2789 -8322 2823
rect -8388 2755 -8322 2789
rect -8388 2721 -8372 2755
rect -8338 2721 -8322 2755
rect -8388 2687 -8322 2721
rect -8388 2653 -8372 2687
rect -8338 2653 -8322 2687
rect -8388 2619 -8322 2653
rect -8388 2585 -8372 2619
rect -8338 2585 -8322 2619
rect -8388 2551 -8322 2585
rect -8388 2517 -8372 2551
rect -8338 2517 -8322 2551
rect -8388 2483 -8322 2517
rect -8388 2449 -8372 2483
rect -8338 2449 -8322 2483
rect -8388 2415 -8322 2449
rect -8388 2381 -8372 2415
rect -8338 2381 -8322 2415
rect -8388 2347 -8322 2381
rect -8388 2313 -8372 2347
rect -8338 2313 -8322 2347
rect -8388 2279 -8322 2313
rect -8388 2245 -8372 2279
rect -8338 2245 -8322 2279
rect -8388 2211 -8322 2245
rect -8388 2177 -8372 2211
rect -8338 2177 -8322 2211
rect -8388 2143 -8322 2177
rect -8388 2109 -8372 2143
rect -8338 2109 -8322 2143
rect -8388 2075 -8322 2109
rect -8388 2041 -8372 2075
rect -8338 2041 -8322 2075
rect -8388 2007 -8322 2041
rect -8388 1973 -8372 2007
rect -8338 1973 -8322 2007
rect -8388 1939 -8322 1973
rect -8388 1905 -8372 1939
rect -8338 1905 -8322 1939
rect -8388 1864 -8322 1905
rect -8292 2823 -8230 2864
rect -1698 2889 -1686 2923
rect -1652 2889 -1636 2923
rect -8292 2789 -8276 2823
rect -8242 2789 -8230 2823
rect -8292 2755 -8230 2789
rect -8292 2721 -8276 2755
rect -8242 2721 -8230 2755
rect -8292 2687 -8230 2721
rect -8292 2653 -8276 2687
rect -8242 2653 -8230 2687
rect -8292 2619 -8230 2653
rect -8292 2585 -8276 2619
rect -8242 2585 -8230 2619
rect -8292 2551 -8230 2585
rect -8292 2517 -8276 2551
rect -8242 2517 -8230 2551
rect -8292 2483 -8230 2517
rect -8292 2449 -8276 2483
rect -8242 2449 -8230 2483
rect -8292 2415 -8230 2449
rect -8292 2381 -8276 2415
rect -8242 2381 -8230 2415
rect -8292 2347 -8230 2381
rect -8292 2313 -8276 2347
rect -8242 2313 -8230 2347
rect -8292 2279 -8230 2313
rect -8292 2245 -8276 2279
rect -8242 2245 -8230 2279
rect -8292 2211 -8230 2245
rect -8292 2177 -8276 2211
rect -8242 2177 -8230 2211
rect -8292 2143 -8230 2177
rect -8292 2109 -8276 2143
rect -8242 2109 -8230 2143
rect -8292 2075 -8230 2109
rect -8292 2041 -8276 2075
rect -8242 2041 -8230 2075
rect -8292 2007 -8230 2041
rect -8292 1973 -8276 2007
rect -8242 1973 -8230 2007
rect -8292 1939 -8230 1973
rect -8292 1905 -8276 1939
rect -8242 1905 -8230 1939
rect -8292 1864 -8230 1905
rect -8060 2815 -7998 2856
rect -8060 2781 -8048 2815
rect -8014 2781 -7998 2815
rect -8060 2747 -7998 2781
rect -8060 2713 -8048 2747
rect -8014 2713 -7998 2747
rect -8060 2679 -7998 2713
rect -8060 2645 -8048 2679
rect -8014 2645 -7998 2679
rect -8060 2611 -7998 2645
rect -8060 2577 -8048 2611
rect -8014 2577 -7998 2611
rect -8060 2543 -7998 2577
rect -8060 2509 -8048 2543
rect -8014 2509 -7998 2543
rect -8060 2475 -7998 2509
rect -8060 2441 -8048 2475
rect -8014 2441 -7998 2475
rect -8060 2407 -7998 2441
rect -8060 2373 -8048 2407
rect -8014 2373 -7998 2407
rect -8060 2339 -7998 2373
rect -8060 2305 -8048 2339
rect -8014 2305 -7998 2339
rect -8060 2271 -7998 2305
rect -8060 2237 -8048 2271
rect -8014 2237 -7998 2271
rect -8060 2203 -7998 2237
rect -8060 2169 -8048 2203
rect -8014 2169 -7998 2203
rect -8060 2135 -7998 2169
rect -8060 2101 -8048 2135
rect -8014 2101 -7998 2135
rect -8060 2067 -7998 2101
rect -8060 2033 -8048 2067
rect -8014 2033 -7998 2067
rect -8060 1999 -7998 2033
rect -8060 1965 -8048 1999
rect -8014 1965 -7998 1999
rect -8060 1931 -7998 1965
rect -8060 1897 -8048 1931
rect -8014 1897 -7998 1931
rect -8060 1856 -7998 1897
rect -7968 2815 -7902 2856
rect -7968 2781 -7952 2815
rect -7918 2781 -7902 2815
rect -7968 2747 -7902 2781
rect -7968 2713 -7952 2747
rect -7918 2713 -7902 2747
rect -7968 2679 -7902 2713
rect -7968 2645 -7952 2679
rect -7918 2645 -7902 2679
rect -7968 2611 -7902 2645
rect -7968 2577 -7952 2611
rect -7918 2577 -7902 2611
rect -7968 2543 -7902 2577
rect -7968 2509 -7952 2543
rect -7918 2509 -7902 2543
rect -7968 2475 -7902 2509
rect -7968 2441 -7952 2475
rect -7918 2441 -7902 2475
rect -7968 2407 -7902 2441
rect -7968 2373 -7952 2407
rect -7918 2373 -7902 2407
rect -7968 2339 -7902 2373
rect -7968 2305 -7952 2339
rect -7918 2305 -7902 2339
rect -7968 2271 -7902 2305
rect -7968 2237 -7952 2271
rect -7918 2237 -7902 2271
rect -7968 2203 -7902 2237
rect -7968 2169 -7952 2203
rect -7918 2169 -7902 2203
rect -7968 2135 -7902 2169
rect -7968 2101 -7952 2135
rect -7918 2101 -7902 2135
rect -7968 2067 -7902 2101
rect -7968 2033 -7952 2067
rect -7918 2033 -7902 2067
rect -7968 1999 -7902 2033
rect -7968 1965 -7952 1999
rect -7918 1965 -7902 1999
rect -7968 1931 -7902 1965
rect -7968 1897 -7952 1931
rect -7918 1897 -7902 1931
rect -7968 1856 -7902 1897
rect -7872 2815 -7806 2856
rect -7872 2781 -7856 2815
rect -7822 2781 -7806 2815
rect -7872 2747 -7806 2781
rect -7872 2713 -7856 2747
rect -7822 2713 -7806 2747
rect -7872 2679 -7806 2713
rect -7872 2645 -7856 2679
rect -7822 2645 -7806 2679
rect -7872 2611 -7806 2645
rect -7872 2577 -7856 2611
rect -7822 2577 -7806 2611
rect -7872 2543 -7806 2577
rect -7872 2509 -7856 2543
rect -7822 2509 -7806 2543
rect -7872 2475 -7806 2509
rect -7872 2441 -7856 2475
rect -7822 2441 -7806 2475
rect -7872 2407 -7806 2441
rect -7872 2373 -7856 2407
rect -7822 2373 -7806 2407
rect -7872 2339 -7806 2373
rect -7872 2305 -7856 2339
rect -7822 2305 -7806 2339
rect -7872 2271 -7806 2305
rect -7872 2237 -7856 2271
rect -7822 2237 -7806 2271
rect -7872 2203 -7806 2237
rect -7872 2169 -7856 2203
rect -7822 2169 -7806 2203
rect -7872 2135 -7806 2169
rect -7872 2101 -7856 2135
rect -7822 2101 -7806 2135
rect -7872 2067 -7806 2101
rect -7872 2033 -7856 2067
rect -7822 2033 -7806 2067
rect -7872 1999 -7806 2033
rect -7872 1965 -7856 1999
rect -7822 1965 -7806 1999
rect -7872 1931 -7806 1965
rect -7872 1897 -7856 1931
rect -7822 1897 -7806 1931
rect -7872 1856 -7806 1897
rect -7776 2815 -7710 2856
rect -7776 2781 -7760 2815
rect -7726 2781 -7710 2815
rect -7776 2747 -7710 2781
rect -7776 2713 -7760 2747
rect -7726 2713 -7710 2747
rect -7776 2679 -7710 2713
rect -7776 2645 -7760 2679
rect -7726 2645 -7710 2679
rect -7776 2611 -7710 2645
rect -7776 2577 -7760 2611
rect -7726 2577 -7710 2611
rect -7776 2543 -7710 2577
rect -7776 2509 -7760 2543
rect -7726 2509 -7710 2543
rect -7776 2475 -7710 2509
rect -7776 2441 -7760 2475
rect -7726 2441 -7710 2475
rect -7776 2407 -7710 2441
rect -7776 2373 -7760 2407
rect -7726 2373 -7710 2407
rect -7776 2339 -7710 2373
rect -7776 2305 -7760 2339
rect -7726 2305 -7710 2339
rect -7776 2271 -7710 2305
rect -7776 2237 -7760 2271
rect -7726 2237 -7710 2271
rect -7776 2203 -7710 2237
rect -7776 2169 -7760 2203
rect -7726 2169 -7710 2203
rect -7776 2135 -7710 2169
rect -7776 2101 -7760 2135
rect -7726 2101 -7710 2135
rect -7776 2067 -7710 2101
rect -7776 2033 -7760 2067
rect -7726 2033 -7710 2067
rect -7776 1999 -7710 2033
rect -7776 1965 -7760 1999
rect -7726 1965 -7710 1999
rect -7776 1931 -7710 1965
rect -7776 1897 -7760 1931
rect -7726 1897 -7710 1931
rect -7776 1856 -7710 1897
rect -7680 2815 -7614 2856
rect -7680 2781 -7664 2815
rect -7630 2781 -7614 2815
rect -7680 2747 -7614 2781
rect -7680 2713 -7664 2747
rect -7630 2713 -7614 2747
rect -7680 2679 -7614 2713
rect -7680 2645 -7664 2679
rect -7630 2645 -7614 2679
rect -7680 2611 -7614 2645
rect -7680 2577 -7664 2611
rect -7630 2577 -7614 2611
rect -7680 2543 -7614 2577
rect -7680 2509 -7664 2543
rect -7630 2509 -7614 2543
rect -7680 2475 -7614 2509
rect -7680 2441 -7664 2475
rect -7630 2441 -7614 2475
rect -7680 2407 -7614 2441
rect -7680 2373 -7664 2407
rect -7630 2373 -7614 2407
rect -7680 2339 -7614 2373
rect -7680 2305 -7664 2339
rect -7630 2305 -7614 2339
rect -7680 2271 -7614 2305
rect -7680 2237 -7664 2271
rect -7630 2237 -7614 2271
rect -7680 2203 -7614 2237
rect -7680 2169 -7664 2203
rect -7630 2169 -7614 2203
rect -7680 2135 -7614 2169
rect -7680 2101 -7664 2135
rect -7630 2101 -7614 2135
rect -7680 2067 -7614 2101
rect -7680 2033 -7664 2067
rect -7630 2033 -7614 2067
rect -7680 1999 -7614 2033
rect -7680 1965 -7664 1999
rect -7630 1965 -7614 1999
rect -7680 1931 -7614 1965
rect -7680 1897 -7664 1931
rect -7630 1897 -7614 1931
rect -7680 1856 -7614 1897
rect -7584 2815 -7518 2856
rect -7584 2781 -7568 2815
rect -7534 2781 -7518 2815
rect -7584 2747 -7518 2781
rect -7584 2713 -7568 2747
rect -7534 2713 -7518 2747
rect -7584 2679 -7518 2713
rect -7584 2645 -7568 2679
rect -7534 2645 -7518 2679
rect -7584 2611 -7518 2645
rect -7584 2577 -7568 2611
rect -7534 2577 -7518 2611
rect -7584 2543 -7518 2577
rect -7584 2509 -7568 2543
rect -7534 2509 -7518 2543
rect -7584 2475 -7518 2509
rect -7584 2441 -7568 2475
rect -7534 2441 -7518 2475
rect -7584 2407 -7518 2441
rect -7584 2373 -7568 2407
rect -7534 2373 -7518 2407
rect -7584 2339 -7518 2373
rect -7584 2305 -7568 2339
rect -7534 2305 -7518 2339
rect -7584 2271 -7518 2305
rect -7584 2237 -7568 2271
rect -7534 2237 -7518 2271
rect -7584 2203 -7518 2237
rect -7584 2169 -7568 2203
rect -7534 2169 -7518 2203
rect -7584 2135 -7518 2169
rect -7584 2101 -7568 2135
rect -7534 2101 -7518 2135
rect -7584 2067 -7518 2101
rect -7584 2033 -7568 2067
rect -7534 2033 -7518 2067
rect -7584 1999 -7518 2033
rect -7584 1965 -7568 1999
rect -7534 1965 -7518 1999
rect -7584 1931 -7518 1965
rect -7584 1897 -7568 1931
rect -7534 1897 -7518 1931
rect -7584 1856 -7518 1897
rect -7488 2815 -7422 2856
rect -7488 2781 -7472 2815
rect -7438 2781 -7422 2815
rect -7488 2747 -7422 2781
rect -7488 2713 -7472 2747
rect -7438 2713 -7422 2747
rect -7488 2679 -7422 2713
rect -7488 2645 -7472 2679
rect -7438 2645 -7422 2679
rect -7488 2611 -7422 2645
rect -7488 2577 -7472 2611
rect -7438 2577 -7422 2611
rect -7488 2543 -7422 2577
rect -7488 2509 -7472 2543
rect -7438 2509 -7422 2543
rect -7488 2475 -7422 2509
rect -7488 2441 -7472 2475
rect -7438 2441 -7422 2475
rect -7488 2407 -7422 2441
rect -7488 2373 -7472 2407
rect -7438 2373 -7422 2407
rect -7488 2339 -7422 2373
rect -7488 2305 -7472 2339
rect -7438 2305 -7422 2339
rect -7488 2271 -7422 2305
rect -7488 2237 -7472 2271
rect -7438 2237 -7422 2271
rect -7488 2203 -7422 2237
rect -7488 2169 -7472 2203
rect -7438 2169 -7422 2203
rect -7488 2135 -7422 2169
rect -7488 2101 -7472 2135
rect -7438 2101 -7422 2135
rect -7488 2067 -7422 2101
rect -7488 2033 -7472 2067
rect -7438 2033 -7422 2067
rect -7488 1999 -7422 2033
rect -7488 1965 -7472 1999
rect -7438 1965 -7422 1999
rect -7488 1931 -7422 1965
rect -7488 1897 -7472 1931
rect -7438 1897 -7422 1931
rect -7488 1856 -7422 1897
rect -7392 2815 -7326 2856
rect -7392 2781 -7376 2815
rect -7342 2781 -7326 2815
rect -7392 2747 -7326 2781
rect -7392 2713 -7376 2747
rect -7342 2713 -7326 2747
rect -7392 2679 -7326 2713
rect -7392 2645 -7376 2679
rect -7342 2645 -7326 2679
rect -7392 2611 -7326 2645
rect -7392 2577 -7376 2611
rect -7342 2577 -7326 2611
rect -7392 2543 -7326 2577
rect -7392 2509 -7376 2543
rect -7342 2509 -7326 2543
rect -7392 2475 -7326 2509
rect -7392 2441 -7376 2475
rect -7342 2441 -7326 2475
rect -7392 2407 -7326 2441
rect -7392 2373 -7376 2407
rect -7342 2373 -7326 2407
rect -7392 2339 -7326 2373
rect -7392 2305 -7376 2339
rect -7342 2305 -7326 2339
rect -7392 2271 -7326 2305
rect -7392 2237 -7376 2271
rect -7342 2237 -7326 2271
rect -7392 2203 -7326 2237
rect -7392 2169 -7376 2203
rect -7342 2169 -7326 2203
rect -7392 2135 -7326 2169
rect -7392 2101 -7376 2135
rect -7342 2101 -7326 2135
rect -7392 2067 -7326 2101
rect -7392 2033 -7376 2067
rect -7342 2033 -7326 2067
rect -7392 1999 -7326 2033
rect -7392 1965 -7376 1999
rect -7342 1965 -7326 1999
rect -7392 1931 -7326 1965
rect -7392 1897 -7376 1931
rect -7342 1897 -7326 1931
rect -7392 1856 -7326 1897
rect -7296 2815 -7230 2856
rect -7296 2781 -7280 2815
rect -7246 2781 -7230 2815
rect -7296 2747 -7230 2781
rect -7296 2713 -7280 2747
rect -7246 2713 -7230 2747
rect -7296 2679 -7230 2713
rect -7296 2645 -7280 2679
rect -7246 2645 -7230 2679
rect -7296 2611 -7230 2645
rect -7296 2577 -7280 2611
rect -7246 2577 -7230 2611
rect -7296 2543 -7230 2577
rect -7296 2509 -7280 2543
rect -7246 2509 -7230 2543
rect -7296 2475 -7230 2509
rect -7296 2441 -7280 2475
rect -7246 2441 -7230 2475
rect -7296 2407 -7230 2441
rect -7296 2373 -7280 2407
rect -7246 2373 -7230 2407
rect -7296 2339 -7230 2373
rect -7296 2305 -7280 2339
rect -7246 2305 -7230 2339
rect -7296 2271 -7230 2305
rect -7296 2237 -7280 2271
rect -7246 2237 -7230 2271
rect -7296 2203 -7230 2237
rect -7296 2169 -7280 2203
rect -7246 2169 -7230 2203
rect -7296 2135 -7230 2169
rect -7296 2101 -7280 2135
rect -7246 2101 -7230 2135
rect -7296 2067 -7230 2101
rect -7296 2033 -7280 2067
rect -7246 2033 -7230 2067
rect -7296 1999 -7230 2033
rect -7296 1965 -7280 1999
rect -7246 1965 -7230 1999
rect -7296 1931 -7230 1965
rect -7296 1897 -7280 1931
rect -7246 1897 -7230 1931
rect -7296 1856 -7230 1897
rect -7200 2815 -7134 2856
rect -7200 2781 -7184 2815
rect -7150 2781 -7134 2815
rect -7200 2747 -7134 2781
rect -7200 2713 -7184 2747
rect -7150 2713 -7134 2747
rect -7200 2679 -7134 2713
rect -7200 2645 -7184 2679
rect -7150 2645 -7134 2679
rect -7200 2611 -7134 2645
rect -7200 2577 -7184 2611
rect -7150 2577 -7134 2611
rect -7200 2543 -7134 2577
rect -7200 2509 -7184 2543
rect -7150 2509 -7134 2543
rect -7200 2475 -7134 2509
rect -7200 2441 -7184 2475
rect -7150 2441 -7134 2475
rect -7200 2407 -7134 2441
rect -7200 2373 -7184 2407
rect -7150 2373 -7134 2407
rect -7200 2339 -7134 2373
rect -7200 2305 -7184 2339
rect -7150 2305 -7134 2339
rect -7200 2271 -7134 2305
rect -7200 2237 -7184 2271
rect -7150 2237 -7134 2271
rect -7200 2203 -7134 2237
rect -7200 2169 -7184 2203
rect -7150 2169 -7134 2203
rect -7200 2135 -7134 2169
rect -7200 2101 -7184 2135
rect -7150 2101 -7134 2135
rect -7200 2067 -7134 2101
rect -7200 2033 -7184 2067
rect -7150 2033 -7134 2067
rect -7200 1999 -7134 2033
rect -7200 1965 -7184 1999
rect -7150 1965 -7134 1999
rect -7200 1931 -7134 1965
rect -7200 1897 -7184 1931
rect -7150 1897 -7134 1931
rect -7200 1856 -7134 1897
rect -7104 2815 -7038 2856
rect -7104 2781 -7088 2815
rect -7054 2781 -7038 2815
rect -7104 2747 -7038 2781
rect -7104 2713 -7088 2747
rect -7054 2713 -7038 2747
rect -7104 2679 -7038 2713
rect -7104 2645 -7088 2679
rect -7054 2645 -7038 2679
rect -7104 2611 -7038 2645
rect -7104 2577 -7088 2611
rect -7054 2577 -7038 2611
rect -7104 2543 -7038 2577
rect -7104 2509 -7088 2543
rect -7054 2509 -7038 2543
rect -7104 2475 -7038 2509
rect -7104 2441 -7088 2475
rect -7054 2441 -7038 2475
rect -7104 2407 -7038 2441
rect -7104 2373 -7088 2407
rect -7054 2373 -7038 2407
rect -7104 2339 -7038 2373
rect -7104 2305 -7088 2339
rect -7054 2305 -7038 2339
rect -7104 2271 -7038 2305
rect -7104 2237 -7088 2271
rect -7054 2237 -7038 2271
rect -7104 2203 -7038 2237
rect -7104 2169 -7088 2203
rect -7054 2169 -7038 2203
rect -7104 2135 -7038 2169
rect -7104 2101 -7088 2135
rect -7054 2101 -7038 2135
rect -7104 2067 -7038 2101
rect -7104 2033 -7088 2067
rect -7054 2033 -7038 2067
rect -7104 1999 -7038 2033
rect -7104 1965 -7088 1999
rect -7054 1965 -7038 1999
rect -7104 1931 -7038 1965
rect -7104 1897 -7088 1931
rect -7054 1897 -7038 1931
rect -7104 1856 -7038 1897
rect -7008 2815 -6942 2856
rect -7008 2781 -6992 2815
rect -6958 2781 -6942 2815
rect -7008 2747 -6942 2781
rect -7008 2713 -6992 2747
rect -6958 2713 -6942 2747
rect -7008 2679 -6942 2713
rect -7008 2645 -6992 2679
rect -6958 2645 -6942 2679
rect -7008 2611 -6942 2645
rect -7008 2577 -6992 2611
rect -6958 2577 -6942 2611
rect -7008 2543 -6942 2577
rect -7008 2509 -6992 2543
rect -6958 2509 -6942 2543
rect -7008 2475 -6942 2509
rect -7008 2441 -6992 2475
rect -6958 2441 -6942 2475
rect -7008 2407 -6942 2441
rect -7008 2373 -6992 2407
rect -6958 2373 -6942 2407
rect -7008 2339 -6942 2373
rect -7008 2305 -6992 2339
rect -6958 2305 -6942 2339
rect -7008 2271 -6942 2305
rect -7008 2237 -6992 2271
rect -6958 2237 -6942 2271
rect -7008 2203 -6942 2237
rect -7008 2169 -6992 2203
rect -6958 2169 -6942 2203
rect -7008 2135 -6942 2169
rect -7008 2101 -6992 2135
rect -6958 2101 -6942 2135
rect -7008 2067 -6942 2101
rect -7008 2033 -6992 2067
rect -6958 2033 -6942 2067
rect -7008 1999 -6942 2033
rect -7008 1965 -6992 1999
rect -6958 1965 -6942 1999
rect -7008 1931 -6942 1965
rect -7008 1897 -6992 1931
rect -6958 1897 -6942 1931
rect -7008 1856 -6942 1897
rect -6912 2815 -6846 2856
rect -6912 2781 -6896 2815
rect -6862 2781 -6846 2815
rect -6912 2747 -6846 2781
rect -6912 2713 -6896 2747
rect -6862 2713 -6846 2747
rect -6912 2679 -6846 2713
rect -6912 2645 -6896 2679
rect -6862 2645 -6846 2679
rect -6912 2611 -6846 2645
rect -6912 2577 -6896 2611
rect -6862 2577 -6846 2611
rect -6912 2543 -6846 2577
rect -6912 2509 -6896 2543
rect -6862 2509 -6846 2543
rect -6912 2475 -6846 2509
rect -6912 2441 -6896 2475
rect -6862 2441 -6846 2475
rect -6912 2407 -6846 2441
rect -6912 2373 -6896 2407
rect -6862 2373 -6846 2407
rect -6912 2339 -6846 2373
rect -6912 2305 -6896 2339
rect -6862 2305 -6846 2339
rect -6912 2271 -6846 2305
rect -6912 2237 -6896 2271
rect -6862 2237 -6846 2271
rect -6912 2203 -6846 2237
rect -6912 2169 -6896 2203
rect -6862 2169 -6846 2203
rect -6912 2135 -6846 2169
rect -6912 2101 -6896 2135
rect -6862 2101 -6846 2135
rect -6912 2067 -6846 2101
rect -6912 2033 -6896 2067
rect -6862 2033 -6846 2067
rect -6912 1999 -6846 2033
rect -6912 1965 -6896 1999
rect -6862 1965 -6846 1999
rect -6912 1931 -6846 1965
rect -6912 1897 -6896 1931
rect -6862 1897 -6846 1931
rect -6912 1856 -6846 1897
rect -6816 2815 -6750 2856
rect -6816 2781 -6800 2815
rect -6766 2781 -6750 2815
rect -6816 2747 -6750 2781
rect -6816 2713 -6800 2747
rect -6766 2713 -6750 2747
rect -6816 2679 -6750 2713
rect -6816 2645 -6800 2679
rect -6766 2645 -6750 2679
rect -6816 2611 -6750 2645
rect -6816 2577 -6800 2611
rect -6766 2577 -6750 2611
rect -6816 2543 -6750 2577
rect -6816 2509 -6800 2543
rect -6766 2509 -6750 2543
rect -6816 2475 -6750 2509
rect -6816 2441 -6800 2475
rect -6766 2441 -6750 2475
rect -6816 2407 -6750 2441
rect -6816 2373 -6800 2407
rect -6766 2373 -6750 2407
rect -6816 2339 -6750 2373
rect -6816 2305 -6800 2339
rect -6766 2305 -6750 2339
rect -6816 2271 -6750 2305
rect -6816 2237 -6800 2271
rect -6766 2237 -6750 2271
rect -6816 2203 -6750 2237
rect -6816 2169 -6800 2203
rect -6766 2169 -6750 2203
rect -6816 2135 -6750 2169
rect -6816 2101 -6800 2135
rect -6766 2101 -6750 2135
rect -6816 2067 -6750 2101
rect -6816 2033 -6800 2067
rect -6766 2033 -6750 2067
rect -6816 1999 -6750 2033
rect -6816 1965 -6800 1999
rect -6766 1965 -6750 1999
rect -6816 1931 -6750 1965
rect -6816 1897 -6800 1931
rect -6766 1897 -6750 1931
rect -6816 1856 -6750 1897
rect -6720 2815 -6654 2856
rect -6720 2781 -6704 2815
rect -6670 2781 -6654 2815
rect -6720 2747 -6654 2781
rect -6720 2713 -6704 2747
rect -6670 2713 -6654 2747
rect -6720 2679 -6654 2713
rect -6720 2645 -6704 2679
rect -6670 2645 -6654 2679
rect -6720 2611 -6654 2645
rect -6720 2577 -6704 2611
rect -6670 2577 -6654 2611
rect -6720 2543 -6654 2577
rect -6720 2509 -6704 2543
rect -6670 2509 -6654 2543
rect -6720 2475 -6654 2509
rect -6720 2441 -6704 2475
rect -6670 2441 -6654 2475
rect -6720 2407 -6654 2441
rect -6720 2373 -6704 2407
rect -6670 2373 -6654 2407
rect -6720 2339 -6654 2373
rect -6720 2305 -6704 2339
rect -6670 2305 -6654 2339
rect -6720 2271 -6654 2305
rect -6720 2237 -6704 2271
rect -6670 2237 -6654 2271
rect -6720 2203 -6654 2237
rect -6720 2169 -6704 2203
rect -6670 2169 -6654 2203
rect -6720 2135 -6654 2169
rect -6720 2101 -6704 2135
rect -6670 2101 -6654 2135
rect -6720 2067 -6654 2101
rect -6720 2033 -6704 2067
rect -6670 2033 -6654 2067
rect -6720 1999 -6654 2033
rect -6720 1965 -6704 1999
rect -6670 1965 -6654 1999
rect -6720 1931 -6654 1965
rect -6720 1897 -6704 1931
rect -6670 1897 -6654 1931
rect -6720 1856 -6654 1897
rect -6624 2815 -6562 2856
rect -6624 2781 -6608 2815
rect -6574 2781 -6562 2815
rect -6624 2747 -6562 2781
rect -6624 2713 -6608 2747
rect -6574 2713 -6562 2747
rect -6624 2679 -6562 2713
rect -6624 2645 -6608 2679
rect -6574 2645 -6562 2679
rect -6624 2611 -6562 2645
rect -6624 2577 -6608 2611
rect -6574 2577 -6562 2611
rect -6624 2543 -6562 2577
rect -6624 2509 -6608 2543
rect -6574 2509 -6562 2543
rect -6624 2475 -6562 2509
rect -6624 2441 -6608 2475
rect -6574 2441 -6562 2475
rect -6624 2407 -6562 2441
rect -6624 2373 -6608 2407
rect -6574 2373 -6562 2407
rect -6624 2339 -6562 2373
rect -6624 2305 -6608 2339
rect -6574 2305 -6562 2339
rect -6624 2271 -6562 2305
rect -6624 2237 -6608 2271
rect -6574 2237 -6562 2271
rect -6624 2203 -6562 2237
rect -6624 2169 -6608 2203
rect -6574 2169 -6562 2203
rect -6624 2135 -6562 2169
rect -6624 2101 -6608 2135
rect -6574 2101 -6562 2135
rect -6624 2067 -6562 2101
rect -6624 2033 -6608 2067
rect -6574 2033 -6562 2067
rect -6624 1999 -6562 2033
rect -6624 1965 -6608 1999
rect -6574 1965 -6562 1999
rect -6624 1931 -6562 1965
rect -6624 1897 -6608 1931
rect -6574 1897 -6562 1931
rect -6624 1856 -6562 1897
rect -6382 2819 -6320 2860
rect -6382 2785 -6370 2819
rect -6336 2785 -6320 2819
rect -6382 2751 -6320 2785
rect -6382 2717 -6370 2751
rect -6336 2717 -6320 2751
rect -6382 2683 -6320 2717
rect -6382 2649 -6370 2683
rect -6336 2649 -6320 2683
rect -6382 2615 -6320 2649
rect -6382 2581 -6370 2615
rect -6336 2581 -6320 2615
rect -6382 2547 -6320 2581
rect -6382 2513 -6370 2547
rect -6336 2513 -6320 2547
rect -6382 2479 -6320 2513
rect -6382 2445 -6370 2479
rect -6336 2445 -6320 2479
rect -6382 2411 -6320 2445
rect -6382 2377 -6370 2411
rect -6336 2377 -6320 2411
rect -6382 2343 -6320 2377
rect -6382 2309 -6370 2343
rect -6336 2309 -6320 2343
rect -6382 2275 -6320 2309
rect -6382 2241 -6370 2275
rect -6336 2241 -6320 2275
rect -6382 2207 -6320 2241
rect -6382 2173 -6370 2207
rect -6336 2173 -6320 2207
rect -6382 2139 -6320 2173
rect -6382 2105 -6370 2139
rect -6336 2105 -6320 2139
rect -6382 2071 -6320 2105
rect -6382 2037 -6370 2071
rect -6336 2037 -6320 2071
rect -6382 2003 -6320 2037
rect -6382 1969 -6370 2003
rect -6336 1969 -6320 2003
rect -6382 1935 -6320 1969
rect -6382 1901 -6370 1935
rect -6336 1901 -6320 1935
rect -6382 1860 -6320 1901
rect -6290 2819 -6224 2860
rect -6290 2785 -6274 2819
rect -6240 2785 -6224 2819
rect -6290 2751 -6224 2785
rect -6290 2717 -6274 2751
rect -6240 2717 -6224 2751
rect -6290 2683 -6224 2717
rect -6290 2649 -6274 2683
rect -6240 2649 -6224 2683
rect -6290 2615 -6224 2649
rect -6290 2581 -6274 2615
rect -6240 2581 -6224 2615
rect -6290 2547 -6224 2581
rect -6290 2513 -6274 2547
rect -6240 2513 -6224 2547
rect -6290 2479 -6224 2513
rect -6290 2445 -6274 2479
rect -6240 2445 -6224 2479
rect -6290 2411 -6224 2445
rect -6290 2377 -6274 2411
rect -6240 2377 -6224 2411
rect -6290 2343 -6224 2377
rect -6290 2309 -6274 2343
rect -6240 2309 -6224 2343
rect -6290 2275 -6224 2309
rect -6290 2241 -6274 2275
rect -6240 2241 -6224 2275
rect -6290 2207 -6224 2241
rect -6290 2173 -6274 2207
rect -6240 2173 -6224 2207
rect -6290 2139 -6224 2173
rect -6290 2105 -6274 2139
rect -6240 2105 -6224 2139
rect -6290 2071 -6224 2105
rect -6290 2037 -6274 2071
rect -6240 2037 -6224 2071
rect -6290 2003 -6224 2037
rect -6290 1969 -6274 2003
rect -6240 1969 -6224 2003
rect -6290 1935 -6224 1969
rect -6290 1901 -6274 1935
rect -6240 1901 -6224 1935
rect -6290 1860 -6224 1901
rect -6194 2819 -6128 2860
rect -6194 2785 -6178 2819
rect -6144 2785 -6128 2819
rect -6194 2751 -6128 2785
rect -6194 2717 -6178 2751
rect -6144 2717 -6128 2751
rect -6194 2683 -6128 2717
rect -6194 2649 -6178 2683
rect -6144 2649 -6128 2683
rect -6194 2615 -6128 2649
rect -6194 2581 -6178 2615
rect -6144 2581 -6128 2615
rect -6194 2547 -6128 2581
rect -6194 2513 -6178 2547
rect -6144 2513 -6128 2547
rect -6194 2479 -6128 2513
rect -6194 2445 -6178 2479
rect -6144 2445 -6128 2479
rect -6194 2411 -6128 2445
rect -6194 2377 -6178 2411
rect -6144 2377 -6128 2411
rect -6194 2343 -6128 2377
rect -6194 2309 -6178 2343
rect -6144 2309 -6128 2343
rect -6194 2275 -6128 2309
rect -6194 2241 -6178 2275
rect -6144 2241 -6128 2275
rect -6194 2207 -6128 2241
rect -6194 2173 -6178 2207
rect -6144 2173 -6128 2207
rect -6194 2139 -6128 2173
rect -6194 2105 -6178 2139
rect -6144 2105 -6128 2139
rect -6194 2071 -6128 2105
rect -6194 2037 -6178 2071
rect -6144 2037 -6128 2071
rect -6194 2003 -6128 2037
rect -6194 1969 -6178 2003
rect -6144 1969 -6128 2003
rect -6194 1935 -6128 1969
rect -6194 1901 -6178 1935
rect -6144 1901 -6128 1935
rect -6194 1860 -6128 1901
rect -6098 2819 -6032 2860
rect -6098 2785 -6082 2819
rect -6048 2785 -6032 2819
rect -6098 2751 -6032 2785
rect -6098 2717 -6082 2751
rect -6048 2717 -6032 2751
rect -6098 2683 -6032 2717
rect -6098 2649 -6082 2683
rect -6048 2649 -6032 2683
rect -6098 2615 -6032 2649
rect -6098 2581 -6082 2615
rect -6048 2581 -6032 2615
rect -6098 2547 -6032 2581
rect -6098 2513 -6082 2547
rect -6048 2513 -6032 2547
rect -6098 2479 -6032 2513
rect -6098 2445 -6082 2479
rect -6048 2445 -6032 2479
rect -6098 2411 -6032 2445
rect -6098 2377 -6082 2411
rect -6048 2377 -6032 2411
rect -6098 2343 -6032 2377
rect -6098 2309 -6082 2343
rect -6048 2309 -6032 2343
rect -6098 2275 -6032 2309
rect -6098 2241 -6082 2275
rect -6048 2241 -6032 2275
rect -6098 2207 -6032 2241
rect -6098 2173 -6082 2207
rect -6048 2173 -6032 2207
rect -6098 2139 -6032 2173
rect -6098 2105 -6082 2139
rect -6048 2105 -6032 2139
rect -6098 2071 -6032 2105
rect -6098 2037 -6082 2071
rect -6048 2037 -6032 2071
rect -6098 2003 -6032 2037
rect -6098 1969 -6082 2003
rect -6048 1969 -6032 2003
rect -6098 1935 -6032 1969
rect -6098 1901 -6082 1935
rect -6048 1901 -6032 1935
rect -6098 1860 -6032 1901
rect -6002 2819 -5936 2860
rect -6002 2785 -5986 2819
rect -5952 2785 -5936 2819
rect -6002 2751 -5936 2785
rect -6002 2717 -5986 2751
rect -5952 2717 -5936 2751
rect -6002 2683 -5936 2717
rect -6002 2649 -5986 2683
rect -5952 2649 -5936 2683
rect -6002 2615 -5936 2649
rect -6002 2581 -5986 2615
rect -5952 2581 -5936 2615
rect -6002 2547 -5936 2581
rect -6002 2513 -5986 2547
rect -5952 2513 -5936 2547
rect -6002 2479 -5936 2513
rect -6002 2445 -5986 2479
rect -5952 2445 -5936 2479
rect -6002 2411 -5936 2445
rect -6002 2377 -5986 2411
rect -5952 2377 -5936 2411
rect -6002 2343 -5936 2377
rect -6002 2309 -5986 2343
rect -5952 2309 -5936 2343
rect -6002 2275 -5936 2309
rect -6002 2241 -5986 2275
rect -5952 2241 -5936 2275
rect -6002 2207 -5936 2241
rect -6002 2173 -5986 2207
rect -5952 2173 -5936 2207
rect -6002 2139 -5936 2173
rect -6002 2105 -5986 2139
rect -5952 2105 -5936 2139
rect -6002 2071 -5936 2105
rect -6002 2037 -5986 2071
rect -5952 2037 -5936 2071
rect -6002 2003 -5936 2037
rect -6002 1969 -5986 2003
rect -5952 1969 -5936 2003
rect -6002 1935 -5936 1969
rect -6002 1901 -5986 1935
rect -5952 1901 -5936 1935
rect -6002 1860 -5936 1901
rect -5906 2819 -5840 2860
rect -5906 2785 -5890 2819
rect -5856 2785 -5840 2819
rect -5906 2751 -5840 2785
rect -5906 2717 -5890 2751
rect -5856 2717 -5840 2751
rect -5906 2683 -5840 2717
rect -5906 2649 -5890 2683
rect -5856 2649 -5840 2683
rect -5906 2615 -5840 2649
rect -5906 2581 -5890 2615
rect -5856 2581 -5840 2615
rect -5906 2547 -5840 2581
rect -5906 2513 -5890 2547
rect -5856 2513 -5840 2547
rect -5906 2479 -5840 2513
rect -5906 2445 -5890 2479
rect -5856 2445 -5840 2479
rect -5906 2411 -5840 2445
rect -5906 2377 -5890 2411
rect -5856 2377 -5840 2411
rect -5906 2343 -5840 2377
rect -5906 2309 -5890 2343
rect -5856 2309 -5840 2343
rect -5906 2275 -5840 2309
rect -5906 2241 -5890 2275
rect -5856 2241 -5840 2275
rect -5906 2207 -5840 2241
rect -5906 2173 -5890 2207
rect -5856 2173 -5840 2207
rect -5906 2139 -5840 2173
rect -5906 2105 -5890 2139
rect -5856 2105 -5840 2139
rect -5906 2071 -5840 2105
rect -5906 2037 -5890 2071
rect -5856 2037 -5840 2071
rect -5906 2003 -5840 2037
rect -5906 1969 -5890 2003
rect -5856 1969 -5840 2003
rect -5906 1935 -5840 1969
rect -5906 1901 -5890 1935
rect -5856 1901 -5840 1935
rect -5906 1860 -5840 1901
rect -5810 2819 -5744 2860
rect -5810 2785 -5794 2819
rect -5760 2785 -5744 2819
rect -5810 2751 -5744 2785
rect -5810 2717 -5794 2751
rect -5760 2717 -5744 2751
rect -5810 2683 -5744 2717
rect -5810 2649 -5794 2683
rect -5760 2649 -5744 2683
rect -5810 2615 -5744 2649
rect -5810 2581 -5794 2615
rect -5760 2581 -5744 2615
rect -5810 2547 -5744 2581
rect -5810 2513 -5794 2547
rect -5760 2513 -5744 2547
rect -5810 2479 -5744 2513
rect -5810 2445 -5794 2479
rect -5760 2445 -5744 2479
rect -5810 2411 -5744 2445
rect -5810 2377 -5794 2411
rect -5760 2377 -5744 2411
rect -5810 2343 -5744 2377
rect -5810 2309 -5794 2343
rect -5760 2309 -5744 2343
rect -5810 2275 -5744 2309
rect -5810 2241 -5794 2275
rect -5760 2241 -5744 2275
rect -5810 2207 -5744 2241
rect -5810 2173 -5794 2207
rect -5760 2173 -5744 2207
rect -5810 2139 -5744 2173
rect -5810 2105 -5794 2139
rect -5760 2105 -5744 2139
rect -5810 2071 -5744 2105
rect -5810 2037 -5794 2071
rect -5760 2037 -5744 2071
rect -5810 2003 -5744 2037
rect -5810 1969 -5794 2003
rect -5760 1969 -5744 2003
rect -5810 1935 -5744 1969
rect -5810 1901 -5794 1935
rect -5760 1901 -5744 1935
rect -5810 1860 -5744 1901
rect -5714 2819 -5648 2860
rect -5714 2785 -5698 2819
rect -5664 2785 -5648 2819
rect -5714 2751 -5648 2785
rect -5714 2717 -5698 2751
rect -5664 2717 -5648 2751
rect -5714 2683 -5648 2717
rect -5714 2649 -5698 2683
rect -5664 2649 -5648 2683
rect -5714 2615 -5648 2649
rect -5714 2581 -5698 2615
rect -5664 2581 -5648 2615
rect -5714 2547 -5648 2581
rect -5714 2513 -5698 2547
rect -5664 2513 -5648 2547
rect -5714 2479 -5648 2513
rect -5714 2445 -5698 2479
rect -5664 2445 -5648 2479
rect -5714 2411 -5648 2445
rect -5714 2377 -5698 2411
rect -5664 2377 -5648 2411
rect -5714 2343 -5648 2377
rect -5714 2309 -5698 2343
rect -5664 2309 -5648 2343
rect -5714 2275 -5648 2309
rect -5714 2241 -5698 2275
rect -5664 2241 -5648 2275
rect -5714 2207 -5648 2241
rect -5714 2173 -5698 2207
rect -5664 2173 -5648 2207
rect -5714 2139 -5648 2173
rect -5714 2105 -5698 2139
rect -5664 2105 -5648 2139
rect -5714 2071 -5648 2105
rect -5714 2037 -5698 2071
rect -5664 2037 -5648 2071
rect -5714 2003 -5648 2037
rect -5714 1969 -5698 2003
rect -5664 1969 -5648 2003
rect -5714 1935 -5648 1969
rect -5714 1901 -5698 1935
rect -5664 1901 -5648 1935
rect -5714 1860 -5648 1901
rect -5618 2819 -5552 2860
rect -5618 2785 -5602 2819
rect -5568 2785 -5552 2819
rect -5618 2751 -5552 2785
rect -5618 2717 -5602 2751
rect -5568 2717 -5552 2751
rect -5618 2683 -5552 2717
rect -5618 2649 -5602 2683
rect -5568 2649 -5552 2683
rect -5618 2615 -5552 2649
rect -5618 2581 -5602 2615
rect -5568 2581 -5552 2615
rect -5618 2547 -5552 2581
rect -5618 2513 -5602 2547
rect -5568 2513 -5552 2547
rect -5618 2479 -5552 2513
rect -5618 2445 -5602 2479
rect -5568 2445 -5552 2479
rect -5618 2411 -5552 2445
rect -5618 2377 -5602 2411
rect -5568 2377 -5552 2411
rect -5618 2343 -5552 2377
rect -5618 2309 -5602 2343
rect -5568 2309 -5552 2343
rect -5618 2275 -5552 2309
rect -5618 2241 -5602 2275
rect -5568 2241 -5552 2275
rect -5618 2207 -5552 2241
rect -5618 2173 -5602 2207
rect -5568 2173 -5552 2207
rect -5618 2139 -5552 2173
rect -5618 2105 -5602 2139
rect -5568 2105 -5552 2139
rect -5618 2071 -5552 2105
rect -5618 2037 -5602 2071
rect -5568 2037 -5552 2071
rect -5618 2003 -5552 2037
rect -5618 1969 -5602 2003
rect -5568 1969 -5552 2003
rect -5618 1935 -5552 1969
rect -5618 1901 -5602 1935
rect -5568 1901 -5552 1935
rect -5618 1860 -5552 1901
rect -5522 2819 -5456 2860
rect -5522 2785 -5506 2819
rect -5472 2785 -5456 2819
rect -5522 2751 -5456 2785
rect -5522 2717 -5506 2751
rect -5472 2717 -5456 2751
rect -5522 2683 -5456 2717
rect -5522 2649 -5506 2683
rect -5472 2649 -5456 2683
rect -5522 2615 -5456 2649
rect -5522 2581 -5506 2615
rect -5472 2581 -5456 2615
rect -5522 2547 -5456 2581
rect -5522 2513 -5506 2547
rect -5472 2513 -5456 2547
rect -5522 2479 -5456 2513
rect -5522 2445 -5506 2479
rect -5472 2445 -5456 2479
rect -5522 2411 -5456 2445
rect -5522 2377 -5506 2411
rect -5472 2377 -5456 2411
rect -5522 2343 -5456 2377
rect -5522 2309 -5506 2343
rect -5472 2309 -5456 2343
rect -5522 2275 -5456 2309
rect -5522 2241 -5506 2275
rect -5472 2241 -5456 2275
rect -5522 2207 -5456 2241
rect -5522 2173 -5506 2207
rect -5472 2173 -5456 2207
rect -5522 2139 -5456 2173
rect -5522 2105 -5506 2139
rect -5472 2105 -5456 2139
rect -5522 2071 -5456 2105
rect -5522 2037 -5506 2071
rect -5472 2037 -5456 2071
rect -5522 2003 -5456 2037
rect -5522 1969 -5506 2003
rect -5472 1969 -5456 2003
rect -5522 1935 -5456 1969
rect -5522 1901 -5506 1935
rect -5472 1901 -5456 1935
rect -5522 1860 -5456 1901
rect -5426 2819 -5364 2860
rect -5426 2785 -5410 2819
rect -5376 2785 -5364 2819
rect -5426 2751 -5364 2785
rect -5426 2717 -5410 2751
rect -5376 2717 -5364 2751
rect -5426 2683 -5364 2717
rect -5426 2649 -5410 2683
rect -5376 2649 -5364 2683
rect -5426 2615 -5364 2649
rect -5426 2581 -5410 2615
rect -5376 2581 -5364 2615
rect -5426 2547 -5364 2581
rect -5426 2513 -5410 2547
rect -5376 2513 -5364 2547
rect -5426 2479 -5364 2513
rect -5426 2445 -5410 2479
rect -5376 2445 -5364 2479
rect -5426 2411 -5364 2445
rect -5426 2377 -5410 2411
rect -5376 2377 -5364 2411
rect -5426 2343 -5364 2377
rect -5426 2309 -5410 2343
rect -5376 2309 -5364 2343
rect -5426 2275 -5364 2309
rect -5426 2241 -5410 2275
rect -5376 2241 -5364 2275
rect -5426 2207 -5364 2241
rect -5426 2173 -5410 2207
rect -5376 2173 -5364 2207
rect -5426 2139 -5364 2173
rect -5426 2105 -5410 2139
rect -5376 2105 -5364 2139
rect -5426 2071 -5364 2105
rect -5426 2037 -5410 2071
rect -5376 2037 -5364 2071
rect -5426 2003 -5364 2037
rect -5426 1969 -5410 2003
rect -5376 1969 -5364 2003
rect -5426 1935 -5364 1969
rect -5426 1901 -5410 1935
rect -5376 1901 -5364 1935
rect -5426 1860 -5364 1901
rect -5210 2829 -5148 2870
rect -5210 2795 -5198 2829
rect -5164 2795 -5148 2829
rect -5210 2761 -5148 2795
rect -5210 2727 -5198 2761
rect -5164 2727 -5148 2761
rect -5210 2693 -5148 2727
rect -5210 2659 -5198 2693
rect -5164 2659 -5148 2693
rect -5210 2625 -5148 2659
rect -5210 2591 -5198 2625
rect -5164 2591 -5148 2625
rect -5210 2557 -5148 2591
rect -5210 2523 -5198 2557
rect -5164 2523 -5148 2557
rect -5210 2489 -5148 2523
rect -5210 2455 -5198 2489
rect -5164 2455 -5148 2489
rect -5210 2421 -5148 2455
rect -5210 2387 -5198 2421
rect -5164 2387 -5148 2421
rect -5210 2353 -5148 2387
rect -5210 2319 -5198 2353
rect -5164 2319 -5148 2353
rect -5210 2285 -5148 2319
rect -5210 2251 -5198 2285
rect -5164 2251 -5148 2285
rect -5210 2217 -5148 2251
rect -5210 2183 -5198 2217
rect -5164 2183 -5148 2217
rect -5210 2149 -5148 2183
rect -5210 2115 -5198 2149
rect -5164 2115 -5148 2149
rect -5210 2081 -5148 2115
rect -5210 2047 -5198 2081
rect -5164 2047 -5148 2081
rect -5210 2013 -5148 2047
rect -5210 1979 -5198 2013
rect -5164 1979 -5148 2013
rect -5210 1945 -5148 1979
rect -5210 1911 -5198 1945
rect -5164 1911 -5148 1945
rect -5210 1870 -5148 1911
rect -5118 2829 -5052 2870
rect -5118 2795 -5102 2829
rect -5068 2795 -5052 2829
rect -5118 2761 -5052 2795
rect -5118 2727 -5102 2761
rect -5068 2727 -5052 2761
rect -5118 2693 -5052 2727
rect -5118 2659 -5102 2693
rect -5068 2659 -5052 2693
rect -5118 2625 -5052 2659
rect -5118 2591 -5102 2625
rect -5068 2591 -5052 2625
rect -5118 2557 -5052 2591
rect -5118 2523 -5102 2557
rect -5068 2523 -5052 2557
rect -5118 2489 -5052 2523
rect -5118 2455 -5102 2489
rect -5068 2455 -5052 2489
rect -5118 2421 -5052 2455
rect -5118 2387 -5102 2421
rect -5068 2387 -5052 2421
rect -5118 2353 -5052 2387
rect -5118 2319 -5102 2353
rect -5068 2319 -5052 2353
rect -5118 2285 -5052 2319
rect -5118 2251 -5102 2285
rect -5068 2251 -5052 2285
rect -5118 2217 -5052 2251
rect -5118 2183 -5102 2217
rect -5068 2183 -5052 2217
rect -5118 2149 -5052 2183
rect -5118 2115 -5102 2149
rect -5068 2115 -5052 2149
rect -5118 2081 -5052 2115
rect -5118 2047 -5102 2081
rect -5068 2047 -5052 2081
rect -5118 2013 -5052 2047
rect -5118 1979 -5102 2013
rect -5068 1979 -5052 2013
rect -5118 1945 -5052 1979
rect -5118 1911 -5102 1945
rect -5068 1911 -5052 1945
rect -5118 1870 -5052 1911
rect -5022 2829 -4956 2870
rect -5022 2795 -5006 2829
rect -4972 2795 -4956 2829
rect -5022 2761 -4956 2795
rect -5022 2727 -5006 2761
rect -4972 2727 -4956 2761
rect -5022 2693 -4956 2727
rect -5022 2659 -5006 2693
rect -4972 2659 -4956 2693
rect -5022 2625 -4956 2659
rect -5022 2591 -5006 2625
rect -4972 2591 -4956 2625
rect -5022 2557 -4956 2591
rect -5022 2523 -5006 2557
rect -4972 2523 -4956 2557
rect -5022 2489 -4956 2523
rect -5022 2455 -5006 2489
rect -4972 2455 -4956 2489
rect -5022 2421 -4956 2455
rect -5022 2387 -5006 2421
rect -4972 2387 -4956 2421
rect -5022 2353 -4956 2387
rect -5022 2319 -5006 2353
rect -4972 2319 -4956 2353
rect -5022 2285 -4956 2319
rect -5022 2251 -5006 2285
rect -4972 2251 -4956 2285
rect -5022 2217 -4956 2251
rect -5022 2183 -5006 2217
rect -4972 2183 -4956 2217
rect -5022 2149 -4956 2183
rect -5022 2115 -5006 2149
rect -4972 2115 -4956 2149
rect -5022 2081 -4956 2115
rect -5022 2047 -5006 2081
rect -4972 2047 -4956 2081
rect -5022 2013 -4956 2047
rect -5022 1979 -5006 2013
rect -4972 1979 -4956 2013
rect -5022 1945 -4956 1979
rect -5022 1911 -5006 1945
rect -4972 1911 -4956 1945
rect -5022 1870 -4956 1911
rect -4926 2829 -4860 2870
rect -4926 2795 -4910 2829
rect -4876 2795 -4860 2829
rect -4926 2761 -4860 2795
rect -4926 2727 -4910 2761
rect -4876 2727 -4860 2761
rect -4926 2693 -4860 2727
rect -4926 2659 -4910 2693
rect -4876 2659 -4860 2693
rect -4926 2625 -4860 2659
rect -4926 2591 -4910 2625
rect -4876 2591 -4860 2625
rect -4926 2557 -4860 2591
rect -4926 2523 -4910 2557
rect -4876 2523 -4860 2557
rect -4926 2489 -4860 2523
rect -4926 2455 -4910 2489
rect -4876 2455 -4860 2489
rect -4926 2421 -4860 2455
rect -4926 2387 -4910 2421
rect -4876 2387 -4860 2421
rect -4926 2353 -4860 2387
rect -4926 2319 -4910 2353
rect -4876 2319 -4860 2353
rect -4926 2285 -4860 2319
rect -4926 2251 -4910 2285
rect -4876 2251 -4860 2285
rect -4926 2217 -4860 2251
rect -4926 2183 -4910 2217
rect -4876 2183 -4860 2217
rect -4926 2149 -4860 2183
rect -4926 2115 -4910 2149
rect -4876 2115 -4860 2149
rect -4926 2081 -4860 2115
rect -4926 2047 -4910 2081
rect -4876 2047 -4860 2081
rect -4926 2013 -4860 2047
rect -4926 1979 -4910 2013
rect -4876 1979 -4860 2013
rect -4926 1945 -4860 1979
rect -4926 1911 -4910 1945
rect -4876 1911 -4860 1945
rect -4926 1870 -4860 1911
rect -4830 2829 -4764 2870
rect -4830 2795 -4814 2829
rect -4780 2795 -4764 2829
rect -4830 2761 -4764 2795
rect -4830 2727 -4814 2761
rect -4780 2727 -4764 2761
rect -4830 2693 -4764 2727
rect -4830 2659 -4814 2693
rect -4780 2659 -4764 2693
rect -4830 2625 -4764 2659
rect -4830 2591 -4814 2625
rect -4780 2591 -4764 2625
rect -4830 2557 -4764 2591
rect -4830 2523 -4814 2557
rect -4780 2523 -4764 2557
rect -4830 2489 -4764 2523
rect -4830 2455 -4814 2489
rect -4780 2455 -4764 2489
rect -4830 2421 -4764 2455
rect -4830 2387 -4814 2421
rect -4780 2387 -4764 2421
rect -4830 2353 -4764 2387
rect -4830 2319 -4814 2353
rect -4780 2319 -4764 2353
rect -4830 2285 -4764 2319
rect -4830 2251 -4814 2285
rect -4780 2251 -4764 2285
rect -4830 2217 -4764 2251
rect -4830 2183 -4814 2217
rect -4780 2183 -4764 2217
rect -4830 2149 -4764 2183
rect -4830 2115 -4814 2149
rect -4780 2115 -4764 2149
rect -4830 2081 -4764 2115
rect -4830 2047 -4814 2081
rect -4780 2047 -4764 2081
rect -4830 2013 -4764 2047
rect -4830 1979 -4814 2013
rect -4780 1979 -4764 2013
rect -4830 1945 -4764 1979
rect -4830 1911 -4814 1945
rect -4780 1911 -4764 1945
rect -4830 1870 -4764 1911
rect -4734 2829 -4672 2870
rect -4734 2795 -4718 2829
rect -4684 2795 -4672 2829
rect -4734 2761 -4672 2795
rect -4734 2727 -4718 2761
rect -4684 2727 -4672 2761
rect -4734 2693 -4672 2727
rect -4734 2659 -4718 2693
rect -4684 2659 -4672 2693
rect -4734 2625 -4672 2659
rect -4734 2591 -4718 2625
rect -4684 2591 -4672 2625
rect -4734 2557 -4672 2591
rect -4734 2523 -4718 2557
rect -4684 2523 -4672 2557
rect -4734 2489 -4672 2523
rect -4734 2455 -4718 2489
rect -4684 2455 -4672 2489
rect -4734 2421 -4672 2455
rect -4734 2387 -4718 2421
rect -4684 2387 -4672 2421
rect -4734 2353 -4672 2387
rect -4734 2319 -4718 2353
rect -4684 2319 -4672 2353
rect -4734 2285 -4672 2319
rect -4734 2251 -4718 2285
rect -4684 2251 -4672 2285
rect -4734 2217 -4672 2251
rect -1698 2855 -1636 2889
rect -1698 2821 -1686 2855
rect -1652 2821 -1636 2855
rect -1698 2787 -1636 2821
rect -1698 2753 -1686 2787
rect -1652 2753 -1636 2787
rect -1698 2719 -1636 2753
rect -1698 2685 -1686 2719
rect -1652 2685 -1636 2719
rect -1698 2651 -1636 2685
rect -1698 2617 -1686 2651
rect -1652 2617 -1636 2651
rect -1698 2583 -1636 2617
rect -1698 2549 -1686 2583
rect -1652 2549 -1636 2583
rect -1698 2515 -1636 2549
rect -1698 2481 -1686 2515
rect -1652 2481 -1636 2515
rect -1698 2447 -1636 2481
rect -1698 2413 -1686 2447
rect -1652 2413 -1636 2447
rect -1698 2379 -1636 2413
rect -1698 2345 -1686 2379
rect -1652 2345 -1636 2379
rect -1698 2311 -1636 2345
rect -1698 2277 -1686 2311
rect -1652 2277 -1636 2311
rect -1698 2236 -1636 2277
rect -1606 3195 -1540 3236
rect -1606 3161 -1590 3195
rect -1556 3161 -1540 3195
rect -1606 3127 -1540 3161
rect -1606 3093 -1590 3127
rect -1556 3093 -1540 3127
rect -1606 3059 -1540 3093
rect -1606 3025 -1590 3059
rect -1556 3025 -1540 3059
rect -1606 2991 -1540 3025
rect -1606 2957 -1590 2991
rect -1556 2957 -1540 2991
rect -1606 2923 -1540 2957
rect -1606 2889 -1590 2923
rect -1556 2889 -1540 2923
rect -1606 2855 -1540 2889
rect -1606 2821 -1590 2855
rect -1556 2821 -1540 2855
rect -1606 2787 -1540 2821
rect -1606 2753 -1590 2787
rect -1556 2753 -1540 2787
rect -1606 2719 -1540 2753
rect -1606 2685 -1590 2719
rect -1556 2685 -1540 2719
rect -1606 2651 -1540 2685
rect -1606 2617 -1590 2651
rect -1556 2617 -1540 2651
rect -1606 2583 -1540 2617
rect -1606 2549 -1590 2583
rect -1556 2549 -1540 2583
rect -1606 2515 -1540 2549
rect -1606 2481 -1590 2515
rect -1556 2481 -1540 2515
rect -1606 2447 -1540 2481
rect -1606 2413 -1590 2447
rect -1556 2413 -1540 2447
rect -1606 2379 -1540 2413
rect -1606 2345 -1590 2379
rect -1556 2345 -1540 2379
rect -1606 2311 -1540 2345
rect -1606 2277 -1590 2311
rect -1556 2277 -1540 2311
rect -1606 2236 -1540 2277
rect -1510 3195 -1444 3236
rect -1510 3161 -1494 3195
rect -1460 3161 -1444 3195
rect -1510 3127 -1444 3161
rect -1510 3093 -1494 3127
rect -1460 3093 -1444 3127
rect -1510 3059 -1444 3093
rect -1510 3025 -1494 3059
rect -1460 3025 -1444 3059
rect -1510 2991 -1444 3025
rect -1510 2957 -1494 2991
rect -1460 2957 -1444 2991
rect -1510 2923 -1444 2957
rect -1510 2889 -1494 2923
rect -1460 2889 -1444 2923
rect -1510 2855 -1444 2889
rect -1510 2821 -1494 2855
rect -1460 2821 -1444 2855
rect -1510 2787 -1444 2821
rect -1510 2753 -1494 2787
rect -1460 2753 -1444 2787
rect -1510 2719 -1444 2753
rect -1510 2685 -1494 2719
rect -1460 2685 -1444 2719
rect -1510 2651 -1444 2685
rect -1510 2617 -1494 2651
rect -1460 2617 -1444 2651
rect -1510 2583 -1444 2617
rect -1510 2549 -1494 2583
rect -1460 2549 -1444 2583
rect -1510 2515 -1444 2549
rect -1510 2481 -1494 2515
rect -1460 2481 -1444 2515
rect -1510 2447 -1444 2481
rect -1510 2413 -1494 2447
rect -1460 2413 -1444 2447
rect -1510 2379 -1444 2413
rect -1510 2345 -1494 2379
rect -1460 2345 -1444 2379
rect -1510 2311 -1444 2345
rect -1510 2277 -1494 2311
rect -1460 2277 -1444 2311
rect -1510 2236 -1444 2277
rect -1414 3195 -1348 3236
rect -1414 3161 -1398 3195
rect -1364 3161 -1348 3195
rect -1414 3127 -1348 3161
rect -1414 3093 -1398 3127
rect -1364 3093 -1348 3127
rect -1414 3059 -1348 3093
rect -1414 3025 -1398 3059
rect -1364 3025 -1348 3059
rect -1414 2991 -1348 3025
rect -1414 2957 -1398 2991
rect -1364 2957 -1348 2991
rect -1414 2923 -1348 2957
rect -1414 2889 -1398 2923
rect -1364 2889 -1348 2923
rect -1414 2855 -1348 2889
rect -1414 2821 -1398 2855
rect -1364 2821 -1348 2855
rect -1414 2787 -1348 2821
rect -1414 2753 -1398 2787
rect -1364 2753 -1348 2787
rect -1414 2719 -1348 2753
rect -1414 2685 -1398 2719
rect -1364 2685 -1348 2719
rect -1414 2651 -1348 2685
rect -1414 2617 -1398 2651
rect -1364 2617 -1348 2651
rect -1414 2583 -1348 2617
rect -1414 2549 -1398 2583
rect -1364 2549 -1348 2583
rect -1414 2515 -1348 2549
rect -1414 2481 -1398 2515
rect -1364 2481 -1348 2515
rect -1414 2447 -1348 2481
rect -1414 2413 -1398 2447
rect -1364 2413 -1348 2447
rect -1414 2379 -1348 2413
rect -1414 2345 -1398 2379
rect -1364 2345 -1348 2379
rect -1414 2311 -1348 2345
rect -1414 2277 -1398 2311
rect -1364 2277 -1348 2311
rect -1414 2236 -1348 2277
rect -1318 3195 -1252 3236
rect -1318 3161 -1302 3195
rect -1268 3161 -1252 3195
rect -1318 3127 -1252 3161
rect -1318 3093 -1302 3127
rect -1268 3093 -1252 3127
rect -1318 3059 -1252 3093
rect -1318 3025 -1302 3059
rect -1268 3025 -1252 3059
rect -1318 2991 -1252 3025
rect -1318 2957 -1302 2991
rect -1268 2957 -1252 2991
rect -1318 2923 -1252 2957
rect -1318 2889 -1302 2923
rect -1268 2889 -1252 2923
rect -1318 2855 -1252 2889
rect -1318 2821 -1302 2855
rect -1268 2821 -1252 2855
rect -1318 2787 -1252 2821
rect -1318 2753 -1302 2787
rect -1268 2753 -1252 2787
rect -1318 2719 -1252 2753
rect -1318 2685 -1302 2719
rect -1268 2685 -1252 2719
rect -1318 2651 -1252 2685
rect -1318 2617 -1302 2651
rect -1268 2617 -1252 2651
rect -1318 2583 -1252 2617
rect -1318 2549 -1302 2583
rect -1268 2549 -1252 2583
rect -1318 2515 -1252 2549
rect -1318 2481 -1302 2515
rect -1268 2481 -1252 2515
rect -1318 2447 -1252 2481
rect -1318 2413 -1302 2447
rect -1268 2413 -1252 2447
rect -1318 2379 -1252 2413
rect -1318 2345 -1302 2379
rect -1268 2345 -1252 2379
rect -1318 2311 -1252 2345
rect -1318 2277 -1302 2311
rect -1268 2277 -1252 2311
rect -1318 2236 -1252 2277
rect -1222 3195 -1156 3236
rect -1222 3161 -1206 3195
rect -1172 3161 -1156 3195
rect -1222 3127 -1156 3161
rect -1222 3093 -1206 3127
rect -1172 3093 -1156 3127
rect -1222 3059 -1156 3093
rect -1222 3025 -1206 3059
rect -1172 3025 -1156 3059
rect -1222 2991 -1156 3025
rect -1222 2957 -1206 2991
rect -1172 2957 -1156 2991
rect -1222 2923 -1156 2957
rect -1222 2889 -1206 2923
rect -1172 2889 -1156 2923
rect -1222 2855 -1156 2889
rect -1222 2821 -1206 2855
rect -1172 2821 -1156 2855
rect -1222 2787 -1156 2821
rect -1222 2753 -1206 2787
rect -1172 2753 -1156 2787
rect -1222 2719 -1156 2753
rect -1222 2685 -1206 2719
rect -1172 2685 -1156 2719
rect -1222 2651 -1156 2685
rect -1222 2617 -1206 2651
rect -1172 2617 -1156 2651
rect -1222 2583 -1156 2617
rect -1222 2549 -1206 2583
rect -1172 2549 -1156 2583
rect -1222 2515 -1156 2549
rect -1222 2481 -1206 2515
rect -1172 2481 -1156 2515
rect -1222 2447 -1156 2481
rect -1222 2413 -1206 2447
rect -1172 2413 -1156 2447
rect -1222 2379 -1156 2413
rect -1222 2345 -1206 2379
rect -1172 2345 -1156 2379
rect -1222 2311 -1156 2345
rect -1222 2277 -1206 2311
rect -1172 2277 -1156 2311
rect -1222 2236 -1156 2277
rect -1126 3195 -1060 3236
rect -1126 3161 -1110 3195
rect -1076 3161 -1060 3195
rect -1126 3127 -1060 3161
rect -1126 3093 -1110 3127
rect -1076 3093 -1060 3127
rect -1126 3059 -1060 3093
rect -1126 3025 -1110 3059
rect -1076 3025 -1060 3059
rect -1126 2991 -1060 3025
rect -1126 2957 -1110 2991
rect -1076 2957 -1060 2991
rect -1126 2923 -1060 2957
rect -1126 2889 -1110 2923
rect -1076 2889 -1060 2923
rect -1126 2855 -1060 2889
rect -1126 2821 -1110 2855
rect -1076 2821 -1060 2855
rect -1126 2787 -1060 2821
rect -1126 2753 -1110 2787
rect -1076 2753 -1060 2787
rect -1126 2719 -1060 2753
rect -1126 2685 -1110 2719
rect -1076 2685 -1060 2719
rect -1126 2651 -1060 2685
rect -1126 2617 -1110 2651
rect -1076 2617 -1060 2651
rect -1126 2583 -1060 2617
rect -1126 2549 -1110 2583
rect -1076 2549 -1060 2583
rect -1126 2515 -1060 2549
rect -1126 2481 -1110 2515
rect -1076 2481 -1060 2515
rect -1126 2447 -1060 2481
rect -1126 2413 -1110 2447
rect -1076 2413 -1060 2447
rect -1126 2379 -1060 2413
rect -1126 2345 -1110 2379
rect -1076 2345 -1060 2379
rect -1126 2311 -1060 2345
rect -1126 2277 -1110 2311
rect -1076 2277 -1060 2311
rect -1126 2236 -1060 2277
rect -1030 3195 -964 3236
rect -1030 3161 -1014 3195
rect -980 3161 -964 3195
rect -1030 3127 -964 3161
rect -1030 3093 -1014 3127
rect -980 3093 -964 3127
rect -1030 3059 -964 3093
rect -1030 3025 -1014 3059
rect -980 3025 -964 3059
rect -1030 2991 -964 3025
rect -1030 2957 -1014 2991
rect -980 2957 -964 2991
rect -1030 2923 -964 2957
rect -1030 2889 -1014 2923
rect -980 2889 -964 2923
rect -1030 2855 -964 2889
rect -1030 2821 -1014 2855
rect -980 2821 -964 2855
rect -1030 2787 -964 2821
rect -1030 2753 -1014 2787
rect -980 2753 -964 2787
rect -1030 2719 -964 2753
rect -1030 2685 -1014 2719
rect -980 2685 -964 2719
rect -1030 2651 -964 2685
rect -1030 2617 -1014 2651
rect -980 2617 -964 2651
rect -1030 2583 -964 2617
rect -1030 2549 -1014 2583
rect -980 2549 -964 2583
rect -1030 2515 -964 2549
rect -1030 2481 -1014 2515
rect -980 2481 -964 2515
rect -1030 2447 -964 2481
rect -1030 2413 -1014 2447
rect -980 2413 -964 2447
rect -1030 2379 -964 2413
rect -1030 2345 -1014 2379
rect -980 2345 -964 2379
rect -1030 2311 -964 2345
rect -1030 2277 -1014 2311
rect -980 2277 -964 2311
rect -1030 2236 -964 2277
rect -934 3195 -872 3236
rect -934 3161 -918 3195
rect -884 3161 -872 3195
rect -934 3127 -872 3161
rect -934 3093 -918 3127
rect -884 3093 -872 3127
rect -934 3059 -872 3093
rect -934 3025 -918 3059
rect -884 3025 -872 3059
rect -934 2991 -872 3025
rect 16674 3221 16736 3255
rect 16674 3187 16686 3221
rect 16720 3187 16736 3221
rect 16674 3153 16736 3187
rect 16674 3119 16686 3153
rect 16720 3119 16736 3153
rect 16674 3085 16736 3119
rect 16674 3051 16686 3085
rect 16720 3051 16736 3085
rect -934 2957 -918 2991
rect -884 2957 -872 2991
rect -934 2923 -872 2957
rect 16674 3017 16736 3051
rect -934 2889 -918 2923
rect -884 2889 -872 2923
rect 16674 2983 16686 3017
rect 16720 2983 16736 3017
rect -934 2855 -872 2889
rect -934 2821 -918 2855
rect -884 2821 -872 2855
rect -934 2787 -872 2821
rect -934 2753 -918 2787
rect -884 2753 -872 2787
rect -934 2719 -872 2753
rect -934 2685 -918 2719
rect -884 2685 -872 2719
rect -934 2651 -872 2685
rect -934 2617 -918 2651
rect -884 2617 -872 2651
rect -934 2583 -872 2617
rect -934 2549 -918 2583
rect -884 2549 -872 2583
rect -934 2515 -872 2549
rect -934 2481 -918 2515
rect -884 2481 -872 2515
rect -934 2447 -872 2481
rect -934 2413 -918 2447
rect -884 2413 -872 2447
rect -934 2379 -872 2413
rect -934 2345 -918 2379
rect -884 2345 -872 2379
rect -934 2311 -872 2345
rect -934 2277 -918 2311
rect -884 2277 -872 2311
rect -934 2236 -872 2277
rect 1470 2789 1532 2830
rect 1470 2755 1482 2789
rect 1516 2755 1532 2789
rect 1470 2721 1532 2755
rect 1470 2687 1482 2721
rect 1516 2687 1532 2721
rect 1470 2653 1532 2687
rect 1470 2619 1482 2653
rect 1516 2619 1532 2653
rect 1470 2585 1532 2619
rect 1470 2551 1482 2585
rect 1516 2551 1532 2585
rect 1470 2517 1532 2551
rect 1470 2483 1482 2517
rect 1516 2483 1532 2517
rect 1470 2449 1532 2483
rect 1470 2415 1482 2449
rect 1516 2415 1532 2449
rect 1470 2381 1532 2415
rect 1470 2347 1482 2381
rect 1516 2347 1532 2381
rect 1470 2313 1532 2347
rect 1470 2279 1482 2313
rect 1516 2279 1532 2313
rect 1470 2245 1532 2279
rect -4734 2183 -4718 2217
rect -4684 2183 -4672 2217
rect 1470 2211 1482 2245
rect 1516 2211 1532 2245
rect -4734 2149 -4672 2183
rect -4734 2115 -4718 2149
rect -4684 2115 -4672 2149
rect -4734 2081 -4672 2115
rect -4734 2047 -4718 2081
rect -4684 2047 -4672 2081
rect -4734 2013 -4672 2047
rect -4734 1979 -4718 2013
rect -4684 1979 -4672 2013
rect -4734 1945 -4672 1979
rect -4734 1911 -4718 1945
rect -4684 1911 -4672 1945
rect -4734 1870 -4672 1911
rect 1470 2177 1532 2211
rect 1470 2143 1482 2177
rect 1516 2143 1532 2177
rect 1470 2109 1532 2143
rect 1470 2075 1482 2109
rect 1516 2075 1532 2109
rect 1470 2041 1532 2075
rect 1470 2007 1482 2041
rect 1516 2007 1532 2041
rect 1470 1973 1532 2007
rect 1470 1939 1482 1973
rect 1516 1939 1532 1973
rect 1470 1905 1532 1939
rect 1470 1871 1482 1905
rect 1516 1871 1532 1905
rect 1470 1830 1532 1871
rect 1562 2789 1628 2830
rect 1562 2755 1578 2789
rect 1612 2755 1628 2789
rect 1562 2721 1628 2755
rect 1562 2687 1578 2721
rect 1612 2687 1628 2721
rect 1562 2653 1628 2687
rect 1562 2619 1578 2653
rect 1612 2619 1628 2653
rect 1562 2585 1628 2619
rect 1562 2551 1578 2585
rect 1612 2551 1628 2585
rect 1562 2517 1628 2551
rect 1562 2483 1578 2517
rect 1612 2483 1628 2517
rect 1562 2449 1628 2483
rect 1562 2415 1578 2449
rect 1612 2415 1628 2449
rect 1562 2381 1628 2415
rect 1562 2347 1578 2381
rect 1612 2347 1628 2381
rect 1562 2313 1628 2347
rect 1562 2279 1578 2313
rect 1612 2279 1628 2313
rect 1562 2245 1628 2279
rect 1562 2211 1578 2245
rect 1612 2211 1628 2245
rect 1562 2177 1628 2211
rect 1562 2143 1578 2177
rect 1612 2143 1628 2177
rect 1562 2109 1628 2143
rect 1562 2075 1578 2109
rect 1612 2075 1628 2109
rect 1562 2041 1628 2075
rect 1562 2007 1578 2041
rect 1612 2007 1628 2041
rect 1562 1973 1628 2007
rect 1562 1939 1578 1973
rect 1612 1939 1628 1973
rect 1562 1905 1628 1939
rect 1562 1871 1578 1905
rect 1612 1871 1628 1905
rect 1562 1830 1628 1871
rect 1658 2789 1724 2830
rect 1658 2755 1674 2789
rect 1708 2755 1724 2789
rect 1658 2721 1724 2755
rect 1658 2687 1674 2721
rect 1708 2687 1724 2721
rect 1658 2653 1724 2687
rect 1658 2619 1674 2653
rect 1708 2619 1724 2653
rect 1658 2585 1724 2619
rect 1658 2551 1674 2585
rect 1708 2551 1724 2585
rect 1658 2517 1724 2551
rect 1658 2483 1674 2517
rect 1708 2483 1724 2517
rect 1658 2449 1724 2483
rect 1658 2415 1674 2449
rect 1708 2415 1724 2449
rect 1658 2381 1724 2415
rect 1658 2347 1674 2381
rect 1708 2347 1724 2381
rect 1658 2313 1724 2347
rect 1658 2279 1674 2313
rect 1708 2279 1724 2313
rect 1658 2245 1724 2279
rect 1658 2211 1674 2245
rect 1708 2211 1724 2245
rect 1658 2177 1724 2211
rect 1658 2143 1674 2177
rect 1708 2143 1724 2177
rect 1658 2109 1724 2143
rect 1658 2075 1674 2109
rect 1708 2075 1724 2109
rect 1658 2041 1724 2075
rect 1658 2007 1674 2041
rect 1708 2007 1724 2041
rect 1658 1973 1724 2007
rect 1658 1939 1674 1973
rect 1708 1939 1724 1973
rect 1658 1905 1724 1939
rect 1658 1871 1674 1905
rect 1708 1871 1724 1905
rect 1658 1830 1724 1871
rect 1754 2789 1820 2830
rect 1754 2755 1770 2789
rect 1804 2755 1820 2789
rect 1754 2721 1820 2755
rect 1754 2687 1770 2721
rect 1804 2687 1820 2721
rect 1754 2653 1820 2687
rect 1754 2619 1770 2653
rect 1804 2619 1820 2653
rect 1754 2585 1820 2619
rect 1754 2551 1770 2585
rect 1804 2551 1820 2585
rect 1754 2517 1820 2551
rect 1754 2483 1770 2517
rect 1804 2483 1820 2517
rect 1754 2449 1820 2483
rect 1754 2415 1770 2449
rect 1804 2415 1820 2449
rect 1754 2381 1820 2415
rect 1754 2347 1770 2381
rect 1804 2347 1820 2381
rect 1754 2313 1820 2347
rect 1754 2279 1770 2313
rect 1804 2279 1820 2313
rect 1754 2245 1820 2279
rect 1754 2211 1770 2245
rect 1804 2211 1820 2245
rect 1754 2177 1820 2211
rect 1754 2143 1770 2177
rect 1804 2143 1820 2177
rect 1754 2109 1820 2143
rect 1754 2075 1770 2109
rect 1804 2075 1820 2109
rect 1754 2041 1820 2075
rect 1754 2007 1770 2041
rect 1804 2007 1820 2041
rect 1754 1973 1820 2007
rect 1754 1939 1770 1973
rect 1804 1939 1820 1973
rect 1754 1905 1820 1939
rect 1754 1871 1770 1905
rect 1804 1871 1820 1905
rect 1754 1830 1820 1871
rect 1850 2789 1912 2830
rect 16674 2949 16736 2983
rect 16674 2915 16686 2949
rect 16720 2915 16736 2949
rect 16674 2881 16736 2915
rect 1850 2755 1866 2789
rect 1900 2755 1912 2789
rect 1850 2721 1912 2755
rect 1850 2687 1866 2721
rect 1900 2687 1912 2721
rect 1850 2653 1912 2687
rect 1850 2619 1866 2653
rect 1900 2619 1912 2653
rect 1850 2585 1912 2619
rect 1850 2551 1866 2585
rect 1900 2551 1912 2585
rect 1850 2517 1912 2551
rect 1850 2483 1866 2517
rect 1900 2483 1912 2517
rect 1850 2449 1912 2483
rect 1850 2415 1866 2449
rect 1900 2415 1912 2449
rect 4426 2773 4488 2814
rect 4426 2739 4438 2773
rect 4472 2739 4488 2773
rect 4426 2705 4488 2739
rect 4426 2671 4438 2705
rect 4472 2671 4488 2705
rect 4426 2637 4488 2671
rect 4426 2603 4438 2637
rect 4472 2603 4488 2637
rect 4426 2569 4488 2603
rect 4426 2535 4438 2569
rect 4472 2535 4488 2569
rect 4426 2501 4488 2535
rect 4426 2467 4438 2501
rect 4472 2467 4488 2501
rect 1850 2381 1912 2415
rect 1850 2347 1866 2381
rect 1900 2347 1912 2381
rect 1850 2313 1912 2347
rect 1850 2279 1866 2313
rect 1900 2279 1912 2313
rect 1850 2245 1912 2279
rect 4426 2433 4488 2467
rect 4426 2399 4438 2433
rect 4472 2399 4488 2433
rect 4426 2365 4488 2399
rect 4426 2331 4438 2365
rect 4472 2331 4488 2365
rect 4426 2297 4488 2331
rect 1850 2211 1866 2245
rect 1900 2211 1912 2245
rect 1850 2177 1912 2211
rect 1850 2143 1866 2177
rect 1900 2143 1912 2177
rect 1850 2109 1912 2143
rect 1850 2075 1866 2109
rect 1900 2075 1912 2109
rect 2488 2261 2546 2276
rect 2488 2227 2500 2261
rect 2534 2227 2546 2261
rect 2488 2193 2546 2227
rect 2488 2159 2500 2193
rect 2534 2159 2546 2193
rect 2488 2125 2546 2159
rect 2488 2091 2500 2125
rect 2534 2091 2546 2125
rect 2488 2076 2546 2091
rect 2646 2261 2704 2276
rect 2646 2227 2658 2261
rect 2692 2227 2704 2261
rect 2646 2193 2704 2227
rect 2646 2159 2658 2193
rect 2692 2159 2704 2193
rect 2646 2125 2704 2159
rect 2646 2091 2658 2125
rect 2692 2091 2704 2125
rect 2646 2076 2704 2091
rect 4426 2263 4438 2297
rect 4472 2263 4488 2297
rect 4426 2229 4488 2263
rect 4426 2195 4438 2229
rect 4472 2195 4488 2229
rect 4426 2161 4488 2195
rect 4426 2127 4438 2161
rect 4472 2127 4488 2161
rect 4426 2093 4488 2127
rect 1850 2041 1912 2075
rect 4426 2059 4438 2093
rect 4472 2059 4488 2093
rect 1850 2007 1866 2041
rect 1900 2007 1912 2041
rect 1850 1973 1912 2007
rect 1850 1939 1866 1973
rect 1900 1939 1912 1973
rect 1850 1905 1912 1939
rect 1850 1871 1866 1905
rect 1900 1871 1912 1905
rect 1850 1830 1912 1871
rect 4426 2025 4488 2059
rect 4426 1991 4438 2025
rect 4472 1991 4488 2025
rect 4426 1957 4488 1991
rect 4426 1923 4438 1957
rect 4472 1923 4488 1957
rect 4426 1889 4488 1923
rect 4426 1855 4438 1889
rect 4472 1855 4488 1889
rect 4426 1814 4488 1855
rect 4518 2773 4584 2814
rect 4518 2739 4534 2773
rect 4568 2739 4584 2773
rect 4518 2705 4584 2739
rect 4518 2671 4534 2705
rect 4568 2671 4584 2705
rect 4518 2637 4584 2671
rect 4518 2603 4534 2637
rect 4568 2603 4584 2637
rect 4518 2569 4584 2603
rect 4518 2535 4534 2569
rect 4568 2535 4584 2569
rect 4518 2501 4584 2535
rect 4518 2467 4534 2501
rect 4568 2467 4584 2501
rect 4518 2433 4584 2467
rect 4518 2399 4534 2433
rect 4568 2399 4584 2433
rect 4518 2365 4584 2399
rect 4518 2331 4534 2365
rect 4568 2331 4584 2365
rect 4518 2297 4584 2331
rect 4518 2263 4534 2297
rect 4568 2263 4584 2297
rect 4518 2229 4584 2263
rect 4518 2195 4534 2229
rect 4568 2195 4584 2229
rect 4518 2161 4584 2195
rect 4518 2127 4534 2161
rect 4568 2127 4584 2161
rect 4518 2093 4584 2127
rect 4518 2059 4534 2093
rect 4568 2059 4584 2093
rect 4518 2025 4584 2059
rect 4518 1991 4534 2025
rect 4568 1991 4584 2025
rect 4518 1957 4584 1991
rect 4518 1923 4534 1957
rect 4568 1923 4584 1957
rect 4518 1889 4584 1923
rect 4518 1855 4534 1889
rect 4568 1855 4584 1889
rect 4518 1814 4584 1855
rect 4614 2773 4680 2814
rect 4614 2739 4630 2773
rect 4664 2739 4680 2773
rect 4614 2705 4680 2739
rect 4614 2671 4630 2705
rect 4664 2671 4680 2705
rect 4614 2637 4680 2671
rect 4614 2603 4630 2637
rect 4664 2603 4680 2637
rect 4614 2569 4680 2603
rect 4614 2535 4630 2569
rect 4664 2535 4680 2569
rect 4614 2501 4680 2535
rect 4614 2467 4630 2501
rect 4664 2467 4680 2501
rect 4614 2433 4680 2467
rect 4614 2399 4630 2433
rect 4664 2399 4680 2433
rect 4614 2365 4680 2399
rect 4614 2331 4630 2365
rect 4664 2331 4680 2365
rect 4614 2297 4680 2331
rect 4614 2263 4630 2297
rect 4664 2263 4680 2297
rect 4614 2229 4680 2263
rect 4614 2195 4630 2229
rect 4664 2195 4680 2229
rect 4614 2161 4680 2195
rect 4614 2127 4630 2161
rect 4664 2127 4680 2161
rect 4614 2093 4680 2127
rect 4614 2059 4630 2093
rect 4664 2059 4680 2093
rect 4614 2025 4680 2059
rect 4614 1991 4630 2025
rect 4664 1991 4680 2025
rect 4614 1957 4680 1991
rect 4614 1923 4630 1957
rect 4664 1923 4680 1957
rect 4614 1889 4680 1923
rect 4614 1855 4630 1889
rect 4664 1855 4680 1889
rect 4614 1814 4680 1855
rect 4710 2773 4776 2814
rect 4710 2739 4726 2773
rect 4760 2739 4776 2773
rect 4710 2705 4776 2739
rect 4710 2671 4726 2705
rect 4760 2671 4776 2705
rect 4710 2637 4776 2671
rect 4710 2603 4726 2637
rect 4760 2603 4776 2637
rect 4710 2569 4776 2603
rect 4710 2535 4726 2569
rect 4760 2535 4776 2569
rect 4710 2501 4776 2535
rect 4710 2467 4726 2501
rect 4760 2467 4776 2501
rect 4710 2433 4776 2467
rect 4710 2399 4726 2433
rect 4760 2399 4776 2433
rect 4710 2365 4776 2399
rect 4710 2331 4726 2365
rect 4760 2331 4776 2365
rect 4710 2297 4776 2331
rect 4710 2263 4726 2297
rect 4760 2263 4776 2297
rect 4710 2229 4776 2263
rect 4710 2195 4726 2229
rect 4760 2195 4776 2229
rect 4710 2161 4776 2195
rect 4710 2127 4726 2161
rect 4760 2127 4776 2161
rect 4710 2093 4776 2127
rect 4710 2059 4726 2093
rect 4760 2059 4776 2093
rect 4710 2025 4776 2059
rect 4710 1991 4726 2025
rect 4760 1991 4776 2025
rect 4710 1957 4776 1991
rect 4710 1923 4726 1957
rect 4760 1923 4776 1957
rect 4710 1889 4776 1923
rect 4710 1855 4726 1889
rect 4760 1855 4776 1889
rect 4710 1814 4776 1855
rect 4806 2773 4868 2814
rect 4806 2739 4822 2773
rect 4856 2739 4868 2773
rect 4806 2705 4868 2739
rect 4806 2671 4822 2705
rect 4856 2671 4868 2705
rect 4806 2637 4868 2671
rect 4806 2603 4822 2637
rect 4856 2603 4868 2637
rect 4806 2569 4868 2603
rect 4806 2535 4822 2569
rect 4856 2535 4868 2569
rect 4806 2501 4868 2535
rect 4806 2467 4822 2501
rect 4856 2467 4868 2501
rect 4806 2433 4868 2467
rect 7456 2773 7518 2814
rect 7456 2739 7468 2773
rect 7502 2739 7518 2773
rect 7456 2705 7518 2739
rect 7456 2671 7468 2705
rect 7502 2671 7518 2705
rect 7456 2637 7518 2671
rect 7456 2603 7468 2637
rect 7502 2603 7518 2637
rect 7456 2569 7518 2603
rect 7456 2535 7468 2569
rect 7502 2535 7518 2569
rect 7456 2501 7518 2535
rect 7456 2467 7468 2501
rect 7502 2467 7518 2501
rect 4806 2399 4822 2433
rect 4856 2399 4868 2433
rect 4806 2365 4868 2399
rect 4806 2331 4822 2365
rect 4856 2331 4868 2365
rect 4806 2297 4868 2331
rect 4806 2263 4822 2297
rect 4856 2263 4868 2297
rect 7456 2433 7518 2467
rect 7456 2399 7468 2433
rect 7502 2399 7518 2433
rect 7456 2365 7518 2399
rect 7456 2331 7468 2365
rect 7502 2331 7518 2365
rect 7456 2297 7518 2331
rect 4806 2229 4868 2263
rect 4806 2195 4822 2229
rect 4856 2195 4868 2229
rect 4806 2161 4868 2195
rect 4806 2127 4822 2161
rect 4856 2127 4868 2161
rect 4806 2093 4868 2127
rect 4806 2059 4822 2093
rect 4856 2059 4868 2093
rect 5488 2261 5546 2276
rect 5488 2227 5500 2261
rect 5534 2227 5546 2261
rect 5488 2193 5546 2227
rect 5488 2159 5500 2193
rect 5534 2159 5546 2193
rect 5488 2125 5546 2159
rect 5488 2091 5500 2125
rect 5534 2091 5546 2125
rect 5488 2076 5546 2091
rect 5646 2261 5704 2276
rect 5646 2227 5658 2261
rect 5692 2227 5704 2261
rect 5646 2193 5704 2227
rect 5646 2159 5658 2193
rect 5692 2159 5704 2193
rect 5646 2125 5704 2159
rect 5646 2091 5658 2125
rect 5692 2091 5704 2125
rect 5646 2076 5704 2091
rect 7456 2263 7468 2297
rect 7502 2263 7518 2297
rect 7456 2229 7518 2263
rect 7456 2195 7468 2229
rect 7502 2195 7518 2229
rect 7456 2161 7518 2195
rect 7456 2127 7468 2161
rect 7502 2127 7518 2161
rect 7456 2093 7518 2127
rect 4806 2025 4868 2059
rect 7456 2059 7468 2093
rect 7502 2059 7518 2093
rect 4806 1991 4822 2025
rect 4856 1991 4868 2025
rect 4806 1957 4868 1991
rect 4806 1923 4822 1957
rect 4856 1923 4868 1957
rect 4806 1889 4868 1923
rect 4806 1855 4822 1889
rect 4856 1855 4868 1889
rect 4806 1814 4868 1855
rect 7456 2025 7518 2059
rect 7456 1991 7468 2025
rect 7502 1991 7518 2025
rect 7456 1957 7518 1991
rect 7456 1923 7468 1957
rect 7502 1923 7518 1957
rect 7456 1889 7518 1923
rect 7456 1855 7468 1889
rect 7502 1855 7518 1889
rect 7456 1814 7518 1855
rect 7548 2773 7614 2814
rect 7548 2739 7564 2773
rect 7598 2739 7614 2773
rect 7548 2705 7614 2739
rect 7548 2671 7564 2705
rect 7598 2671 7614 2705
rect 7548 2637 7614 2671
rect 7548 2603 7564 2637
rect 7598 2603 7614 2637
rect 7548 2569 7614 2603
rect 7548 2535 7564 2569
rect 7598 2535 7614 2569
rect 7548 2501 7614 2535
rect 7548 2467 7564 2501
rect 7598 2467 7614 2501
rect 7548 2433 7614 2467
rect 7548 2399 7564 2433
rect 7598 2399 7614 2433
rect 7548 2365 7614 2399
rect 7548 2331 7564 2365
rect 7598 2331 7614 2365
rect 7548 2297 7614 2331
rect 7548 2263 7564 2297
rect 7598 2263 7614 2297
rect 7548 2229 7614 2263
rect 7548 2195 7564 2229
rect 7598 2195 7614 2229
rect 7548 2161 7614 2195
rect 7548 2127 7564 2161
rect 7598 2127 7614 2161
rect 7548 2093 7614 2127
rect 7548 2059 7564 2093
rect 7598 2059 7614 2093
rect 7548 2025 7614 2059
rect 7548 1991 7564 2025
rect 7598 1991 7614 2025
rect 7548 1957 7614 1991
rect 7548 1923 7564 1957
rect 7598 1923 7614 1957
rect 7548 1889 7614 1923
rect 7548 1855 7564 1889
rect 7598 1855 7614 1889
rect 7548 1814 7614 1855
rect 7644 2773 7710 2814
rect 7644 2739 7660 2773
rect 7694 2739 7710 2773
rect 7644 2705 7710 2739
rect 7644 2671 7660 2705
rect 7694 2671 7710 2705
rect 7644 2637 7710 2671
rect 7644 2603 7660 2637
rect 7694 2603 7710 2637
rect 7644 2569 7710 2603
rect 7644 2535 7660 2569
rect 7694 2535 7710 2569
rect 7644 2501 7710 2535
rect 7644 2467 7660 2501
rect 7694 2467 7710 2501
rect 7644 2433 7710 2467
rect 7644 2399 7660 2433
rect 7694 2399 7710 2433
rect 7644 2365 7710 2399
rect 7644 2331 7660 2365
rect 7694 2331 7710 2365
rect 7644 2297 7710 2331
rect 7644 2263 7660 2297
rect 7694 2263 7710 2297
rect 7644 2229 7710 2263
rect 7644 2195 7660 2229
rect 7694 2195 7710 2229
rect 7644 2161 7710 2195
rect 7644 2127 7660 2161
rect 7694 2127 7710 2161
rect 7644 2093 7710 2127
rect 7644 2059 7660 2093
rect 7694 2059 7710 2093
rect 7644 2025 7710 2059
rect 7644 1991 7660 2025
rect 7694 1991 7710 2025
rect 7644 1957 7710 1991
rect 7644 1923 7660 1957
rect 7694 1923 7710 1957
rect 7644 1889 7710 1923
rect 7644 1855 7660 1889
rect 7694 1855 7710 1889
rect 7644 1814 7710 1855
rect 7740 2773 7806 2814
rect 7740 2739 7756 2773
rect 7790 2739 7806 2773
rect 7740 2705 7806 2739
rect 7740 2671 7756 2705
rect 7790 2671 7806 2705
rect 7740 2637 7806 2671
rect 7740 2603 7756 2637
rect 7790 2603 7806 2637
rect 7740 2569 7806 2603
rect 7740 2535 7756 2569
rect 7790 2535 7806 2569
rect 7740 2501 7806 2535
rect 7740 2467 7756 2501
rect 7790 2467 7806 2501
rect 7740 2433 7806 2467
rect 7740 2399 7756 2433
rect 7790 2399 7806 2433
rect 7740 2365 7806 2399
rect 7740 2331 7756 2365
rect 7790 2331 7806 2365
rect 7740 2297 7806 2331
rect 7740 2263 7756 2297
rect 7790 2263 7806 2297
rect 7740 2229 7806 2263
rect 7740 2195 7756 2229
rect 7790 2195 7806 2229
rect 7740 2161 7806 2195
rect 7740 2127 7756 2161
rect 7790 2127 7806 2161
rect 7740 2093 7806 2127
rect 7740 2059 7756 2093
rect 7790 2059 7806 2093
rect 7740 2025 7806 2059
rect 7740 1991 7756 2025
rect 7790 1991 7806 2025
rect 7740 1957 7806 1991
rect 7740 1923 7756 1957
rect 7790 1923 7806 1957
rect 7740 1889 7806 1923
rect 7740 1855 7756 1889
rect 7790 1855 7806 1889
rect 7740 1814 7806 1855
rect 7836 2773 7898 2814
rect 7836 2739 7852 2773
rect 7886 2739 7898 2773
rect 7836 2705 7898 2739
rect 7836 2671 7852 2705
rect 7886 2671 7898 2705
rect 7836 2637 7898 2671
rect 7836 2603 7852 2637
rect 7886 2603 7898 2637
rect 7836 2569 7898 2603
rect 7836 2535 7852 2569
rect 7886 2535 7898 2569
rect 7836 2501 7898 2535
rect 7836 2467 7852 2501
rect 7886 2467 7898 2501
rect 7836 2433 7898 2467
rect 10544 2771 10606 2812
rect 10544 2737 10556 2771
rect 10590 2737 10606 2771
rect 10544 2703 10606 2737
rect 10544 2669 10556 2703
rect 10590 2669 10606 2703
rect 10544 2635 10606 2669
rect 10544 2601 10556 2635
rect 10590 2601 10606 2635
rect 10544 2567 10606 2601
rect 10544 2533 10556 2567
rect 10590 2533 10606 2567
rect 10544 2499 10606 2533
rect 10544 2465 10556 2499
rect 10590 2465 10606 2499
rect 7836 2399 7852 2433
rect 7886 2399 7898 2433
rect 7836 2365 7898 2399
rect 7836 2331 7852 2365
rect 7886 2331 7898 2365
rect 7836 2297 7898 2331
rect 7836 2263 7852 2297
rect 7886 2263 7898 2297
rect 10544 2431 10606 2465
rect 10544 2397 10556 2431
rect 10590 2397 10606 2431
rect 10544 2363 10606 2397
rect 10544 2329 10556 2363
rect 10590 2329 10606 2363
rect 10544 2295 10606 2329
rect 7836 2229 7898 2263
rect 7836 2195 7852 2229
rect 7886 2195 7898 2229
rect 7836 2161 7898 2195
rect 7836 2127 7852 2161
rect 7886 2127 7898 2161
rect 7836 2093 7898 2127
rect 7836 2059 7852 2093
rect 7886 2059 7898 2093
rect 8488 2261 8546 2276
rect 8488 2227 8500 2261
rect 8534 2227 8546 2261
rect 8488 2193 8546 2227
rect 8488 2159 8500 2193
rect 8534 2159 8546 2193
rect 8488 2125 8546 2159
rect 8488 2091 8500 2125
rect 8534 2091 8546 2125
rect 8488 2076 8546 2091
rect 8646 2261 8704 2276
rect 8646 2227 8658 2261
rect 8692 2227 8704 2261
rect 8646 2193 8704 2227
rect 8646 2159 8658 2193
rect 8692 2159 8704 2193
rect 8646 2125 8704 2159
rect 8646 2091 8658 2125
rect 8692 2091 8704 2125
rect 8646 2076 8704 2091
rect 10544 2261 10556 2295
rect 10590 2261 10606 2295
rect 10544 2227 10606 2261
rect 10544 2193 10556 2227
rect 10590 2193 10606 2227
rect 10544 2159 10606 2193
rect 10544 2125 10556 2159
rect 10590 2125 10606 2159
rect 10544 2091 10606 2125
rect 7836 2025 7898 2059
rect 10544 2057 10556 2091
rect 10590 2057 10606 2091
rect 7836 1991 7852 2025
rect 7886 1991 7898 2025
rect 7836 1957 7898 1991
rect 7836 1923 7852 1957
rect 7886 1923 7898 1957
rect 7836 1889 7898 1923
rect 7836 1855 7852 1889
rect 7886 1855 7898 1889
rect 7836 1814 7898 1855
rect 10544 2023 10606 2057
rect 10544 1989 10556 2023
rect 10590 1989 10606 2023
rect 10544 1955 10606 1989
rect 10544 1921 10556 1955
rect 10590 1921 10606 1955
rect 10544 1887 10606 1921
rect 10544 1853 10556 1887
rect 10590 1853 10606 1887
rect 10544 1812 10606 1853
rect 10636 2771 10702 2812
rect 10636 2737 10652 2771
rect 10686 2737 10702 2771
rect 10636 2703 10702 2737
rect 10636 2669 10652 2703
rect 10686 2669 10702 2703
rect 10636 2635 10702 2669
rect 10636 2601 10652 2635
rect 10686 2601 10702 2635
rect 10636 2567 10702 2601
rect 10636 2533 10652 2567
rect 10686 2533 10702 2567
rect 10636 2499 10702 2533
rect 10636 2465 10652 2499
rect 10686 2465 10702 2499
rect 10636 2431 10702 2465
rect 10636 2397 10652 2431
rect 10686 2397 10702 2431
rect 10636 2363 10702 2397
rect 10636 2329 10652 2363
rect 10686 2329 10702 2363
rect 10636 2295 10702 2329
rect 10636 2261 10652 2295
rect 10686 2261 10702 2295
rect 10636 2227 10702 2261
rect 10636 2193 10652 2227
rect 10686 2193 10702 2227
rect 10636 2159 10702 2193
rect 10636 2125 10652 2159
rect 10686 2125 10702 2159
rect 10636 2091 10702 2125
rect 10636 2057 10652 2091
rect 10686 2057 10702 2091
rect 10636 2023 10702 2057
rect 10636 1989 10652 2023
rect 10686 1989 10702 2023
rect 10636 1955 10702 1989
rect 10636 1921 10652 1955
rect 10686 1921 10702 1955
rect 10636 1887 10702 1921
rect 10636 1853 10652 1887
rect 10686 1853 10702 1887
rect 10636 1812 10702 1853
rect 10732 2771 10798 2812
rect 10732 2737 10748 2771
rect 10782 2737 10798 2771
rect 10732 2703 10798 2737
rect 10732 2669 10748 2703
rect 10782 2669 10798 2703
rect 10732 2635 10798 2669
rect 10732 2601 10748 2635
rect 10782 2601 10798 2635
rect 10732 2567 10798 2601
rect 10732 2533 10748 2567
rect 10782 2533 10798 2567
rect 10732 2499 10798 2533
rect 10732 2465 10748 2499
rect 10782 2465 10798 2499
rect 10732 2431 10798 2465
rect 10732 2397 10748 2431
rect 10782 2397 10798 2431
rect 10732 2363 10798 2397
rect 10732 2329 10748 2363
rect 10782 2329 10798 2363
rect 10732 2295 10798 2329
rect 10732 2261 10748 2295
rect 10782 2261 10798 2295
rect 10732 2227 10798 2261
rect 10732 2193 10748 2227
rect 10782 2193 10798 2227
rect 10732 2159 10798 2193
rect 10732 2125 10748 2159
rect 10782 2125 10798 2159
rect 10732 2091 10798 2125
rect 10732 2057 10748 2091
rect 10782 2057 10798 2091
rect 10732 2023 10798 2057
rect 10732 1989 10748 2023
rect 10782 1989 10798 2023
rect 10732 1955 10798 1989
rect 10732 1921 10748 1955
rect 10782 1921 10798 1955
rect 10732 1887 10798 1921
rect 10732 1853 10748 1887
rect 10782 1853 10798 1887
rect 10732 1812 10798 1853
rect 10828 2771 10894 2812
rect 10828 2737 10844 2771
rect 10878 2737 10894 2771
rect 10828 2703 10894 2737
rect 10828 2669 10844 2703
rect 10878 2669 10894 2703
rect 10828 2635 10894 2669
rect 10828 2601 10844 2635
rect 10878 2601 10894 2635
rect 10828 2567 10894 2601
rect 10828 2533 10844 2567
rect 10878 2533 10894 2567
rect 10828 2499 10894 2533
rect 10828 2465 10844 2499
rect 10878 2465 10894 2499
rect 10828 2431 10894 2465
rect 10828 2397 10844 2431
rect 10878 2397 10894 2431
rect 10828 2363 10894 2397
rect 10828 2329 10844 2363
rect 10878 2329 10894 2363
rect 10828 2295 10894 2329
rect 10828 2261 10844 2295
rect 10878 2261 10894 2295
rect 10828 2227 10894 2261
rect 10828 2193 10844 2227
rect 10878 2193 10894 2227
rect 10828 2159 10894 2193
rect 10828 2125 10844 2159
rect 10878 2125 10894 2159
rect 10828 2091 10894 2125
rect 10828 2057 10844 2091
rect 10878 2057 10894 2091
rect 10828 2023 10894 2057
rect 10828 1989 10844 2023
rect 10878 1989 10894 2023
rect 10828 1955 10894 1989
rect 10828 1921 10844 1955
rect 10878 1921 10894 1955
rect 10828 1887 10894 1921
rect 10828 1853 10844 1887
rect 10878 1853 10894 1887
rect 10828 1812 10894 1853
rect 10924 2771 10986 2812
rect 16674 2847 16686 2881
rect 16720 2847 16736 2881
rect 16674 2813 16736 2847
rect 10924 2737 10940 2771
rect 10974 2737 10986 2771
rect 10924 2703 10986 2737
rect 10924 2669 10940 2703
rect 10974 2669 10986 2703
rect 10924 2635 10986 2669
rect 10924 2601 10940 2635
rect 10974 2601 10986 2635
rect 10924 2567 10986 2601
rect 10924 2533 10940 2567
rect 10974 2533 10986 2567
rect 10924 2499 10986 2533
rect 10924 2465 10940 2499
rect 10974 2465 10986 2499
rect 10924 2431 10986 2465
rect 13700 2745 13762 2786
rect 13700 2711 13712 2745
rect 13746 2711 13762 2745
rect 13700 2677 13762 2711
rect 13700 2643 13712 2677
rect 13746 2643 13762 2677
rect 13700 2609 13762 2643
rect 13700 2575 13712 2609
rect 13746 2575 13762 2609
rect 13700 2541 13762 2575
rect 13700 2507 13712 2541
rect 13746 2507 13762 2541
rect 13700 2473 13762 2507
rect 10924 2397 10940 2431
rect 10974 2397 10986 2431
rect 10924 2363 10986 2397
rect 10924 2329 10940 2363
rect 10974 2329 10986 2363
rect 10924 2295 10986 2329
rect 10924 2261 10940 2295
rect 10974 2261 10986 2295
rect 13700 2439 13712 2473
rect 13746 2439 13762 2473
rect 13700 2405 13762 2439
rect 13700 2371 13712 2405
rect 13746 2371 13762 2405
rect 13700 2337 13762 2371
rect 13700 2303 13712 2337
rect 13746 2303 13762 2337
rect 10924 2227 10986 2261
rect 10924 2193 10940 2227
rect 10974 2193 10986 2227
rect 10924 2159 10986 2193
rect 10924 2125 10940 2159
rect 10974 2125 10986 2159
rect 10924 2091 10986 2125
rect 10924 2057 10940 2091
rect 10974 2057 10986 2091
rect 11488 2261 11546 2276
rect 11488 2227 11500 2261
rect 11534 2227 11546 2261
rect 11488 2193 11546 2227
rect 11488 2159 11500 2193
rect 11534 2159 11546 2193
rect 11488 2125 11546 2159
rect 11488 2091 11500 2125
rect 11534 2091 11546 2125
rect 11488 2076 11546 2091
rect 11646 2261 11704 2276
rect 11646 2227 11658 2261
rect 11692 2227 11704 2261
rect 11646 2193 11704 2227
rect 11646 2159 11658 2193
rect 11692 2159 11704 2193
rect 11646 2125 11704 2159
rect 11646 2091 11658 2125
rect 11692 2091 11704 2125
rect 11646 2076 11704 2091
rect 13700 2269 13762 2303
rect 13700 2235 13712 2269
rect 13746 2235 13762 2269
rect 13700 2201 13762 2235
rect 13700 2167 13712 2201
rect 13746 2167 13762 2201
rect 13700 2133 13762 2167
rect 13700 2099 13712 2133
rect 13746 2099 13762 2133
rect 10924 2023 10986 2057
rect 13700 2065 13762 2099
rect 10924 1989 10940 2023
rect 10974 1989 10986 2023
rect 10924 1955 10986 1989
rect 10924 1921 10940 1955
rect 10974 1921 10986 1955
rect 10924 1887 10986 1921
rect 10924 1853 10940 1887
rect 10974 1853 10986 1887
rect 10924 1812 10986 1853
rect 13700 2031 13712 2065
rect 13746 2031 13762 2065
rect 13700 1997 13762 2031
rect 13700 1963 13712 1997
rect 13746 1963 13762 1997
rect 13700 1929 13762 1963
rect 13700 1895 13712 1929
rect 13746 1895 13762 1929
rect 13700 1861 13762 1895
rect 13700 1827 13712 1861
rect 13746 1827 13762 1861
rect 13700 1786 13762 1827
rect 13792 2745 13858 2786
rect 13792 2711 13808 2745
rect 13842 2711 13858 2745
rect 13792 2677 13858 2711
rect 13792 2643 13808 2677
rect 13842 2643 13858 2677
rect 13792 2609 13858 2643
rect 13792 2575 13808 2609
rect 13842 2575 13858 2609
rect 13792 2541 13858 2575
rect 13792 2507 13808 2541
rect 13842 2507 13858 2541
rect 13792 2473 13858 2507
rect 13792 2439 13808 2473
rect 13842 2439 13858 2473
rect 13792 2405 13858 2439
rect 13792 2371 13808 2405
rect 13842 2371 13858 2405
rect 13792 2337 13858 2371
rect 13792 2303 13808 2337
rect 13842 2303 13858 2337
rect 13792 2269 13858 2303
rect 13792 2235 13808 2269
rect 13842 2235 13858 2269
rect 13792 2201 13858 2235
rect 13792 2167 13808 2201
rect 13842 2167 13858 2201
rect 13792 2133 13858 2167
rect 13792 2099 13808 2133
rect 13842 2099 13858 2133
rect 13792 2065 13858 2099
rect 13792 2031 13808 2065
rect 13842 2031 13858 2065
rect 13792 1997 13858 2031
rect 13792 1963 13808 1997
rect 13842 1963 13858 1997
rect 13792 1929 13858 1963
rect 13792 1895 13808 1929
rect 13842 1895 13858 1929
rect 13792 1861 13858 1895
rect 13792 1827 13808 1861
rect 13842 1827 13858 1861
rect 13792 1786 13858 1827
rect 13888 2745 13954 2786
rect 13888 2711 13904 2745
rect 13938 2711 13954 2745
rect 13888 2677 13954 2711
rect 13888 2643 13904 2677
rect 13938 2643 13954 2677
rect 13888 2609 13954 2643
rect 13888 2575 13904 2609
rect 13938 2575 13954 2609
rect 13888 2541 13954 2575
rect 13888 2507 13904 2541
rect 13938 2507 13954 2541
rect 13888 2473 13954 2507
rect 13888 2439 13904 2473
rect 13938 2439 13954 2473
rect 13888 2405 13954 2439
rect 13888 2371 13904 2405
rect 13938 2371 13954 2405
rect 13888 2337 13954 2371
rect 13888 2303 13904 2337
rect 13938 2303 13954 2337
rect 13888 2269 13954 2303
rect 13888 2235 13904 2269
rect 13938 2235 13954 2269
rect 13888 2201 13954 2235
rect 13888 2167 13904 2201
rect 13938 2167 13954 2201
rect 13888 2133 13954 2167
rect 13888 2099 13904 2133
rect 13938 2099 13954 2133
rect 13888 2065 13954 2099
rect 13888 2031 13904 2065
rect 13938 2031 13954 2065
rect 13888 1997 13954 2031
rect 13888 1963 13904 1997
rect 13938 1963 13954 1997
rect 13888 1929 13954 1963
rect 13888 1895 13904 1929
rect 13938 1895 13954 1929
rect 13888 1861 13954 1895
rect 13888 1827 13904 1861
rect 13938 1827 13954 1861
rect 13888 1786 13954 1827
rect 13984 2745 14050 2786
rect 13984 2711 14000 2745
rect 14034 2711 14050 2745
rect 13984 2677 14050 2711
rect 13984 2643 14000 2677
rect 14034 2643 14050 2677
rect 13984 2609 14050 2643
rect 13984 2575 14000 2609
rect 14034 2575 14050 2609
rect 13984 2541 14050 2575
rect 13984 2507 14000 2541
rect 14034 2507 14050 2541
rect 13984 2473 14050 2507
rect 13984 2439 14000 2473
rect 14034 2439 14050 2473
rect 13984 2405 14050 2439
rect 13984 2371 14000 2405
rect 14034 2371 14050 2405
rect 13984 2337 14050 2371
rect 13984 2303 14000 2337
rect 14034 2303 14050 2337
rect 13984 2269 14050 2303
rect 13984 2235 14000 2269
rect 14034 2235 14050 2269
rect 13984 2201 14050 2235
rect 13984 2167 14000 2201
rect 14034 2167 14050 2201
rect 13984 2133 14050 2167
rect 13984 2099 14000 2133
rect 14034 2099 14050 2133
rect 13984 2065 14050 2099
rect 13984 2031 14000 2065
rect 14034 2031 14050 2065
rect 13984 1997 14050 2031
rect 13984 1963 14000 1997
rect 14034 1963 14050 1997
rect 13984 1929 14050 1963
rect 13984 1895 14000 1929
rect 14034 1895 14050 1929
rect 13984 1861 14050 1895
rect 13984 1827 14000 1861
rect 14034 1827 14050 1861
rect 13984 1786 14050 1827
rect 14080 2745 14142 2786
rect 14080 2711 14096 2745
rect 14130 2711 14142 2745
rect 14080 2677 14142 2711
rect 14080 2643 14096 2677
rect 14130 2643 14142 2677
rect 14080 2609 14142 2643
rect 14080 2575 14096 2609
rect 14130 2575 14142 2609
rect 14080 2541 14142 2575
rect 14080 2507 14096 2541
rect 14130 2507 14142 2541
rect 16674 2779 16686 2813
rect 16720 2779 16736 2813
rect 16674 2745 16736 2779
rect 16674 2711 16686 2745
rect 16720 2711 16736 2745
rect 16674 2677 16736 2711
rect 16674 2643 16686 2677
rect 16720 2643 16736 2677
rect 16674 2609 16736 2643
rect 16674 2575 16686 2609
rect 16720 2575 16736 2609
rect 16674 2534 16736 2575
rect 16766 3493 16832 3534
rect 16766 3459 16782 3493
rect 16816 3459 16832 3493
rect 16766 3425 16832 3459
rect 16766 3391 16782 3425
rect 16816 3391 16832 3425
rect 16766 3357 16832 3391
rect 16766 3323 16782 3357
rect 16816 3323 16832 3357
rect 16766 3289 16832 3323
rect 16766 3255 16782 3289
rect 16816 3255 16832 3289
rect 16766 3221 16832 3255
rect 16766 3187 16782 3221
rect 16816 3187 16832 3221
rect 16766 3153 16832 3187
rect 16766 3119 16782 3153
rect 16816 3119 16832 3153
rect 16766 3085 16832 3119
rect 16766 3051 16782 3085
rect 16816 3051 16832 3085
rect 16766 3017 16832 3051
rect 16766 2983 16782 3017
rect 16816 2983 16832 3017
rect 16766 2949 16832 2983
rect 16766 2915 16782 2949
rect 16816 2915 16832 2949
rect 16766 2881 16832 2915
rect 16766 2847 16782 2881
rect 16816 2847 16832 2881
rect 16766 2813 16832 2847
rect 16766 2779 16782 2813
rect 16816 2779 16832 2813
rect 16766 2745 16832 2779
rect 16766 2711 16782 2745
rect 16816 2711 16832 2745
rect 16766 2677 16832 2711
rect 16766 2643 16782 2677
rect 16816 2643 16832 2677
rect 16766 2609 16832 2643
rect 16766 2575 16782 2609
rect 16816 2575 16832 2609
rect 16766 2534 16832 2575
rect 16862 3493 16928 3534
rect 16862 3459 16878 3493
rect 16912 3459 16928 3493
rect 16862 3425 16928 3459
rect 16862 3391 16878 3425
rect 16912 3391 16928 3425
rect 16862 3357 16928 3391
rect 16862 3323 16878 3357
rect 16912 3323 16928 3357
rect 16862 3289 16928 3323
rect 16862 3255 16878 3289
rect 16912 3255 16928 3289
rect 16862 3221 16928 3255
rect 16862 3187 16878 3221
rect 16912 3187 16928 3221
rect 16862 3153 16928 3187
rect 16862 3119 16878 3153
rect 16912 3119 16928 3153
rect 16862 3085 16928 3119
rect 16862 3051 16878 3085
rect 16912 3051 16928 3085
rect 16862 3017 16928 3051
rect 16862 2983 16878 3017
rect 16912 2983 16928 3017
rect 16862 2949 16928 2983
rect 16862 2915 16878 2949
rect 16912 2915 16928 2949
rect 16862 2881 16928 2915
rect 16862 2847 16878 2881
rect 16912 2847 16928 2881
rect 16862 2813 16928 2847
rect 16862 2779 16878 2813
rect 16912 2779 16928 2813
rect 16862 2745 16928 2779
rect 16862 2711 16878 2745
rect 16912 2711 16928 2745
rect 16862 2677 16928 2711
rect 16862 2643 16878 2677
rect 16912 2643 16928 2677
rect 16862 2609 16928 2643
rect 16862 2575 16878 2609
rect 16912 2575 16928 2609
rect 16862 2534 16928 2575
rect 16958 3493 17024 3534
rect 16958 3459 16974 3493
rect 17008 3459 17024 3493
rect 16958 3425 17024 3459
rect 16958 3391 16974 3425
rect 17008 3391 17024 3425
rect 16958 3357 17024 3391
rect 16958 3323 16974 3357
rect 17008 3323 17024 3357
rect 16958 3289 17024 3323
rect 16958 3255 16974 3289
rect 17008 3255 17024 3289
rect 16958 3221 17024 3255
rect 16958 3187 16974 3221
rect 17008 3187 17024 3221
rect 16958 3153 17024 3187
rect 16958 3119 16974 3153
rect 17008 3119 17024 3153
rect 16958 3085 17024 3119
rect 16958 3051 16974 3085
rect 17008 3051 17024 3085
rect 16958 3017 17024 3051
rect 16958 2983 16974 3017
rect 17008 2983 17024 3017
rect 16958 2949 17024 2983
rect 16958 2915 16974 2949
rect 17008 2915 17024 2949
rect 16958 2881 17024 2915
rect 16958 2847 16974 2881
rect 17008 2847 17024 2881
rect 16958 2813 17024 2847
rect 16958 2779 16974 2813
rect 17008 2779 17024 2813
rect 16958 2745 17024 2779
rect 16958 2711 16974 2745
rect 17008 2711 17024 2745
rect 16958 2677 17024 2711
rect 16958 2643 16974 2677
rect 17008 2643 17024 2677
rect 16958 2609 17024 2643
rect 16958 2575 16974 2609
rect 17008 2575 17024 2609
rect 16958 2534 17024 2575
rect 17054 3493 17120 3534
rect 17054 3459 17070 3493
rect 17104 3459 17120 3493
rect 17054 3425 17120 3459
rect 17054 3391 17070 3425
rect 17104 3391 17120 3425
rect 17054 3357 17120 3391
rect 17054 3323 17070 3357
rect 17104 3323 17120 3357
rect 17054 3289 17120 3323
rect 17054 3255 17070 3289
rect 17104 3255 17120 3289
rect 17054 3221 17120 3255
rect 17054 3187 17070 3221
rect 17104 3187 17120 3221
rect 17054 3153 17120 3187
rect 17054 3119 17070 3153
rect 17104 3119 17120 3153
rect 17054 3085 17120 3119
rect 17054 3051 17070 3085
rect 17104 3051 17120 3085
rect 17054 3017 17120 3051
rect 17054 2983 17070 3017
rect 17104 2983 17120 3017
rect 17054 2949 17120 2983
rect 17054 2915 17070 2949
rect 17104 2915 17120 2949
rect 17054 2881 17120 2915
rect 17054 2847 17070 2881
rect 17104 2847 17120 2881
rect 17054 2813 17120 2847
rect 17054 2779 17070 2813
rect 17104 2779 17120 2813
rect 17054 2745 17120 2779
rect 17054 2711 17070 2745
rect 17104 2711 17120 2745
rect 17054 2677 17120 2711
rect 17054 2643 17070 2677
rect 17104 2643 17120 2677
rect 17054 2609 17120 2643
rect 17054 2575 17070 2609
rect 17104 2575 17120 2609
rect 17054 2534 17120 2575
rect 17150 3493 17212 3534
rect 17150 3459 17166 3493
rect 17200 3459 17212 3493
rect 17150 3425 17212 3459
rect 17150 3391 17166 3425
rect 17200 3391 17212 3425
rect 17150 3357 17212 3391
rect 17150 3323 17166 3357
rect 17200 3323 17212 3357
rect 17150 3289 17212 3323
rect 17150 3255 17166 3289
rect 17200 3255 17212 3289
rect 17150 3221 17212 3255
rect 17150 3187 17166 3221
rect 17200 3187 17212 3221
rect 17150 3153 17212 3187
rect 17150 3119 17166 3153
rect 17200 3119 17212 3153
rect 17150 3085 17212 3119
rect 17150 3051 17166 3085
rect 17200 3051 17212 3085
rect 17150 3017 17212 3051
rect 17150 2983 17166 3017
rect 17200 2983 17212 3017
rect 17150 2949 17212 2983
rect 17150 2915 17166 2949
rect 17200 2915 17212 2949
rect 17150 2881 17212 2915
rect 17150 2847 17166 2881
rect 17200 2847 17212 2881
rect 17150 2813 17212 2847
rect 17150 2779 17166 2813
rect 17200 2779 17212 2813
rect 17150 2745 17212 2779
rect 17150 2711 17166 2745
rect 17200 2711 17212 2745
rect 17150 2677 17212 2711
rect 17150 2643 17166 2677
rect 17200 2643 17212 2677
rect 17150 2609 17212 2643
rect 17150 2575 17166 2609
rect 17200 2575 17212 2609
rect 17150 2534 17212 2575
rect 17366 3483 17428 3524
rect 17366 3449 17378 3483
rect 17412 3449 17428 3483
rect 17366 3415 17428 3449
rect 17366 3381 17378 3415
rect 17412 3381 17428 3415
rect 17366 3347 17428 3381
rect 17366 3313 17378 3347
rect 17412 3313 17428 3347
rect 17366 3279 17428 3313
rect 17366 3245 17378 3279
rect 17412 3245 17428 3279
rect 17366 3211 17428 3245
rect 17366 3177 17378 3211
rect 17412 3177 17428 3211
rect 17366 3143 17428 3177
rect 17366 3109 17378 3143
rect 17412 3109 17428 3143
rect 17366 3075 17428 3109
rect 17366 3041 17378 3075
rect 17412 3041 17428 3075
rect 17366 3007 17428 3041
rect 17366 2973 17378 3007
rect 17412 2973 17428 3007
rect 17366 2939 17428 2973
rect 17366 2905 17378 2939
rect 17412 2905 17428 2939
rect 17366 2871 17428 2905
rect 17366 2837 17378 2871
rect 17412 2837 17428 2871
rect 17366 2803 17428 2837
rect 17366 2769 17378 2803
rect 17412 2769 17428 2803
rect 17366 2735 17428 2769
rect 17366 2701 17378 2735
rect 17412 2701 17428 2735
rect 17366 2667 17428 2701
rect 17366 2633 17378 2667
rect 17412 2633 17428 2667
rect 17366 2599 17428 2633
rect 17366 2565 17378 2599
rect 17412 2565 17428 2599
rect 17366 2524 17428 2565
rect 17458 3483 17524 3524
rect 17458 3449 17474 3483
rect 17508 3449 17524 3483
rect 17458 3415 17524 3449
rect 17458 3381 17474 3415
rect 17508 3381 17524 3415
rect 17458 3347 17524 3381
rect 17458 3313 17474 3347
rect 17508 3313 17524 3347
rect 17458 3279 17524 3313
rect 17458 3245 17474 3279
rect 17508 3245 17524 3279
rect 17458 3211 17524 3245
rect 17458 3177 17474 3211
rect 17508 3177 17524 3211
rect 17458 3143 17524 3177
rect 17458 3109 17474 3143
rect 17508 3109 17524 3143
rect 17458 3075 17524 3109
rect 17458 3041 17474 3075
rect 17508 3041 17524 3075
rect 17458 3007 17524 3041
rect 17458 2973 17474 3007
rect 17508 2973 17524 3007
rect 17458 2939 17524 2973
rect 17458 2905 17474 2939
rect 17508 2905 17524 2939
rect 17458 2871 17524 2905
rect 17458 2837 17474 2871
rect 17508 2837 17524 2871
rect 17458 2803 17524 2837
rect 17458 2769 17474 2803
rect 17508 2769 17524 2803
rect 17458 2735 17524 2769
rect 17458 2701 17474 2735
rect 17508 2701 17524 2735
rect 17458 2667 17524 2701
rect 17458 2633 17474 2667
rect 17508 2633 17524 2667
rect 17458 2599 17524 2633
rect 17458 2565 17474 2599
rect 17508 2565 17524 2599
rect 17458 2524 17524 2565
rect 17554 3483 17620 3524
rect 17554 3449 17570 3483
rect 17604 3449 17620 3483
rect 17554 3415 17620 3449
rect 17554 3381 17570 3415
rect 17604 3381 17620 3415
rect 17554 3347 17620 3381
rect 17554 3313 17570 3347
rect 17604 3313 17620 3347
rect 17554 3279 17620 3313
rect 17554 3245 17570 3279
rect 17604 3245 17620 3279
rect 17554 3211 17620 3245
rect 17554 3177 17570 3211
rect 17604 3177 17620 3211
rect 17554 3143 17620 3177
rect 17554 3109 17570 3143
rect 17604 3109 17620 3143
rect 17554 3075 17620 3109
rect 17554 3041 17570 3075
rect 17604 3041 17620 3075
rect 17554 3007 17620 3041
rect 17554 2973 17570 3007
rect 17604 2973 17620 3007
rect 17554 2939 17620 2973
rect 17554 2905 17570 2939
rect 17604 2905 17620 2939
rect 17554 2871 17620 2905
rect 17554 2837 17570 2871
rect 17604 2837 17620 2871
rect 17554 2803 17620 2837
rect 17554 2769 17570 2803
rect 17604 2769 17620 2803
rect 17554 2735 17620 2769
rect 17554 2701 17570 2735
rect 17604 2701 17620 2735
rect 17554 2667 17620 2701
rect 17554 2633 17570 2667
rect 17604 2633 17620 2667
rect 17554 2599 17620 2633
rect 17554 2565 17570 2599
rect 17604 2565 17620 2599
rect 17554 2524 17620 2565
rect 17650 3483 17716 3524
rect 17650 3449 17666 3483
rect 17700 3449 17716 3483
rect 17650 3415 17716 3449
rect 17650 3381 17666 3415
rect 17700 3381 17716 3415
rect 17650 3347 17716 3381
rect 17650 3313 17666 3347
rect 17700 3313 17716 3347
rect 17650 3279 17716 3313
rect 17650 3245 17666 3279
rect 17700 3245 17716 3279
rect 17650 3211 17716 3245
rect 17650 3177 17666 3211
rect 17700 3177 17716 3211
rect 17650 3143 17716 3177
rect 17650 3109 17666 3143
rect 17700 3109 17716 3143
rect 17650 3075 17716 3109
rect 17650 3041 17666 3075
rect 17700 3041 17716 3075
rect 17650 3007 17716 3041
rect 17650 2973 17666 3007
rect 17700 2973 17716 3007
rect 17650 2939 17716 2973
rect 17650 2905 17666 2939
rect 17700 2905 17716 2939
rect 17650 2871 17716 2905
rect 17650 2837 17666 2871
rect 17700 2837 17716 2871
rect 17650 2803 17716 2837
rect 17650 2769 17666 2803
rect 17700 2769 17716 2803
rect 17650 2735 17716 2769
rect 17650 2701 17666 2735
rect 17700 2701 17716 2735
rect 17650 2667 17716 2701
rect 17650 2633 17666 2667
rect 17700 2633 17716 2667
rect 17650 2599 17716 2633
rect 17650 2565 17666 2599
rect 17700 2565 17716 2599
rect 17650 2524 17716 2565
rect 17746 3483 17812 3524
rect 17746 3449 17762 3483
rect 17796 3449 17812 3483
rect 17746 3415 17812 3449
rect 17746 3381 17762 3415
rect 17796 3381 17812 3415
rect 17746 3347 17812 3381
rect 17746 3313 17762 3347
rect 17796 3313 17812 3347
rect 17746 3279 17812 3313
rect 17746 3245 17762 3279
rect 17796 3245 17812 3279
rect 17746 3211 17812 3245
rect 17746 3177 17762 3211
rect 17796 3177 17812 3211
rect 17746 3143 17812 3177
rect 17746 3109 17762 3143
rect 17796 3109 17812 3143
rect 17746 3075 17812 3109
rect 17746 3041 17762 3075
rect 17796 3041 17812 3075
rect 17746 3007 17812 3041
rect 17746 2973 17762 3007
rect 17796 2973 17812 3007
rect 17746 2939 17812 2973
rect 17746 2905 17762 2939
rect 17796 2905 17812 2939
rect 17746 2871 17812 2905
rect 17746 2837 17762 2871
rect 17796 2837 17812 2871
rect 17746 2803 17812 2837
rect 17746 2769 17762 2803
rect 17796 2769 17812 2803
rect 17746 2735 17812 2769
rect 17746 2701 17762 2735
rect 17796 2701 17812 2735
rect 17746 2667 17812 2701
rect 17746 2633 17762 2667
rect 17796 2633 17812 2667
rect 17746 2599 17812 2633
rect 17746 2565 17762 2599
rect 17796 2565 17812 2599
rect 17746 2524 17812 2565
rect 17842 3483 17908 3524
rect 17842 3449 17858 3483
rect 17892 3449 17908 3483
rect 17842 3415 17908 3449
rect 17842 3381 17858 3415
rect 17892 3381 17908 3415
rect 17842 3347 17908 3381
rect 17842 3313 17858 3347
rect 17892 3313 17908 3347
rect 17842 3279 17908 3313
rect 17842 3245 17858 3279
rect 17892 3245 17908 3279
rect 17842 3211 17908 3245
rect 17842 3177 17858 3211
rect 17892 3177 17908 3211
rect 17842 3143 17908 3177
rect 17842 3109 17858 3143
rect 17892 3109 17908 3143
rect 17842 3075 17908 3109
rect 17842 3041 17858 3075
rect 17892 3041 17908 3075
rect 17842 3007 17908 3041
rect 17842 2973 17858 3007
rect 17892 2973 17908 3007
rect 17842 2939 17908 2973
rect 17842 2905 17858 2939
rect 17892 2905 17908 2939
rect 17842 2871 17908 2905
rect 17842 2837 17858 2871
rect 17892 2837 17908 2871
rect 17842 2803 17908 2837
rect 17842 2769 17858 2803
rect 17892 2769 17908 2803
rect 17842 2735 17908 2769
rect 17842 2701 17858 2735
rect 17892 2701 17908 2735
rect 17842 2667 17908 2701
rect 17842 2633 17858 2667
rect 17892 2633 17908 2667
rect 17842 2599 17908 2633
rect 17842 2565 17858 2599
rect 17892 2565 17908 2599
rect 17842 2524 17908 2565
rect 17938 3483 18004 3524
rect 17938 3449 17954 3483
rect 17988 3449 18004 3483
rect 17938 3415 18004 3449
rect 17938 3381 17954 3415
rect 17988 3381 18004 3415
rect 17938 3347 18004 3381
rect 17938 3313 17954 3347
rect 17988 3313 18004 3347
rect 17938 3279 18004 3313
rect 17938 3245 17954 3279
rect 17988 3245 18004 3279
rect 17938 3211 18004 3245
rect 17938 3177 17954 3211
rect 17988 3177 18004 3211
rect 17938 3143 18004 3177
rect 17938 3109 17954 3143
rect 17988 3109 18004 3143
rect 17938 3075 18004 3109
rect 17938 3041 17954 3075
rect 17988 3041 18004 3075
rect 17938 3007 18004 3041
rect 17938 2973 17954 3007
rect 17988 2973 18004 3007
rect 17938 2939 18004 2973
rect 17938 2905 17954 2939
rect 17988 2905 18004 2939
rect 17938 2871 18004 2905
rect 17938 2837 17954 2871
rect 17988 2837 18004 2871
rect 17938 2803 18004 2837
rect 17938 2769 17954 2803
rect 17988 2769 18004 2803
rect 17938 2735 18004 2769
rect 17938 2701 17954 2735
rect 17988 2701 18004 2735
rect 17938 2667 18004 2701
rect 17938 2633 17954 2667
rect 17988 2633 18004 2667
rect 17938 2599 18004 2633
rect 17938 2565 17954 2599
rect 17988 2565 18004 2599
rect 17938 2524 18004 2565
rect 18034 3483 18100 3524
rect 18034 3449 18050 3483
rect 18084 3449 18100 3483
rect 18034 3415 18100 3449
rect 18034 3381 18050 3415
rect 18084 3381 18100 3415
rect 18034 3347 18100 3381
rect 18034 3313 18050 3347
rect 18084 3313 18100 3347
rect 18034 3279 18100 3313
rect 18034 3245 18050 3279
rect 18084 3245 18100 3279
rect 18034 3211 18100 3245
rect 18034 3177 18050 3211
rect 18084 3177 18100 3211
rect 18034 3143 18100 3177
rect 18034 3109 18050 3143
rect 18084 3109 18100 3143
rect 18034 3075 18100 3109
rect 18034 3041 18050 3075
rect 18084 3041 18100 3075
rect 18034 3007 18100 3041
rect 18034 2973 18050 3007
rect 18084 2973 18100 3007
rect 18034 2939 18100 2973
rect 18034 2905 18050 2939
rect 18084 2905 18100 2939
rect 18034 2871 18100 2905
rect 18034 2837 18050 2871
rect 18084 2837 18100 2871
rect 18034 2803 18100 2837
rect 18034 2769 18050 2803
rect 18084 2769 18100 2803
rect 18034 2735 18100 2769
rect 18034 2701 18050 2735
rect 18084 2701 18100 2735
rect 18034 2667 18100 2701
rect 18034 2633 18050 2667
rect 18084 2633 18100 2667
rect 18034 2599 18100 2633
rect 18034 2565 18050 2599
rect 18084 2565 18100 2599
rect 18034 2524 18100 2565
rect 18130 3483 18196 3524
rect 18130 3449 18146 3483
rect 18180 3449 18196 3483
rect 18130 3415 18196 3449
rect 18130 3381 18146 3415
rect 18180 3381 18196 3415
rect 18130 3347 18196 3381
rect 18130 3313 18146 3347
rect 18180 3313 18196 3347
rect 18130 3279 18196 3313
rect 18130 3245 18146 3279
rect 18180 3245 18196 3279
rect 18130 3211 18196 3245
rect 18130 3177 18146 3211
rect 18180 3177 18196 3211
rect 18130 3143 18196 3177
rect 18130 3109 18146 3143
rect 18180 3109 18196 3143
rect 18130 3075 18196 3109
rect 18130 3041 18146 3075
rect 18180 3041 18196 3075
rect 18130 3007 18196 3041
rect 18130 2973 18146 3007
rect 18180 2973 18196 3007
rect 18130 2939 18196 2973
rect 18130 2905 18146 2939
rect 18180 2905 18196 2939
rect 18130 2871 18196 2905
rect 18130 2837 18146 2871
rect 18180 2837 18196 2871
rect 18130 2803 18196 2837
rect 18130 2769 18146 2803
rect 18180 2769 18196 2803
rect 18130 2735 18196 2769
rect 18130 2701 18146 2735
rect 18180 2701 18196 2735
rect 18130 2667 18196 2701
rect 18130 2633 18146 2667
rect 18180 2633 18196 2667
rect 18130 2599 18196 2633
rect 18130 2565 18146 2599
rect 18180 2565 18196 2599
rect 18130 2524 18196 2565
rect 18226 3483 18292 3524
rect 18226 3449 18242 3483
rect 18276 3449 18292 3483
rect 18226 3415 18292 3449
rect 18226 3381 18242 3415
rect 18276 3381 18292 3415
rect 18226 3347 18292 3381
rect 18226 3313 18242 3347
rect 18276 3313 18292 3347
rect 18226 3279 18292 3313
rect 18226 3245 18242 3279
rect 18276 3245 18292 3279
rect 18226 3211 18292 3245
rect 18226 3177 18242 3211
rect 18276 3177 18292 3211
rect 18226 3143 18292 3177
rect 18226 3109 18242 3143
rect 18276 3109 18292 3143
rect 18226 3075 18292 3109
rect 18226 3041 18242 3075
rect 18276 3041 18292 3075
rect 18226 3007 18292 3041
rect 18226 2973 18242 3007
rect 18276 2973 18292 3007
rect 18226 2939 18292 2973
rect 18226 2905 18242 2939
rect 18276 2905 18292 2939
rect 18226 2871 18292 2905
rect 18226 2837 18242 2871
rect 18276 2837 18292 2871
rect 18226 2803 18292 2837
rect 18226 2769 18242 2803
rect 18276 2769 18292 2803
rect 18226 2735 18292 2769
rect 18226 2701 18242 2735
rect 18276 2701 18292 2735
rect 18226 2667 18292 2701
rect 18226 2633 18242 2667
rect 18276 2633 18292 2667
rect 18226 2599 18292 2633
rect 18226 2565 18242 2599
rect 18276 2565 18292 2599
rect 18226 2524 18292 2565
rect 18322 3483 18384 3524
rect 18322 3449 18338 3483
rect 18372 3449 18384 3483
rect 18322 3415 18384 3449
rect 18322 3381 18338 3415
rect 18372 3381 18384 3415
rect 18322 3347 18384 3381
rect 18322 3313 18338 3347
rect 18372 3313 18384 3347
rect 18322 3279 18384 3313
rect 18322 3245 18338 3279
rect 18372 3245 18384 3279
rect 18322 3211 18384 3245
rect 18322 3177 18338 3211
rect 18372 3177 18384 3211
rect 18322 3143 18384 3177
rect 18322 3109 18338 3143
rect 18372 3109 18384 3143
rect 18322 3075 18384 3109
rect 18322 3041 18338 3075
rect 18372 3041 18384 3075
rect 18322 3007 18384 3041
rect 18322 2973 18338 3007
rect 18372 2973 18384 3007
rect 18322 2939 18384 2973
rect 18322 2905 18338 2939
rect 18372 2905 18384 2939
rect 18322 2871 18384 2905
rect 18322 2837 18338 2871
rect 18372 2837 18384 2871
rect 18322 2803 18384 2837
rect 18322 2769 18338 2803
rect 18372 2769 18384 2803
rect 18322 2735 18384 2769
rect 18322 2701 18338 2735
rect 18372 2701 18384 2735
rect 18322 2667 18384 2701
rect 18322 2633 18338 2667
rect 18372 2633 18384 2667
rect 18322 2599 18384 2633
rect 18322 2565 18338 2599
rect 18372 2565 18384 2599
rect 18322 2524 18384 2565
rect 18564 3479 18626 3520
rect 18564 3445 18576 3479
rect 18610 3445 18626 3479
rect 18564 3411 18626 3445
rect 18564 3377 18576 3411
rect 18610 3377 18626 3411
rect 18564 3343 18626 3377
rect 18564 3309 18576 3343
rect 18610 3309 18626 3343
rect 18564 3275 18626 3309
rect 18564 3241 18576 3275
rect 18610 3241 18626 3275
rect 18564 3207 18626 3241
rect 18564 3173 18576 3207
rect 18610 3173 18626 3207
rect 18564 3139 18626 3173
rect 18564 3105 18576 3139
rect 18610 3105 18626 3139
rect 18564 3071 18626 3105
rect 18564 3037 18576 3071
rect 18610 3037 18626 3071
rect 18564 3003 18626 3037
rect 18564 2969 18576 3003
rect 18610 2969 18626 3003
rect 18564 2935 18626 2969
rect 18564 2901 18576 2935
rect 18610 2901 18626 2935
rect 18564 2867 18626 2901
rect 18564 2833 18576 2867
rect 18610 2833 18626 2867
rect 18564 2799 18626 2833
rect 18564 2765 18576 2799
rect 18610 2765 18626 2799
rect 18564 2731 18626 2765
rect 18564 2697 18576 2731
rect 18610 2697 18626 2731
rect 18564 2663 18626 2697
rect 18564 2629 18576 2663
rect 18610 2629 18626 2663
rect 18564 2595 18626 2629
rect 18564 2561 18576 2595
rect 18610 2561 18626 2595
rect 14080 2473 14142 2507
rect 18564 2520 18626 2561
rect 18656 3479 18722 3520
rect 18656 3445 18672 3479
rect 18706 3445 18722 3479
rect 18656 3411 18722 3445
rect 18656 3377 18672 3411
rect 18706 3377 18722 3411
rect 18656 3343 18722 3377
rect 18656 3309 18672 3343
rect 18706 3309 18722 3343
rect 18656 3275 18722 3309
rect 18656 3241 18672 3275
rect 18706 3241 18722 3275
rect 18656 3207 18722 3241
rect 18656 3173 18672 3207
rect 18706 3173 18722 3207
rect 18656 3139 18722 3173
rect 18656 3105 18672 3139
rect 18706 3105 18722 3139
rect 18656 3071 18722 3105
rect 18656 3037 18672 3071
rect 18706 3037 18722 3071
rect 18656 3003 18722 3037
rect 18656 2969 18672 3003
rect 18706 2969 18722 3003
rect 18656 2935 18722 2969
rect 18656 2901 18672 2935
rect 18706 2901 18722 2935
rect 18656 2867 18722 2901
rect 18656 2833 18672 2867
rect 18706 2833 18722 2867
rect 18656 2799 18722 2833
rect 18656 2765 18672 2799
rect 18706 2765 18722 2799
rect 18656 2731 18722 2765
rect 18656 2697 18672 2731
rect 18706 2697 18722 2731
rect 18656 2663 18722 2697
rect 18656 2629 18672 2663
rect 18706 2629 18722 2663
rect 18656 2595 18722 2629
rect 18656 2561 18672 2595
rect 18706 2561 18722 2595
rect 18656 2520 18722 2561
rect 18752 3479 18818 3520
rect 18752 3445 18768 3479
rect 18802 3445 18818 3479
rect 18752 3411 18818 3445
rect 18752 3377 18768 3411
rect 18802 3377 18818 3411
rect 18752 3343 18818 3377
rect 18752 3309 18768 3343
rect 18802 3309 18818 3343
rect 18752 3275 18818 3309
rect 18752 3241 18768 3275
rect 18802 3241 18818 3275
rect 18752 3207 18818 3241
rect 18752 3173 18768 3207
rect 18802 3173 18818 3207
rect 18752 3139 18818 3173
rect 18752 3105 18768 3139
rect 18802 3105 18818 3139
rect 18752 3071 18818 3105
rect 18752 3037 18768 3071
rect 18802 3037 18818 3071
rect 18752 3003 18818 3037
rect 18752 2969 18768 3003
rect 18802 2969 18818 3003
rect 18752 2935 18818 2969
rect 18752 2901 18768 2935
rect 18802 2901 18818 2935
rect 18752 2867 18818 2901
rect 18752 2833 18768 2867
rect 18802 2833 18818 2867
rect 18752 2799 18818 2833
rect 18752 2765 18768 2799
rect 18802 2765 18818 2799
rect 18752 2731 18818 2765
rect 18752 2697 18768 2731
rect 18802 2697 18818 2731
rect 18752 2663 18818 2697
rect 18752 2629 18768 2663
rect 18802 2629 18818 2663
rect 18752 2595 18818 2629
rect 18752 2561 18768 2595
rect 18802 2561 18818 2595
rect 18752 2520 18818 2561
rect 18848 3479 18914 3520
rect 18848 3445 18864 3479
rect 18898 3445 18914 3479
rect 18848 3411 18914 3445
rect 18848 3377 18864 3411
rect 18898 3377 18914 3411
rect 18848 3343 18914 3377
rect 18848 3309 18864 3343
rect 18898 3309 18914 3343
rect 18848 3275 18914 3309
rect 18848 3241 18864 3275
rect 18898 3241 18914 3275
rect 18848 3207 18914 3241
rect 18848 3173 18864 3207
rect 18898 3173 18914 3207
rect 18848 3139 18914 3173
rect 18848 3105 18864 3139
rect 18898 3105 18914 3139
rect 18848 3071 18914 3105
rect 18848 3037 18864 3071
rect 18898 3037 18914 3071
rect 18848 3003 18914 3037
rect 18848 2969 18864 3003
rect 18898 2969 18914 3003
rect 18848 2935 18914 2969
rect 18848 2901 18864 2935
rect 18898 2901 18914 2935
rect 18848 2867 18914 2901
rect 18848 2833 18864 2867
rect 18898 2833 18914 2867
rect 18848 2799 18914 2833
rect 18848 2765 18864 2799
rect 18898 2765 18914 2799
rect 18848 2731 18914 2765
rect 18848 2697 18864 2731
rect 18898 2697 18914 2731
rect 18848 2663 18914 2697
rect 18848 2629 18864 2663
rect 18898 2629 18914 2663
rect 18848 2595 18914 2629
rect 18848 2561 18864 2595
rect 18898 2561 18914 2595
rect 18848 2520 18914 2561
rect 18944 3479 19010 3520
rect 18944 3445 18960 3479
rect 18994 3445 19010 3479
rect 18944 3411 19010 3445
rect 18944 3377 18960 3411
rect 18994 3377 19010 3411
rect 18944 3343 19010 3377
rect 18944 3309 18960 3343
rect 18994 3309 19010 3343
rect 18944 3275 19010 3309
rect 18944 3241 18960 3275
rect 18994 3241 19010 3275
rect 18944 3207 19010 3241
rect 18944 3173 18960 3207
rect 18994 3173 19010 3207
rect 18944 3139 19010 3173
rect 18944 3105 18960 3139
rect 18994 3105 19010 3139
rect 18944 3071 19010 3105
rect 18944 3037 18960 3071
rect 18994 3037 19010 3071
rect 18944 3003 19010 3037
rect 18944 2969 18960 3003
rect 18994 2969 19010 3003
rect 18944 2935 19010 2969
rect 18944 2901 18960 2935
rect 18994 2901 19010 2935
rect 18944 2867 19010 2901
rect 18944 2833 18960 2867
rect 18994 2833 19010 2867
rect 18944 2799 19010 2833
rect 18944 2765 18960 2799
rect 18994 2765 19010 2799
rect 18944 2731 19010 2765
rect 18944 2697 18960 2731
rect 18994 2697 19010 2731
rect 18944 2663 19010 2697
rect 18944 2629 18960 2663
rect 18994 2629 19010 2663
rect 18944 2595 19010 2629
rect 18944 2561 18960 2595
rect 18994 2561 19010 2595
rect 18944 2520 19010 2561
rect 19040 3479 19106 3520
rect 19040 3445 19056 3479
rect 19090 3445 19106 3479
rect 19040 3411 19106 3445
rect 19040 3377 19056 3411
rect 19090 3377 19106 3411
rect 19040 3343 19106 3377
rect 19040 3309 19056 3343
rect 19090 3309 19106 3343
rect 19040 3275 19106 3309
rect 19040 3241 19056 3275
rect 19090 3241 19106 3275
rect 19040 3207 19106 3241
rect 19040 3173 19056 3207
rect 19090 3173 19106 3207
rect 19040 3139 19106 3173
rect 19040 3105 19056 3139
rect 19090 3105 19106 3139
rect 19040 3071 19106 3105
rect 19040 3037 19056 3071
rect 19090 3037 19106 3071
rect 19040 3003 19106 3037
rect 19040 2969 19056 3003
rect 19090 2969 19106 3003
rect 19040 2935 19106 2969
rect 19040 2901 19056 2935
rect 19090 2901 19106 2935
rect 19040 2867 19106 2901
rect 19040 2833 19056 2867
rect 19090 2833 19106 2867
rect 19040 2799 19106 2833
rect 19040 2765 19056 2799
rect 19090 2765 19106 2799
rect 19040 2731 19106 2765
rect 19040 2697 19056 2731
rect 19090 2697 19106 2731
rect 19040 2663 19106 2697
rect 19040 2629 19056 2663
rect 19090 2629 19106 2663
rect 19040 2595 19106 2629
rect 19040 2561 19056 2595
rect 19090 2561 19106 2595
rect 19040 2520 19106 2561
rect 19136 3479 19202 3520
rect 19136 3445 19152 3479
rect 19186 3445 19202 3479
rect 19136 3411 19202 3445
rect 19136 3377 19152 3411
rect 19186 3377 19202 3411
rect 19136 3343 19202 3377
rect 19136 3309 19152 3343
rect 19186 3309 19202 3343
rect 19136 3275 19202 3309
rect 19136 3241 19152 3275
rect 19186 3241 19202 3275
rect 19136 3207 19202 3241
rect 19136 3173 19152 3207
rect 19186 3173 19202 3207
rect 19136 3139 19202 3173
rect 19136 3105 19152 3139
rect 19186 3105 19202 3139
rect 19136 3071 19202 3105
rect 19136 3037 19152 3071
rect 19186 3037 19202 3071
rect 19136 3003 19202 3037
rect 19136 2969 19152 3003
rect 19186 2969 19202 3003
rect 19136 2935 19202 2969
rect 19136 2901 19152 2935
rect 19186 2901 19202 2935
rect 19136 2867 19202 2901
rect 19136 2833 19152 2867
rect 19186 2833 19202 2867
rect 19136 2799 19202 2833
rect 19136 2765 19152 2799
rect 19186 2765 19202 2799
rect 19136 2731 19202 2765
rect 19136 2697 19152 2731
rect 19186 2697 19202 2731
rect 19136 2663 19202 2697
rect 19136 2629 19152 2663
rect 19186 2629 19202 2663
rect 19136 2595 19202 2629
rect 19136 2561 19152 2595
rect 19186 2561 19202 2595
rect 19136 2520 19202 2561
rect 19232 3479 19298 3520
rect 19232 3445 19248 3479
rect 19282 3445 19298 3479
rect 19232 3411 19298 3445
rect 19232 3377 19248 3411
rect 19282 3377 19298 3411
rect 19232 3343 19298 3377
rect 19232 3309 19248 3343
rect 19282 3309 19298 3343
rect 19232 3275 19298 3309
rect 19232 3241 19248 3275
rect 19282 3241 19298 3275
rect 19232 3207 19298 3241
rect 19232 3173 19248 3207
rect 19282 3173 19298 3207
rect 19232 3139 19298 3173
rect 19232 3105 19248 3139
rect 19282 3105 19298 3139
rect 19232 3071 19298 3105
rect 19232 3037 19248 3071
rect 19282 3037 19298 3071
rect 19232 3003 19298 3037
rect 19232 2969 19248 3003
rect 19282 2969 19298 3003
rect 19232 2935 19298 2969
rect 19232 2901 19248 2935
rect 19282 2901 19298 2935
rect 19232 2867 19298 2901
rect 19232 2833 19248 2867
rect 19282 2833 19298 2867
rect 19232 2799 19298 2833
rect 19232 2765 19248 2799
rect 19282 2765 19298 2799
rect 19232 2731 19298 2765
rect 19232 2697 19248 2731
rect 19282 2697 19298 2731
rect 19232 2663 19298 2697
rect 19232 2629 19248 2663
rect 19282 2629 19298 2663
rect 19232 2595 19298 2629
rect 19232 2561 19248 2595
rect 19282 2561 19298 2595
rect 19232 2520 19298 2561
rect 19328 3479 19394 3520
rect 19328 3445 19344 3479
rect 19378 3445 19394 3479
rect 19328 3411 19394 3445
rect 19328 3377 19344 3411
rect 19378 3377 19394 3411
rect 19328 3343 19394 3377
rect 19328 3309 19344 3343
rect 19378 3309 19394 3343
rect 19328 3275 19394 3309
rect 19328 3241 19344 3275
rect 19378 3241 19394 3275
rect 19328 3207 19394 3241
rect 19328 3173 19344 3207
rect 19378 3173 19394 3207
rect 19328 3139 19394 3173
rect 19328 3105 19344 3139
rect 19378 3105 19394 3139
rect 19328 3071 19394 3105
rect 19328 3037 19344 3071
rect 19378 3037 19394 3071
rect 19328 3003 19394 3037
rect 19328 2969 19344 3003
rect 19378 2969 19394 3003
rect 19328 2935 19394 2969
rect 19328 2901 19344 2935
rect 19378 2901 19394 2935
rect 19328 2867 19394 2901
rect 19328 2833 19344 2867
rect 19378 2833 19394 2867
rect 19328 2799 19394 2833
rect 19328 2765 19344 2799
rect 19378 2765 19394 2799
rect 19328 2731 19394 2765
rect 19328 2697 19344 2731
rect 19378 2697 19394 2731
rect 19328 2663 19394 2697
rect 19328 2629 19344 2663
rect 19378 2629 19394 2663
rect 19328 2595 19394 2629
rect 19328 2561 19344 2595
rect 19378 2561 19394 2595
rect 19328 2520 19394 2561
rect 19424 3479 19490 3520
rect 19424 3445 19440 3479
rect 19474 3445 19490 3479
rect 19424 3411 19490 3445
rect 19424 3377 19440 3411
rect 19474 3377 19490 3411
rect 19424 3343 19490 3377
rect 19424 3309 19440 3343
rect 19474 3309 19490 3343
rect 19424 3275 19490 3309
rect 19424 3241 19440 3275
rect 19474 3241 19490 3275
rect 19424 3207 19490 3241
rect 19424 3173 19440 3207
rect 19474 3173 19490 3207
rect 19424 3139 19490 3173
rect 19424 3105 19440 3139
rect 19474 3105 19490 3139
rect 19424 3071 19490 3105
rect 19424 3037 19440 3071
rect 19474 3037 19490 3071
rect 19424 3003 19490 3037
rect 19424 2969 19440 3003
rect 19474 2969 19490 3003
rect 19424 2935 19490 2969
rect 19424 2901 19440 2935
rect 19474 2901 19490 2935
rect 19424 2867 19490 2901
rect 19424 2833 19440 2867
rect 19474 2833 19490 2867
rect 19424 2799 19490 2833
rect 19424 2765 19440 2799
rect 19474 2765 19490 2799
rect 19424 2731 19490 2765
rect 19424 2697 19440 2731
rect 19474 2697 19490 2731
rect 19424 2663 19490 2697
rect 19424 2629 19440 2663
rect 19474 2629 19490 2663
rect 19424 2595 19490 2629
rect 19424 2561 19440 2595
rect 19474 2561 19490 2595
rect 19424 2520 19490 2561
rect 19520 3479 19586 3520
rect 19520 3445 19536 3479
rect 19570 3445 19586 3479
rect 19520 3411 19586 3445
rect 19520 3377 19536 3411
rect 19570 3377 19586 3411
rect 19520 3343 19586 3377
rect 19520 3309 19536 3343
rect 19570 3309 19586 3343
rect 19520 3275 19586 3309
rect 19520 3241 19536 3275
rect 19570 3241 19586 3275
rect 19520 3207 19586 3241
rect 19520 3173 19536 3207
rect 19570 3173 19586 3207
rect 19520 3139 19586 3173
rect 19520 3105 19536 3139
rect 19570 3105 19586 3139
rect 19520 3071 19586 3105
rect 19520 3037 19536 3071
rect 19570 3037 19586 3071
rect 19520 3003 19586 3037
rect 19520 2969 19536 3003
rect 19570 2969 19586 3003
rect 19520 2935 19586 2969
rect 19520 2901 19536 2935
rect 19570 2901 19586 2935
rect 19520 2867 19586 2901
rect 19520 2833 19536 2867
rect 19570 2833 19586 2867
rect 19520 2799 19586 2833
rect 19520 2765 19536 2799
rect 19570 2765 19586 2799
rect 19520 2731 19586 2765
rect 19520 2697 19536 2731
rect 19570 2697 19586 2731
rect 19520 2663 19586 2697
rect 19520 2629 19536 2663
rect 19570 2629 19586 2663
rect 19520 2595 19586 2629
rect 19520 2561 19536 2595
rect 19570 2561 19586 2595
rect 19520 2520 19586 2561
rect 19616 3479 19682 3520
rect 19616 3445 19632 3479
rect 19666 3445 19682 3479
rect 19616 3411 19682 3445
rect 19616 3377 19632 3411
rect 19666 3377 19682 3411
rect 19616 3343 19682 3377
rect 19616 3309 19632 3343
rect 19666 3309 19682 3343
rect 19616 3275 19682 3309
rect 19616 3241 19632 3275
rect 19666 3241 19682 3275
rect 19616 3207 19682 3241
rect 19616 3173 19632 3207
rect 19666 3173 19682 3207
rect 19616 3139 19682 3173
rect 19616 3105 19632 3139
rect 19666 3105 19682 3139
rect 19616 3071 19682 3105
rect 19616 3037 19632 3071
rect 19666 3037 19682 3071
rect 19616 3003 19682 3037
rect 19616 2969 19632 3003
rect 19666 2969 19682 3003
rect 19616 2935 19682 2969
rect 19616 2901 19632 2935
rect 19666 2901 19682 2935
rect 19616 2867 19682 2901
rect 19616 2833 19632 2867
rect 19666 2833 19682 2867
rect 19616 2799 19682 2833
rect 19616 2765 19632 2799
rect 19666 2765 19682 2799
rect 19616 2731 19682 2765
rect 19616 2697 19632 2731
rect 19666 2697 19682 2731
rect 19616 2663 19682 2697
rect 19616 2629 19632 2663
rect 19666 2629 19682 2663
rect 19616 2595 19682 2629
rect 19616 2561 19632 2595
rect 19666 2561 19682 2595
rect 19616 2520 19682 2561
rect 19712 3479 19778 3520
rect 19712 3445 19728 3479
rect 19762 3445 19778 3479
rect 19712 3411 19778 3445
rect 19712 3377 19728 3411
rect 19762 3377 19778 3411
rect 19712 3343 19778 3377
rect 19712 3309 19728 3343
rect 19762 3309 19778 3343
rect 19712 3275 19778 3309
rect 19712 3241 19728 3275
rect 19762 3241 19778 3275
rect 19712 3207 19778 3241
rect 19712 3173 19728 3207
rect 19762 3173 19778 3207
rect 19712 3139 19778 3173
rect 19712 3105 19728 3139
rect 19762 3105 19778 3139
rect 19712 3071 19778 3105
rect 19712 3037 19728 3071
rect 19762 3037 19778 3071
rect 19712 3003 19778 3037
rect 19712 2969 19728 3003
rect 19762 2969 19778 3003
rect 19712 2935 19778 2969
rect 19712 2901 19728 2935
rect 19762 2901 19778 2935
rect 19712 2867 19778 2901
rect 19712 2833 19728 2867
rect 19762 2833 19778 2867
rect 19712 2799 19778 2833
rect 19712 2765 19728 2799
rect 19762 2765 19778 2799
rect 19712 2731 19778 2765
rect 19712 2697 19728 2731
rect 19762 2697 19778 2731
rect 19712 2663 19778 2697
rect 19712 2629 19728 2663
rect 19762 2629 19778 2663
rect 19712 2595 19778 2629
rect 19712 2561 19728 2595
rect 19762 2561 19778 2595
rect 19712 2520 19778 2561
rect 19808 3479 19874 3520
rect 19808 3445 19824 3479
rect 19858 3445 19874 3479
rect 19808 3411 19874 3445
rect 19808 3377 19824 3411
rect 19858 3377 19874 3411
rect 19808 3343 19874 3377
rect 19808 3309 19824 3343
rect 19858 3309 19874 3343
rect 19808 3275 19874 3309
rect 19808 3241 19824 3275
rect 19858 3241 19874 3275
rect 19808 3207 19874 3241
rect 19808 3173 19824 3207
rect 19858 3173 19874 3207
rect 19808 3139 19874 3173
rect 19808 3105 19824 3139
rect 19858 3105 19874 3139
rect 19808 3071 19874 3105
rect 19808 3037 19824 3071
rect 19858 3037 19874 3071
rect 19808 3003 19874 3037
rect 19808 2969 19824 3003
rect 19858 2969 19874 3003
rect 19808 2935 19874 2969
rect 19808 2901 19824 2935
rect 19858 2901 19874 2935
rect 19808 2867 19874 2901
rect 19808 2833 19824 2867
rect 19858 2833 19874 2867
rect 19808 2799 19874 2833
rect 19808 2765 19824 2799
rect 19858 2765 19874 2799
rect 19808 2731 19874 2765
rect 19808 2697 19824 2731
rect 19858 2697 19874 2731
rect 19808 2663 19874 2697
rect 19808 2629 19824 2663
rect 19858 2629 19874 2663
rect 19808 2595 19874 2629
rect 19808 2561 19824 2595
rect 19858 2561 19874 2595
rect 19808 2520 19874 2561
rect 19904 3479 19970 3520
rect 19904 3445 19920 3479
rect 19954 3445 19970 3479
rect 19904 3411 19970 3445
rect 19904 3377 19920 3411
rect 19954 3377 19970 3411
rect 19904 3343 19970 3377
rect 19904 3309 19920 3343
rect 19954 3309 19970 3343
rect 19904 3275 19970 3309
rect 19904 3241 19920 3275
rect 19954 3241 19970 3275
rect 19904 3207 19970 3241
rect 19904 3173 19920 3207
rect 19954 3173 19970 3207
rect 19904 3139 19970 3173
rect 19904 3105 19920 3139
rect 19954 3105 19970 3139
rect 19904 3071 19970 3105
rect 19904 3037 19920 3071
rect 19954 3037 19970 3071
rect 19904 3003 19970 3037
rect 19904 2969 19920 3003
rect 19954 2969 19970 3003
rect 19904 2935 19970 2969
rect 19904 2901 19920 2935
rect 19954 2901 19970 2935
rect 19904 2867 19970 2901
rect 19904 2833 19920 2867
rect 19954 2833 19970 2867
rect 19904 2799 19970 2833
rect 19904 2765 19920 2799
rect 19954 2765 19970 2799
rect 19904 2731 19970 2765
rect 19904 2697 19920 2731
rect 19954 2697 19970 2731
rect 19904 2663 19970 2697
rect 19904 2629 19920 2663
rect 19954 2629 19970 2663
rect 19904 2595 19970 2629
rect 19904 2561 19920 2595
rect 19954 2561 19970 2595
rect 19904 2520 19970 2561
rect 20000 3479 20062 3520
rect 20000 3445 20016 3479
rect 20050 3445 20062 3479
rect 20000 3411 20062 3445
rect 20000 3377 20016 3411
rect 20050 3377 20062 3411
rect 20000 3343 20062 3377
rect 20000 3309 20016 3343
rect 20050 3309 20062 3343
rect 20000 3275 20062 3309
rect 20000 3241 20016 3275
rect 20050 3241 20062 3275
rect 20000 3207 20062 3241
rect 20000 3173 20016 3207
rect 20050 3173 20062 3207
rect 20000 3139 20062 3173
rect 20000 3105 20016 3139
rect 20050 3105 20062 3139
rect 20000 3071 20062 3105
rect 20000 3037 20016 3071
rect 20050 3037 20062 3071
rect 20000 3003 20062 3037
rect 20000 2969 20016 3003
rect 20050 2969 20062 3003
rect 20000 2935 20062 2969
rect 20000 2901 20016 2935
rect 20050 2901 20062 2935
rect 20000 2867 20062 2901
rect 20000 2833 20016 2867
rect 20050 2833 20062 2867
rect 20000 2799 20062 2833
rect 20000 2765 20016 2799
rect 20050 2765 20062 2799
rect 20000 2731 20062 2765
rect 20000 2697 20016 2731
rect 20050 2697 20062 2731
rect 20000 2663 20062 2697
rect 20000 2629 20016 2663
rect 20050 2629 20062 2663
rect 20000 2595 20062 2629
rect 20000 2561 20016 2595
rect 20050 2561 20062 2595
rect 20000 2520 20062 2561
rect 20232 3487 20294 3528
rect 20232 3453 20244 3487
rect 20278 3453 20294 3487
rect 20232 3419 20294 3453
rect 20232 3385 20244 3419
rect 20278 3385 20294 3419
rect 20232 3351 20294 3385
rect 20232 3317 20244 3351
rect 20278 3317 20294 3351
rect 20232 3283 20294 3317
rect 20232 3249 20244 3283
rect 20278 3249 20294 3283
rect 20232 3215 20294 3249
rect 20232 3181 20244 3215
rect 20278 3181 20294 3215
rect 20232 3147 20294 3181
rect 20232 3113 20244 3147
rect 20278 3113 20294 3147
rect 20232 3079 20294 3113
rect 20232 3045 20244 3079
rect 20278 3045 20294 3079
rect 20232 3011 20294 3045
rect 20232 2977 20244 3011
rect 20278 2977 20294 3011
rect 20232 2943 20294 2977
rect 20232 2909 20244 2943
rect 20278 2909 20294 2943
rect 20232 2875 20294 2909
rect 20232 2841 20244 2875
rect 20278 2841 20294 2875
rect 20232 2807 20294 2841
rect 20232 2773 20244 2807
rect 20278 2773 20294 2807
rect 20232 2739 20294 2773
rect 20232 2705 20244 2739
rect 20278 2705 20294 2739
rect 20232 2671 20294 2705
rect 20232 2637 20244 2671
rect 20278 2637 20294 2671
rect 20232 2603 20294 2637
rect 20232 2569 20244 2603
rect 20278 2569 20294 2603
rect 20232 2528 20294 2569
rect 20324 3487 20390 3528
rect 20324 3453 20340 3487
rect 20374 3453 20390 3487
rect 20324 3419 20390 3453
rect 20324 3385 20340 3419
rect 20374 3385 20390 3419
rect 20324 3351 20390 3385
rect 20324 3317 20340 3351
rect 20374 3317 20390 3351
rect 20324 3283 20390 3317
rect 20324 3249 20340 3283
rect 20374 3249 20390 3283
rect 20324 3215 20390 3249
rect 20324 3181 20340 3215
rect 20374 3181 20390 3215
rect 20324 3147 20390 3181
rect 20324 3113 20340 3147
rect 20374 3113 20390 3147
rect 20324 3079 20390 3113
rect 20324 3045 20340 3079
rect 20374 3045 20390 3079
rect 20324 3011 20390 3045
rect 20324 2977 20340 3011
rect 20374 2977 20390 3011
rect 20324 2943 20390 2977
rect 20324 2909 20340 2943
rect 20374 2909 20390 2943
rect 20324 2875 20390 2909
rect 20324 2841 20340 2875
rect 20374 2841 20390 2875
rect 20324 2807 20390 2841
rect 20324 2773 20340 2807
rect 20374 2773 20390 2807
rect 20324 2739 20390 2773
rect 20324 2705 20340 2739
rect 20374 2705 20390 2739
rect 20324 2671 20390 2705
rect 20324 2637 20340 2671
rect 20374 2637 20390 2671
rect 20324 2603 20390 2637
rect 20324 2569 20340 2603
rect 20374 2569 20390 2603
rect 20324 2528 20390 2569
rect 20420 3487 20486 3528
rect 20420 3453 20436 3487
rect 20470 3453 20486 3487
rect 20420 3419 20486 3453
rect 20420 3385 20436 3419
rect 20470 3385 20486 3419
rect 20420 3351 20486 3385
rect 20420 3317 20436 3351
rect 20470 3317 20486 3351
rect 20420 3283 20486 3317
rect 20420 3249 20436 3283
rect 20470 3249 20486 3283
rect 20420 3215 20486 3249
rect 20420 3181 20436 3215
rect 20470 3181 20486 3215
rect 20420 3147 20486 3181
rect 20420 3113 20436 3147
rect 20470 3113 20486 3147
rect 20420 3079 20486 3113
rect 20420 3045 20436 3079
rect 20470 3045 20486 3079
rect 20420 3011 20486 3045
rect 20420 2977 20436 3011
rect 20470 2977 20486 3011
rect 20420 2943 20486 2977
rect 20420 2909 20436 2943
rect 20470 2909 20486 2943
rect 20420 2875 20486 2909
rect 20420 2841 20436 2875
rect 20470 2841 20486 2875
rect 20420 2807 20486 2841
rect 20420 2773 20436 2807
rect 20470 2773 20486 2807
rect 20420 2739 20486 2773
rect 20420 2705 20436 2739
rect 20470 2705 20486 2739
rect 20420 2671 20486 2705
rect 20420 2637 20436 2671
rect 20470 2637 20486 2671
rect 20420 2603 20486 2637
rect 20420 2569 20436 2603
rect 20470 2569 20486 2603
rect 20420 2528 20486 2569
rect 20516 3487 20582 3528
rect 20516 3453 20532 3487
rect 20566 3453 20582 3487
rect 20516 3419 20582 3453
rect 20516 3385 20532 3419
rect 20566 3385 20582 3419
rect 20516 3351 20582 3385
rect 20516 3317 20532 3351
rect 20566 3317 20582 3351
rect 20516 3283 20582 3317
rect 20516 3249 20532 3283
rect 20566 3249 20582 3283
rect 20516 3215 20582 3249
rect 20516 3181 20532 3215
rect 20566 3181 20582 3215
rect 20516 3147 20582 3181
rect 20516 3113 20532 3147
rect 20566 3113 20582 3147
rect 20516 3079 20582 3113
rect 20516 3045 20532 3079
rect 20566 3045 20582 3079
rect 20516 3011 20582 3045
rect 20516 2977 20532 3011
rect 20566 2977 20582 3011
rect 20516 2943 20582 2977
rect 20516 2909 20532 2943
rect 20566 2909 20582 2943
rect 20516 2875 20582 2909
rect 20516 2841 20532 2875
rect 20566 2841 20582 2875
rect 20516 2807 20582 2841
rect 20516 2773 20532 2807
rect 20566 2773 20582 2807
rect 20516 2739 20582 2773
rect 20516 2705 20532 2739
rect 20566 2705 20582 2739
rect 20516 2671 20582 2705
rect 20516 2637 20532 2671
rect 20566 2637 20582 2671
rect 20516 2603 20582 2637
rect 20516 2569 20532 2603
rect 20566 2569 20582 2603
rect 20516 2528 20582 2569
rect 20612 3487 20678 3528
rect 20612 3453 20628 3487
rect 20662 3453 20678 3487
rect 20612 3419 20678 3453
rect 20612 3385 20628 3419
rect 20662 3385 20678 3419
rect 20612 3351 20678 3385
rect 20612 3317 20628 3351
rect 20662 3317 20678 3351
rect 20612 3283 20678 3317
rect 20612 3249 20628 3283
rect 20662 3249 20678 3283
rect 20612 3215 20678 3249
rect 20612 3181 20628 3215
rect 20662 3181 20678 3215
rect 20612 3147 20678 3181
rect 20612 3113 20628 3147
rect 20662 3113 20678 3147
rect 20612 3079 20678 3113
rect 20612 3045 20628 3079
rect 20662 3045 20678 3079
rect 20612 3011 20678 3045
rect 20612 2977 20628 3011
rect 20662 2977 20678 3011
rect 20612 2943 20678 2977
rect 20612 2909 20628 2943
rect 20662 2909 20678 2943
rect 20612 2875 20678 2909
rect 20612 2841 20628 2875
rect 20662 2841 20678 2875
rect 20612 2807 20678 2841
rect 20612 2773 20628 2807
rect 20662 2773 20678 2807
rect 20612 2739 20678 2773
rect 20612 2705 20628 2739
rect 20662 2705 20678 2739
rect 20612 2671 20678 2705
rect 20612 2637 20628 2671
rect 20662 2637 20678 2671
rect 20612 2603 20678 2637
rect 20612 2569 20628 2603
rect 20662 2569 20678 2603
rect 20612 2528 20678 2569
rect 20708 3487 20774 3528
rect 20708 3453 20724 3487
rect 20758 3453 20774 3487
rect 20708 3419 20774 3453
rect 20708 3385 20724 3419
rect 20758 3385 20774 3419
rect 20708 3351 20774 3385
rect 20708 3317 20724 3351
rect 20758 3317 20774 3351
rect 20708 3283 20774 3317
rect 20708 3249 20724 3283
rect 20758 3249 20774 3283
rect 20708 3215 20774 3249
rect 20708 3181 20724 3215
rect 20758 3181 20774 3215
rect 20708 3147 20774 3181
rect 20708 3113 20724 3147
rect 20758 3113 20774 3147
rect 20708 3079 20774 3113
rect 20708 3045 20724 3079
rect 20758 3045 20774 3079
rect 20708 3011 20774 3045
rect 20708 2977 20724 3011
rect 20758 2977 20774 3011
rect 20708 2943 20774 2977
rect 20708 2909 20724 2943
rect 20758 2909 20774 2943
rect 20708 2875 20774 2909
rect 20708 2841 20724 2875
rect 20758 2841 20774 2875
rect 20708 2807 20774 2841
rect 20708 2773 20724 2807
rect 20758 2773 20774 2807
rect 20708 2739 20774 2773
rect 20708 2705 20724 2739
rect 20758 2705 20774 2739
rect 20708 2671 20774 2705
rect 20708 2637 20724 2671
rect 20758 2637 20774 2671
rect 20708 2603 20774 2637
rect 20708 2569 20724 2603
rect 20758 2569 20774 2603
rect 20708 2528 20774 2569
rect 20804 3487 20870 3528
rect 20804 3453 20820 3487
rect 20854 3453 20870 3487
rect 20804 3419 20870 3453
rect 20804 3385 20820 3419
rect 20854 3385 20870 3419
rect 20804 3351 20870 3385
rect 20804 3317 20820 3351
rect 20854 3317 20870 3351
rect 20804 3283 20870 3317
rect 20804 3249 20820 3283
rect 20854 3249 20870 3283
rect 20804 3215 20870 3249
rect 20804 3181 20820 3215
rect 20854 3181 20870 3215
rect 20804 3147 20870 3181
rect 20804 3113 20820 3147
rect 20854 3113 20870 3147
rect 20804 3079 20870 3113
rect 20804 3045 20820 3079
rect 20854 3045 20870 3079
rect 20804 3011 20870 3045
rect 20804 2977 20820 3011
rect 20854 2977 20870 3011
rect 20804 2943 20870 2977
rect 20804 2909 20820 2943
rect 20854 2909 20870 2943
rect 20804 2875 20870 2909
rect 20804 2841 20820 2875
rect 20854 2841 20870 2875
rect 20804 2807 20870 2841
rect 20804 2773 20820 2807
rect 20854 2773 20870 2807
rect 20804 2739 20870 2773
rect 20804 2705 20820 2739
rect 20854 2705 20870 2739
rect 20804 2671 20870 2705
rect 20804 2637 20820 2671
rect 20854 2637 20870 2671
rect 20804 2603 20870 2637
rect 20804 2569 20820 2603
rect 20854 2569 20870 2603
rect 20804 2528 20870 2569
rect 20900 3487 20966 3528
rect 20900 3453 20916 3487
rect 20950 3453 20966 3487
rect 20900 3419 20966 3453
rect 20900 3385 20916 3419
rect 20950 3385 20966 3419
rect 20900 3351 20966 3385
rect 20900 3317 20916 3351
rect 20950 3317 20966 3351
rect 20900 3283 20966 3317
rect 20900 3249 20916 3283
rect 20950 3249 20966 3283
rect 20900 3215 20966 3249
rect 20900 3181 20916 3215
rect 20950 3181 20966 3215
rect 20900 3147 20966 3181
rect 20900 3113 20916 3147
rect 20950 3113 20966 3147
rect 20900 3079 20966 3113
rect 20900 3045 20916 3079
rect 20950 3045 20966 3079
rect 20900 3011 20966 3045
rect 20900 2977 20916 3011
rect 20950 2977 20966 3011
rect 20900 2943 20966 2977
rect 20900 2909 20916 2943
rect 20950 2909 20966 2943
rect 20900 2875 20966 2909
rect 20900 2841 20916 2875
rect 20950 2841 20966 2875
rect 20900 2807 20966 2841
rect 20900 2773 20916 2807
rect 20950 2773 20966 2807
rect 20900 2739 20966 2773
rect 20900 2705 20916 2739
rect 20950 2705 20966 2739
rect 20900 2671 20966 2705
rect 20900 2637 20916 2671
rect 20950 2637 20966 2671
rect 20900 2603 20966 2637
rect 20900 2569 20916 2603
rect 20950 2569 20966 2603
rect 20900 2528 20966 2569
rect 20996 3487 21062 3528
rect 20996 3453 21012 3487
rect 21046 3453 21062 3487
rect 20996 3419 21062 3453
rect 20996 3385 21012 3419
rect 21046 3385 21062 3419
rect 20996 3351 21062 3385
rect 20996 3317 21012 3351
rect 21046 3317 21062 3351
rect 20996 3283 21062 3317
rect 20996 3249 21012 3283
rect 21046 3249 21062 3283
rect 20996 3215 21062 3249
rect 20996 3181 21012 3215
rect 21046 3181 21062 3215
rect 20996 3147 21062 3181
rect 20996 3113 21012 3147
rect 21046 3113 21062 3147
rect 20996 3079 21062 3113
rect 20996 3045 21012 3079
rect 21046 3045 21062 3079
rect 20996 3011 21062 3045
rect 20996 2977 21012 3011
rect 21046 2977 21062 3011
rect 20996 2943 21062 2977
rect 20996 2909 21012 2943
rect 21046 2909 21062 2943
rect 20996 2875 21062 2909
rect 20996 2841 21012 2875
rect 21046 2841 21062 2875
rect 20996 2807 21062 2841
rect 20996 2773 21012 2807
rect 21046 2773 21062 2807
rect 20996 2739 21062 2773
rect 20996 2705 21012 2739
rect 21046 2705 21062 2739
rect 20996 2671 21062 2705
rect 20996 2637 21012 2671
rect 21046 2637 21062 2671
rect 20996 2603 21062 2637
rect 20996 2569 21012 2603
rect 21046 2569 21062 2603
rect 20996 2528 21062 2569
rect 21092 3487 21158 3528
rect 21092 3453 21108 3487
rect 21142 3453 21158 3487
rect 21092 3419 21158 3453
rect 21092 3385 21108 3419
rect 21142 3385 21158 3419
rect 21092 3351 21158 3385
rect 21092 3317 21108 3351
rect 21142 3317 21158 3351
rect 21092 3283 21158 3317
rect 21092 3249 21108 3283
rect 21142 3249 21158 3283
rect 21092 3215 21158 3249
rect 21092 3181 21108 3215
rect 21142 3181 21158 3215
rect 21092 3147 21158 3181
rect 21092 3113 21108 3147
rect 21142 3113 21158 3147
rect 21092 3079 21158 3113
rect 21092 3045 21108 3079
rect 21142 3045 21158 3079
rect 21092 3011 21158 3045
rect 21092 2977 21108 3011
rect 21142 2977 21158 3011
rect 21092 2943 21158 2977
rect 21092 2909 21108 2943
rect 21142 2909 21158 2943
rect 21092 2875 21158 2909
rect 21092 2841 21108 2875
rect 21142 2841 21158 2875
rect 21092 2807 21158 2841
rect 21092 2773 21108 2807
rect 21142 2773 21158 2807
rect 21092 2739 21158 2773
rect 21092 2705 21108 2739
rect 21142 2705 21158 2739
rect 21092 2671 21158 2705
rect 21092 2637 21108 2671
rect 21142 2637 21158 2671
rect 21092 2603 21158 2637
rect 21092 2569 21108 2603
rect 21142 2569 21158 2603
rect 21092 2528 21158 2569
rect 21188 3487 21254 3528
rect 21188 3453 21204 3487
rect 21238 3453 21254 3487
rect 21188 3419 21254 3453
rect 21188 3385 21204 3419
rect 21238 3385 21254 3419
rect 21188 3351 21254 3385
rect 21188 3317 21204 3351
rect 21238 3317 21254 3351
rect 21188 3283 21254 3317
rect 21188 3249 21204 3283
rect 21238 3249 21254 3283
rect 21188 3215 21254 3249
rect 21188 3181 21204 3215
rect 21238 3181 21254 3215
rect 21188 3147 21254 3181
rect 21188 3113 21204 3147
rect 21238 3113 21254 3147
rect 21188 3079 21254 3113
rect 21188 3045 21204 3079
rect 21238 3045 21254 3079
rect 21188 3011 21254 3045
rect 21188 2977 21204 3011
rect 21238 2977 21254 3011
rect 21188 2943 21254 2977
rect 21188 2909 21204 2943
rect 21238 2909 21254 2943
rect 21188 2875 21254 2909
rect 21188 2841 21204 2875
rect 21238 2841 21254 2875
rect 21188 2807 21254 2841
rect 21188 2773 21204 2807
rect 21238 2773 21254 2807
rect 21188 2739 21254 2773
rect 21188 2705 21204 2739
rect 21238 2705 21254 2739
rect 21188 2671 21254 2705
rect 21188 2637 21204 2671
rect 21238 2637 21254 2671
rect 21188 2603 21254 2637
rect 21188 2569 21204 2603
rect 21238 2569 21254 2603
rect 21188 2528 21254 2569
rect 21284 3487 21350 3528
rect 21284 3453 21300 3487
rect 21334 3453 21350 3487
rect 21284 3419 21350 3453
rect 21284 3385 21300 3419
rect 21334 3385 21350 3419
rect 21284 3351 21350 3385
rect 21284 3317 21300 3351
rect 21334 3317 21350 3351
rect 21284 3283 21350 3317
rect 21284 3249 21300 3283
rect 21334 3249 21350 3283
rect 21284 3215 21350 3249
rect 21284 3181 21300 3215
rect 21334 3181 21350 3215
rect 21284 3147 21350 3181
rect 21284 3113 21300 3147
rect 21334 3113 21350 3147
rect 21284 3079 21350 3113
rect 21284 3045 21300 3079
rect 21334 3045 21350 3079
rect 21284 3011 21350 3045
rect 21284 2977 21300 3011
rect 21334 2977 21350 3011
rect 21284 2943 21350 2977
rect 21284 2909 21300 2943
rect 21334 2909 21350 2943
rect 21284 2875 21350 2909
rect 21284 2841 21300 2875
rect 21334 2841 21350 2875
rect 21284 2807 21350 2841
rect 21284 2773 21300 2807
rect 21334 2773 21350 2807
rect 21284 2739 21350 2773
rect 21284 2705 21300 2739
rect 21334 2705 21350 2739
rect 21284 2671 21350 2705
rect 21284 2637 21300 2671
rect 21334 2637 21350 2671
rect 21284 2603 21350 2637
rect 21284 2569 21300 2603
rect 21334 2569 21350 2603
rect 21284 2528 21350 2569
rect 21380 3487 21446 3528
rect 21380 3453 21396 3487
rect 21430 3453 21446 3487
rect 21380 3419 21446 3453
rect 21380 3385 21396 3419
rect 21430 3385 21446 3419
rect 21380 3351 21446 3385
rect 21380 3317 21396 3351
rect 21430 3317 21446 3351
rect 21380 3283 21446 3317
rect 21380 3249 21396 3283
rect 21430 3249 21446 3283
rect 21380 3215 21446 3249
rect 21380 3181 21396 3215
rect 21430 3181 21446 3215
rect 21380 3147 21446 3181
rect 21380 3113 21396 3147
rect 21430 3113 21446 3147
rect 21380 3079 21446 3113
rect 21380 3045 21396 3079
rect 21430 3045 21446 3079
rect 21380 3011 21446 3045
rect 21380 2977 21396 3011
rect 21430 2977 21446 3011
rect 21380 2943 21446 2977
rect 21380 2909 21396 2943
rect 21430 2909 21446 2943
rect 21380 2875 21446 2909
rect 21380 2841 21396 2875
rect 21430 2841 21446 2875
rect 21380 2807 21446 2841
rect 21380 2773 21396 2807
rect 21430 2773 21446 2807
rect 21380 2739 21446 2773
rect 21380 2705 21396 2739
rect 21430 2705 21446 2739
rect 21380 2671 21446 2705
rect 21380 2637 21396 2671
rect 21430 2637 21446 2671
rect 21380 2603 21446 2637
rect 21380 2569 21396 2603
rect 21430 2569 21446 2603
rect 21380 2528 21446 2569
rect 21476 3487 21542 3528
rect 21476 3453 21492 3487
rect 21526 3453 21542 3487
rect 21476 3419 21542 3453
rect 21476 3385 21492 3419
rect 21526 3385 21542 3419
rect 21476 3351 21542 3385
rect 21476 3317 21492 3351
rect 21526 3317 21542 3351
rect 21476 3283 21542 3317
rect 21476 3249 21492 3283
rect 21526 3249 21542 3283
rect 21476 3215 21542 3249
rect 21476 3181 21492 3215
rect 21526 3181 21542 3215
rect 21476 3147 21542 3181
rect 21476 3113 21492 3147
rect 21526 3113 21542 3147
rect 21476 3079 21542 3113
rect 21476 3045 21492 3079
rect 21526 3045 21542 3079
rect 21476 3011 21542 3045
rect 21476 2977 21492 3011
rect 21526 2977 21542 3011
rect 21476 2943 21542 2977
rect 21476 2909 21492 2943
rect 21526 2909 21542 2943
rect 21476 2875 21542 2909
rect 21476 2841 21492 2875
rect 21526 2841 21542 2875
rect 21476 2807 21542 2841
rect 21476 2773 21492 2807
rect 21526 2773 21542 2807
rect 21476 2739 21542 2773
rect 21476 2705 21492 2739
rect 21526 2705 21542 2739
rect 21476 2671 21542 2705
rect 21476 2637 21492 2671
rect 21526 2637 21542 2671
rect 21476 2603 21542 2637
rect 21476 2569 21492 2603
rect 21526 2569 21542 2603
rect 21476 2528 21542 2569
rect 21572 3487 21638 3528
rect 21572 3453 21588 3487
rect 21622 3453 21638 3487
rect 21572 3419 21638 3453
rect 21572 3385 21588 3419
rect 21622 3385 21638 3419
rect 21572 3351 21638 3385
rect 21572 3317 21588 3351
rect 21622 3317 21638 3351
rect 21572 3283 21638 3317
rect 21572 3249 21588 3283
rect 21622 3249 21638 3283
rect 21572 3215 21638 3249
rect 21572 3181 21588 3215
rect 21622 3181 21638 3215
rect 21572 3147 21638 3181
rect 21572 3113 21588 3147
rect 21622 3113 21638 3147
rect 21572 3079 21638 3113
rect 21572 3045 21588 3079
rect 21622 3045 21638 3079
rect 21572 3011 21638 3045
rect 21572 2977 21588 3011
rect 21622 2977 21638 3011
rect 21572 2943 21638 2977
rect 21572 2909 21588 2943
rect 21622 2909 21638 2943
rect 21572 2875 21638 2909
rect 21572 2841 21588 2875
rect 21622 2841 21638 2875
rect 21572 2807 21638 2841
rect 21572 2773 21588 2807
rect 21622 2773 21638 2807
rect 21572 2739 21638 2773
rect 21572 2705 21588 2739
rect 21622 2705 21638 2739
rect 21572 2671 21638 2705
rect 21572 2637 21588 2671
rect 21622 2637 21638 2671
rect 21572 2603 21638 2637
rect 21572 2569 21588 2603
rect 21622 2569 21638 2603
rect 21572 2528 21638 2569
rect 21668 3487 21734 3528
rect 21668 3453 21684 3487
rect 21718 3453 21734 3487
rect 21668 3419 21734 3453
rect 21668 3385 21684 3419
rect 21718 3385 21734 3419
rect 21668 3351 21734 3385
rect 21668 3317 21684 3351
rect 21718 3317 21734 3351
rect 21668 3283 21734 3317
rect 21668 3249 21684 3283
rect 21718 3249 21734 3283
rect 21668 3215 21734 3249
rect 21668 3181 21684 3215
rect 21718 3181 21734 3215
rect 21668 3147 21734 3181
rect 21668 3113 21684 3147
rect 21718 3113 21734 3147
rect 21668 3079 21734 3113
rect 21668 3045 21684 3079
rect 21718 3045 21734 3079
rect 21668 3011 21734 3045
rect 21668 2977 21684 3011
rect 21718 2977 21734 3011
rect 21668 2943 21734 2977
rect 21668 2909 21684 2943
rect 21718 2909 21734 2943
rect 21668 2875 21734 2909
rect 21668 2841 21684 2875
rect 21718 2841 21734 2875
rect 21668 2807 21734 2841
rect 21668 2773 21684 2807
rect 21718 2773 21734 2807
rect 21668 2739 21734 2773
rect 21668 2705 21684 2739
rect 21718 2705 21734 2739
rect 21668 2671 21734 2705
rect 21668 2637 21684 2671
rect 21718 2637 21734 2671
rect 21668 2603 21734 2637
rect 21668 2569 21684 2603
rect 21718 2569 21734 2603
rect 21668 2528 21734 2569
rect 21764 3487 21830 3528
rect 21764 3453 21780 3487
rect 21814 3453 21830 3487
rect 21764 3419 21830 3453
rect 21764 3385 21780 3419
rect 21814 3385 21830 3419
rect 21764 3351 21830 3385
rect 21764 3317 21780 3351
rect 21814 3317 21830 3351
rect 21764 3283 21830 3317
rect 21764 3249 21780 3283
rect 21814 3249 21830 3283
rect 21764 3215 21830 3249
rect 21764 3181 21780 3215
rect 21814 3181 21830 3215
rect 21764 3147 21830 3181
rect 21764 3113 21780 3147
rect 21814 3113 21830 3147
rect 21764 3079 21830 3113
rect 21764 3045 21780 3079
rect 21814 3045 21830 3079
rect 21764 3011 21830 3045
rect 21764 2977 21780 3011
rect 21814 2977 21830 3011
rect 21764 2943 21830 2977
rect 21764 2909 21780 2943
rect 21814 2909 21830 2943
rect 21764 2875 21830 2909
rect 21764 2841 21780 2875
rect 21814 2841 21830 2875
rect 21764 2807 21830 2841
rect 21764 2773 21780 2807
rect 21814 2773 21830 2807
rect 21764 2739 21830 2773
rect 21764 2705 21780 2739
rect 21814 2705 21830 2739
rect 21764 2671 21830 2705
rect 21764 2637 21780 2671
rect 21814 2637 21830 2671
rect 21764 2603 21830 2637
rect 21764 2569 21780 2603
rect 21814 2569 21830 2603
rect 21764 2528 21830 2569
rect 21860 3487 21926 3528
rect 21860 3453 21876 3487
rect 21910 3453 21926 3487
rect 21860 3419 21926 3453
rect 21860 3385 21876 3419
rect 21910 3385 21926 3419
rect 21860 3351 21926 3385
rect 21860 3317 21876 3351
rect 21910 3317 21926 3351
rect 21860 3283 21926 3317
rect 21860 3249 21876 3283
rect 21910 3249 21926 3283
rect 21860 3215 21926 3249
rect 21860 3181 21876 3215
rect 21910 3181 21926 3215
rect 21860 3147 21926 3181
rect 21860 3113 21876 3147
rect 21910 3113 21926 3147
rect 21860 3079 21926 3113
rect 21860 3045 21876 3079
rect 21910 3045 21926 3079
rect 21860 3011 21926 3045
rect 21860 2977 21876 3011
rect 21910 2977 21926 3011
rect 21860 2943 21926 2977
rect 21860 2909 21876 2943
rect 21910 2909 21926 2943
rect 21860 2875 21926 2909
rect 21860 2841 21876 2875
rect 21910 2841 21926 2875
rect 21860 2807 21926 2841
rect 21860 2773 21876 2807
rect 21910 2773 21926 2807
rect 21860 2739 21926 2773
rect 21860 2705 21876 2739
rect 21910 2705 21926 2739
rect 21860 2671 21926 2705
rect 21860 2637 21876 2671
rect 21910 2637 21926 2671
rect 21860 2603 21926 2637
rect 21860 2569 21876 2603
rect 21910 2569 21926 2603
rect 21860 2528 21926 2569
rect 21956 3487 22022 3528
rect 21956 3453 21972 3487
rect 22006 3453 22022 3487
rect 21956 3419 22022 3453
rect 21956 3385 21972 3419
rect 22006 3385 22022 3419
rect 21956 3351 22022 3385
rect 21956 3317 21972 3351
rect 22006 3317 22022 3351
rect 21956 3283 22022 3317
rect 21956 3249 21972 3283
rect 22006 3249 22022 3283
rect 21956 3215 22022 3249
rect 21956 3181 21972 3215
rect 22006 3181 22022 3215
rect 21956 3147 22022 3181
rect 21956 3113 21972 3147
rect 22006 3113 22022 3147
rect 21956 3079 22022 3113
rect 21956 3045 21972 3079
rect 22006 3045 22022 3079
rect 21956 3011 22022 3045
rect 21956 2977 21972 3011
rect 22006 2977 22022 3011
rect 21956 2943 22022 2977
rect 21956 2909 21972 2943
rect 22006 2909 22022 2943
rect 21956 2875 22022 2909
rect 21956 2841 21972 2875
rect 22006 2841 22022 2875
rect 21956 2807 22022 2841
rect 21956 2773 21972 2807
rect 22006 2773 22022 2807
rect 21956 2739 22022 2773
rect 21956 2705 21972 2739
rect 22006 2705 22022 2739
rect 21956 2671 22022 2705
rect 21956 2637 21972 2671
rect 22006 2637 22022 2671
rect 21956 2603 22022 2637
rect 21956 2569 21972 2603
rect 22006 2569 22022 2603
rect 21956 2528 22022 2569
rect 22052 3487 22118 3528
rect 22052 3453 22068 3487
rect 22102 3453 22118 3487
rect 22052 3419 22118 3453
rect 22052 3385 22068 3419
rect 22102 3385 22118 3419
rect 22052 3351 22118 3385
rect 22052 3317 22068 3351
rect 22102 3317 22118 3351
rect 22052 3283 22118 3317
rect 22052 3249 22068 3283
rect 22102 3249 22118 3283
rect 22052 3215 22118 3249
rect 22052 3181 22068 3215
rect 22102 3181 22118 3215
rect 22052 3147 22118 3181
rect 22052 3113 22068 3147
rect 22102 3113 22118 3147
rect 22052 3079 22118 3113
rect 22052 3045 22068 3079
rect 22102 3045 22118 3079
rect 22052 3011 22118 3045
rect 22052 2977 22068 3011
rect 22102 2977 22118 3011
rect 22052 2943 22118 2977
rect 22052 2909 22068 2943
rect 22102 2909 22118 2943
rect 22052 2875 22118 2909
rect 22052 2841 22068 2875
rect 22102 2841 22118 2875
rect 22052 2807 22118 2841
rect 22052 2773 22068 2807
rect 22102 2773 22118 2807
rect 22052 2739 22118 2773
rect 22052 2705 22068 2739
rect 22102 2705 22118 2739
rect 22052 2671 22118 2705
rect 22052 2637 22068 2671
rect 22102 2637 22118 2671
rect 22052 2603 22118 2637
rect 22052 2569 22068 2603
rect 22102 2569 22118 2603
rect 22052 2528 22118 2569
rect 22148 3487 22210 3528
rect 22148 3453 22164 3487
rect 22198 3453 22210 3487
rect 22148 3419 22210 3453
rect 22148 3385 22164 3419
rect 22198 3385 22210 3419
rect 22148 3351 22210 3385
rect 22148 3317 22164 3351
rect 22198 3317 22210 3351
rect 22148 3283 22210 3317
rect 22148 3249 22164 3283
rect 22198 3249 22210 3283
rect 22148 3215 22210 3249
rect 22148 3181 22164 3215
rect 22198 3181 22210 3215
rect 22148 3147 22210 3181
rect 22148 3113 22164 3147
rect 22198 3113 22210 3147
rect 22148 3079 22210 3113
rect 22148 3045 22164 3079
rect 22198 3045 22210 3079
rect 22148 3011 22210 3045
rect 22148 2977 22164 3011
rect 22198 2977 22210 3011
rect 22148 2943 22210 2977
rect 22148 2909 22164 2943
rect 22198 2909 22210 2943
rect 22148 2875 22210 2909
rect 22148 2841 22164 2875
rect 22198 2841 22210 2875
rect 22148 2807 22210 2841
rect 22148 2773 22164 2807
rect 22198 2773 22210 2807
rect 22148 2739 22210 2773
rect 22148 2705 22164 2739
rect 22198 2705 22210 2739
rect 22148 2671 22210 2705
rect 22148 2637 22164 2671
rect 22198 2637 22210 2671
rect 22148 2603 22210 2637
rect 22148 2569 22164 2603
rect 22198 2569 22210 2603
rect 22148 2528 22210 2569
rect 23162 3491 23224 3532
rect 23162 3457 23174 3491
rect 23208 3457 23224 3491
rect 23162 3423 23224 3457
rect 23162 3389 23174 3423
rect 23208 3389 23224 3423
rect 23162 3355 23224 3389
rect 23162 3321 23174 3355
rect 23208 3321 23224 3355
rect 23162 3287 23224 3321
rect 23162 3253 23174 3287
rect 23208 3253 23224 3287
rect 23162 3219 23224 3253
rect 23162 3185 23174 3219
rect 23208 3185 23224 3219
rect 23162 3151 23224 3185
rect 23162 3117 23174 3151
rect 23208 3117 23224 3151
rect 23162 3083 23224 3117
rect 23162 3049 23174 3083
rect 23208 3049 23224 3083
rect 23162 3015 23224 3049
rect 23162 2981 23174 3015
rect 23208 2981 23224 3015
rect 23162 2947 23224 2981
rect 23162 2913 23174 2947
rect 23208 2913 23224 2947
rect 23162 2879 23224 2913
rect 23162 2845 23174 2879
rect 23208 2845 23224 2879
rect 23162 2811 23224 2845
rect 23162 2777 23174 2811
rect 23208 2777 23224 2811
rect 23162 2743 23224 2777
rect 23162 2709 23174 2743
rect 23208 2709 23224 2743
rect 23162 2675 23224 2709
rect 23162 2641 23174 2675
rect 23208 2641 23224 2675
rect 23162 2607 23224 2641
rect 23162 2573 23174 2607
rect 23208 2573 23224 2607
rect 23162 2532 23224 2573
rect 23254 3491 23320 3532
rect 23254 3457 23270 3491
rect 23304 3457 23320 3491
rect 23254 3423 23320 3457
rect 23254 3389 23270 3423
rect 23304 3389 23320 3423
rect 23254 3355 23320 3389
rect 23254 3321 23270 3355
rect 23304 3321 23320 3355
rect 23254 3287 23320 3321
rect 23254 3253 23270 3287
rect 23304 3253 23320 3287
rect 23254 3219 23320 3253
rect 23254 3185 23270 3219
rect 23304 3185 23320 3219
rect 23254 3151 23320 3185
rect 23254 3117 23270 3151
rect 23304 3117 23320 3151
rect 23254 3083 23320 3117
rect 23254 3049 23270 3083
rect 23304 3049 23320 3083
rect 23254 3015 23320 3049
rect 23254 2981 23270 3015
rect 23304 2981 23320 3015
rect 23254 2947 23320 2981
rect 23254 2913 23270 2947
rect 23304 2913 23320 2947
rect 23254 2879 23320 2913
rect 23254 2845 23270 2879
rect 23304 2845 23320 2879
rect 23254 2811 23320 2845
rect 23254 2777 23270 2811
rect 23304 2777 23320 2811
rect 23254 2743 23320 2777
rect 23254 2709 23270 2743
rect 23304 2709 23320 2743
rect 23254 2675 23320 2709
rect 23254 2641 23270 2675
rect 23304 2641 23320 2675
rect 23254 2607 23320 2641
rect 23254 2573 23270 2607
rect 23304 2573 23320 2607
rect 23254 2532 23320 2573
rect 23350 3491 23416 3532
rect 23350 3457 23366 3491
rect 23400 3457 23416 3491
rect 23350 3423 23416 3457
rect 23350 3389 23366 3423
rect 23400 3389 23416 3423
rect 23350 3355 23416 3389
rect 23350 3321 23366 3355
rect 23400 3321 23416 3355
rect 23350 3287 23416 3321
rect 23350 3253 23366 3287
rect 23400 3253 23416 3287
rect 23350 3219 23416 3253
rect 23350 3185 23366 3219
rect 23400 3185 23416 3219
rect 23350 3151 23416 3185
rect 23350 3117 23366 3151
rect 23400 3117 23416 3151
rect 23350 3083 23416 3117
rect 23350 3049 23366 3083
rect 23400 3049 23416 3083
rect 23350 3015 23416 3049
rect 23350 2981 23366 3015
rect 23400 2981 23416 3015
rect 23350 2947 23416 2981
rect 23350 2913 23366 2947
rect 23400 2913 23416 2947
rect 23350 2879 23416 2913
rect 23350 2845 23366 2879
rect 23400 2845 23416 2879
rect 23350 2811 23416 2845
rect 23350 2777 23366 2811
rect 23400 2777 23416 2811
rect 23350 2743 23416 2777
rect 23350 2709 23366 2743
rect 23400 2709 23416 2743
rect 23350 2675 23416 2709
rect 23350 2641 23366 2675
rect 23400 2641 23416 2675
rect 23350 2607 23416 2641
rect 23350 2573 23366 2607
rect 23400 2573 23416 2607
rect 23350 2532 23416 2573
rect 23446 3491 23512 3532
rect 23446 3457 23462 3491
rect 23496 3457 23512 3491
rect 23446 3423 23512 3457
rect 23446 3389 23462 3423
rect 23496 3389 23512 3423
rect 23446 3355 23512 3389
rect 23446 3321 23462 3355
rect 23496 3321 23512 3355
rect 23446 3287 23512 3321
rect 23446 3253 23462 3287
rect 23496 3253 23512 3287
rect 23446 3219 23512 3253
rect 23446 3185 23462 3219
rect 23496 3185 23512 3219
rect 23446 3151 23512 3185
rect 23446 3117 23462 3151
rect 23496 3117 23512 3151
rect 23446 3083 23512 3117
rect 23446 3049 23462 3083
rect 23496 3049 23512 3083
rect 23446 3015 23512 3049
rect 23446 2981 23462 3015
rect 23496 2981 23512 3015
rect 23446 2947 23512 2981
rect 23446 2913 23462 2947
rect 23496 2913 23512 2947
rect 23446 2879 23512 2913
rect 23446 2845 23462 2879
rect 23496 2845 23512 2879
rect 23446 2811 23512 2845
rect 23446 2777 23462 2811
rect 23496 2777 23512 2811
rect 23446 2743 23512 2777
rect 23446 2709 23462 2743
rect 23496 2709 23512 2743
rect 23446 2675 23512 2709
rect 23446 2641 23462 2675
rect 23496 2641 23512 2675
rect 23446 2607 23512 2641
rect 23446 2573 23462 2607
rect 23496 2573 23512 2607
rect 23446 2532 23512 2573
rect 23542 3491 23608 3532
rect 23542 3457 23558 3491
rect 23592 3457 23608 3491
rect 23542 3423 23608 3457
rect 23542 3389 23558 3423
rect 23592 3389 23608 3423
rect 23542 3355 23608 3389
rect 23542 3321 23558 3355
rect 23592 3321 23608 3355
rect 23542 3287 23608 3321
rect 23542 3253 23558 3287
rect 23592 3253 23608 3287
rect 23542 3219 23608 3253
rect 23542 3185 23558 3219
rect 23592 3185 23608 3219
rect 23542 3151 23608 3185
rect 23542 3117 23558 3151
rect 23592 3117 23608 3151
rect 23542 3083 23608 3117
rect 23542 3049 23558 3083
rect 23592 3049 23608 3083
rect 23542 3015 23608 3049
rect 23542 2981 23558 3015
rect 23592 2981 23608 3015
rect 23542 2947 23608 2981
rect 23542 2913 23558 2947
rect 23592 2913 23608 2947
rect 23542 2879 23608 2913
rect 23542 2845 23558 2879
rect 23592 2845 23608 2879
rect 23542 2811 23608 2845
rect 23542 2777 23558 2811
rect 23592 2777 23608 2811
rect 23542 2743 23608 2777
rect 23542 2709 23558 2743
rect 23592 2709 23608 2743
rect 23542 2675 23608 2709
rect 23542 2641 23558 2675
rect 23592 2641 23608 2675
rect 23542 2607 23608 2641
rect 23542 2573 23558 2607
rect 23592 2573 23608 2607
rect 23542 2532 23608 2573
rect 23638 3491 23700 3532
rect 23638 3457 23654 3491
rect 23688 3457 23700 3491
rect 23638 3423 23700 3457
rect 23638 3389 23654 3423
rect 23688 3389 23700 3423
rect 23638 3355 23700 3389
rect 23638 3321 23654 3355
rect 23688 3321 23700 3355
rect 23638 3287 23700 3321
rect 23638 3253 23654 3287
rect 23688 3253 23700 3287
rect 23638 3219 23700 3253
rect 23638 3185 23654 3219
rect 23688 3185 23700 3219
rect 23638 3151 23700 3185
rect 23638 3117 23654 3151
rect 23688 3117 23700 3151
rect 23638 3083 23700 3117
rect 23638 3049 23654 3083
rect 23688 3049 23700 3083
rect 23638 3015 23700 3049
rect 23638 2981 23654 3015
rect 23688 2981 23700 3015
rect 23638 2947 23700 2981
rect 23638 2913 23654 2947
rect 23688 2913 23700 2947
rect 23638 2879 23700 2913
rect 23638 2845 23654 2879
rect 23688 2845 23700 2879
rect 23638 2811 23700 2845
rect 23638 2777 23654 2811
rect 23688 2777 23700 2811
rect 23638 2743 23700 2777
rect 23638 2709 23654 2743
rect 23688 2709 23700 2743
rect 23638 2675 23700 2709
rect 23638 2641 23654 2675
rect 23688 2641 23700 2675
rect 23638 2607 23700 2641
rect 23638 2573 23654 2607
rect 23688 2573 23700 2607
rect 23638 2532 23700 2573
rect 23854 3481 23916 3522
rect 23854 3447 23866 3481
rect 23900 3447 23916 3481
rect 23854 3413 23916 3447
rect 23854 3379 23866 3413
rect 23900 3379 23916 3413
rect 23854 3345 23916 3379
rect 23854 3311 23866 3345
rect 23900 3311 23916 3345
rect 23854 3277 23916 3311
rect 23854 3243 23866 3277
rect 23900 3243 23916 3277
rect 23854 3209 23916 3243
rect 23854 3175 23866 3209
rect 23900 3175 23916 3209
rect 23854 3141 23916 3175
rect 23854 3107 23866 3141
rect 23900 3107 23916 3141
rect 23854 3073 23916 3107
rect 23854 3039 23866 3073
rect 23900 3039 23916 3073
rect 23854 3005 23916 3039
rect 23854 2971 23866 3005
rect 23900 2971 23916 3005
rect 23854 2937 23916 2971
rect 23854 2903 23866 2937
rect 23900 2903 23916 2937
rect 23854 2869 23916 2903
rect 23854 2835 23866 2869
rect 23900 2835 23916 2869
rect 23854 2801 23916 2835
rect 23854 2767 23866 2801
rect 23900 2767 23916 2801
rect 23854 2733 23916 2767
rect 23854 2699 23866 2733
rect 23900 2699 23916 2733
rect 23854 2665 23916 2699
rect 23854 2631 23866 2665
rect 23900 2631 23916 2665
rect 23854 2597 23916 2631
rect 23854 2563 23866 2597
rect 23900 2563 23916 2597
rect 23854 2522 23916 2563
rect 23946 3481 24012 3522
rect 23946 3447 23962 3481
rect 23996 3447 24012 3481
rect 23946 3413 24012 3447
rect 23946 3379 23962 3413
rect 23996 3379 24012 3413
rect 23946 3345 24012 3379
rect 23946 3311 23962 3345
rect 23996 3311 24012 3345
rect 23946 3277 24012 3311
rect 23946 3243 23962 3277
rect 23996 3243 24012 3277
rect 23946 3209 24012 3243
rect 23946 3175 23962 3209
rect 23996 3175 24012 3209
rect 23946 3141 24012 3175
rect 23946 3107 23962 3141
rect 23996 3107 24012 3141
rect 23946 3073 24012 3107
rect 23946 3039 23962 3073
rect 23996 3039 24012 3073
rect 23946 3005 24012 3039
rect 23946 2971 23962 3005
rect 23996 2971 24012 3005
rect 23946 2937 24012 2971
rect 23946 2903 23962 2937
rect 23996 2903 24012 2937
rect 23946 2869 24012 2903
rect 23946 2835 23962 2869
rect 23996 2835 24012 2869
rect 23946 2801 24012 2835
rect 23946 2767 23962 2801
rect 23996 2767 24012 2801
rect 23946 2733 24012 2767
rect 23946 2699 23962 2733
rect 23996 2699 24012 2733
rect 23946 2665 24012 2699
rect 23946 2631 23962 2665
rect 23996 2631 24012 2665
rect 23946 2597 24012 2631
rect 23946 2563 23962 2597
rect 23996 2563 24012 2597
rect 23946 2522 24012 2563
rect 24042 3481 24108 3522
rect 24042 3447 24058 3481
rect 24092 3447 24108 3481
rect 24042 3413 24108 3447
rect 24042 3379 24058 3413
rect 24092 3379 24108 3413
rect 24042 3345 24108 3379
rect 24042 3311 24058 3345
rect 24092 3311 24108 3345
rect 24042 3277 24108 3311
rect 24042 3243 24058 3277
rect 24092 3243 24108 3277
rect 24042 3209 24108 3243
rect 24042 3175 24058 3209
rect 24092 3175 24108 3209
rect 24042 3141 24108 3175
rect 24042 3107 24058 3141
rect 24092 3107 24108 3141
rect 24042 3073 24108 3107
rect 24042 3039 24058 3073
rect 24092 3039 24108 3073
rect 24042 3005 24108 3039
rect 24042 2971 24058 3005
rect 24092 2971 24108 3005
rect 24042 2937 24108 2971
rect 24042 2903 24058 2937
rect 24092 2903 24108 2937
rect 24042 2869 24108 2903
rect 24042 2835 24058 2869
rect 24092 2835 24108 2869
rect 24042 2801 24108 2835
rect 24042 2767 24058 2801
rect 24092 2767 24108 2801
rect 24042 2733 24108 2767
rect 24042 2699 24058 2733
rect 24092 2699 24108 2733
rect 24042 2665 24108 2699
rect 24042 2631 24058 2665
rect 24092 2631 24108 2665
rect 24042 2597 24108 2631
rect 24042 2563 24058 2597
rect 24092 2563 24108 2597
rect 24042 2522 24108 2563
rect 24138 3481 24204 3522
rect 24138 3447 24154 3481
rect 24188 3447 24204 3481
rect 24138 3413 24204 3447
rect 24138 3379 24154 3413
rect 24188 3379 24204 3413
rect 24138 3345 24204 3379
rect 24138 3311 24154 3345
rect 24188 3311 24204 3345
rect 24138 3277 24204 3311
rect 24138 3243 24154 3277
rect 24188 3243 24204 3277
rect 24138 3209 24204 3243
rect 24138 3175 24154 3209
rect 24188 3175 24204 3209
rect 24138 3141 24204 3175
rect 24138 3107 24154 3141
rect 24188 3107 24204 3141
rect 24138 3073 24204 3107
rect 24138 3039 24154 3073
rect 24188 3039 24204 3073
rect 24138 3005 24204 3039
rect 24138 2971 24154 3005
rect 24188 2971 24204 3005
rect 24138 2937 24204 2971
rect 24138 2903 24154 2937
rect 24188 2903 24204 2937
rect 24138 2869 24204 2903
rect 24138 2835 24154 2869
rect 24188 2835 24204 2869
rect 24138 2801 24204 2835
rect 24138 2767 24154 2801
rect 24188 2767 24204 2801
rect 24138 2733 24204 2767
rect 24138 2699 24154 2733
rect 24188 2699 24204 2733
rect 24138 2665 24204 2699
rect 24138 2631 24154 2665
rect 24188 2631 24204 2665
rect 24138 2597 24204 2631
rect 24138 2563 24154 2597
rect 24188 2563 24204 2597
rect 24138 2522 24204 2563
rect 24234 3481 24300 3522
rect 24234 3447 24250 3481
rect 24284 3447 24300 3481
rect 24234 3413 24300 3447
rect 24234 3379 24250 3413
rect 24284 3379 24300 3413
rect 24234 3345 24300 3379
rect 24234 3311 24250 3345
rect 24284 3311 24300 3345
rect 24234 3277 24300 3311
rect 24234 3243 24250 3277
rect 24284 3243 24300 3277
rect 24234 3209 24300 3243
rect 24234 3175 24250 3209
rect 24284 3175 24300 3209
rect 24234 3141 24300 3175
rect 24234 3107 24250 3141
rect 24284 3107 24300 3141
rect 24234 3073 24300 3107
rect 24234 3039 24250 3073
rect 24284 3039 24300 3073
rect 24234 3005 24300 3039
rect 24234 2971 24250 3005
rect 24284 2971 24300 3005
rect 24234 2937 24300 2971
rect 24234 2903 24250 2937
rect 24284 2903 24300 2937
rect 24234 2869 24300 2903
rect 24234 2835 24250 2869
rect 24284 2835 24300 2869
rect 24234 2801 24300 2835
rect 24234 2767 24250 2801
rect 24284 2767 24300 2801
rect 24234 2733 24300 2767
rect 24234 2699 24250 2733
rect 24284 2699 24300 2733
rect 24234 2665 24300 2699
rect 24234 2631 24250 2665
rect 24284 2631 24300 2665
rect 24234 2597 24300 2631
rect 24234 2563 24250 2597
rect 24284 2563 24300 2597
rect 24234 2522 24300 2563
rect 24330 3481 24396 3522
rect 24330 3447 24346 3481
rect 24380 3447 24396 3481
rect 24330 3413 24396 3447
rect 24330 3379 24346 3413
rect 24380 3379 24396 3413
rect 24330 3345 24396 3379
rect 24330 3311 24346 3345
rect 24380 3311 24396 3345
rect 24330 3277 24396 3311
rect 24330 3243 24346 3277
rect 24380 3243 24396 3277
rect 24330 3209 24396 3243
rect 24330 3175 24346 3209
rect 24380 3175 24396 3209
rect 24330 3141 24396 3175
rect 24330 3107 24346 3141
rect 24380 3107 24396 3141
rect 24330 3073 24396 3107
rect 24330 3039 24346 3073
rect 24380 3039 24396 3073
rect 24330 3005 24396 3039
rect 24330 2971 24346 3005
rect 24380 2971 24396 3005
rect 24330 2937 24396 2971
rect 24330 2903 24346 2937
rect 24380 2903 24396 2937
rect 24330 2869 24396 2903
rect 24330 2835 24346 2869
rect 24380 2835 24396 2869
rect 24330 2801 24396 2835
rect 24330 2767 24346 2801
rect 24380 2767 24396 2801
rect 24330 2733 24396 2767
rect 24330 2699 24346 2733
rect 24380 2699 24396 2733
rect 24330 2665 24396 2699
rect 24330 2631 24346 2665
rect 24380 2631 24396 2665
rect 24330 2597 24396 2631
rect 24330 2563 24346 2597
rect 24380 2563 24396 2597
rect 24330 2522 24396 2563
rect 24426 3481 24492 3522
rect 24426 3447 24442 3481
rect 24476 3447 24492 3481
rect 24426 3413 24492 3447
rect 24426 3379 24442 3413
rect 24476 3379 24492 3413
rect 24426 3345 24492 3379
rect 24426 3311 24442 3345
rect 24476 3311 24492 3345
rect 24426 3277 24492 3311
rect 24426 3243 24442 3277
rect 24476 3243 24492 3277
rect 24426 3209 24492 3243
rect 24426 3175 24442 3209
rect 24476 3175 24492 3209
rect 24426 3141 24492 3175
rect 24426 3107 24442 3141
rect 24476 3107 24492 3141
rect 24426 3073 24492 3107
rect 24426 3039 24442 3073
rect 24476 3039 24492 3073
rect 24426 3005 24492 3039
rect 24426 2971 24442 3005
rect 24476 2971 24492 3005
rect 24426 2937 24492 2971
rect 24426 2903 24442 2937
rect 24476 2903 24492 2937
rect 24426 2869 24492 2903
rect 24426 2835 24442 2869
rect 24476 2835 24492 2869
rect 24426 2801 24492 2835
rect 24426 2767 24442 2801
rect 24476 2767 24492 2801
rect 24426 2733 24492 2767
rect 24426 2699 24442 2733
rect 24476 2699 24492 2733
rect 24426 2665 24492 2699
rect 24426 2631 24442 2665
rect 24476 2631 24492 2665
rect 24426 2597 24492 2631
rect 24426 2563 24442 2597
rect 24476 2563 24492 2597
rect 24426 2522 24492 2563
rect 24522 3481 24588 3522
rect 24522 3447 24538 3481
rect 24572 3447 24588 3481
rect 24522 3413 24588 3447
rect 24522 3379 24538 3413
rect 24572 3379 24588 3413
rect 24522 3345 24588 3379
rect 24522 3311 24538 3345
rect 24572 3311 24588 3345
rect 24522 3277 24588 3311
rect 24522 3243 24538 3277
rect 24572 3243 24588 3277
rect 24522 3209 24588 3243
rect 24522 3175 24538 3209
rect 24572 3175 24588 3209
rect 24522 3141 24588 3175
rect 24522 3107 24538 3141
rect 24572 3107 24588 3141
rect 24522 3073 24588 3107
rect 24522 3039 24538 3073
rect 24572 3039 24588 3073
rect 24522 3005 24588 3039
rect 24522 2971 24538 3005
rect 24572 2971 24588 3005
rect 24522 2937 24588 2971
rect 24522 2903 24538 2937
rect 24572 2903 24588 2937
rect 24522 2869 24588 2903
rect 24522 2835 24538 2869
rect 24572 2835 24588 2869
rect 24522 2801 24588 2835
rect 24522 2767 24538 2801
rect 24572 2767 24588 2801
rect 24522 2733 24588 2767
rect 24522 2699 24538 2733
rect 24572 2699 24588 2733
rect 24522 2665 24588 2699
rect 24522 2631 24538 2665
rect 24572 2631 24588 2665
rect 24522 2597 24588 2631
rect 24522 2563 24538 2597
rect 24572 2563 24588 2597
rect 24522 2522 24588 2563
rect 24618 3481 24684 3522
rect 24618 3447 24634 3481
rect 24668 3447 24684 3481
rect 24618 3413 24684 3447
rect 24618 3379 24634 3413
rect 24668 3379 24684 3413
rect 24618 3345 24684 3379
rect 24618 3311 24634 3345
rect 24668 3311 24684 3345
rect 24618 3277 24684 3311
rect 24618 3243 24634 3277
rect 24668 3243 24684 3277
rect 24618 3209 24684 3243
rect 24618 3175 24634 3209
rect 24668 3175 24684 3209
rect 24618 3141 24684 3175
rect 24618 3107 24634 3141
rect 24668 3107 24684 3141
rect 24618 3073 24684 3107
rect 24618 3039 24634 3073
rect 24668 3039 24684 3073
rect 24618 3005 24684 3039
rect 24618 2971 24634 3005
rect 24668 2971 24684 3005
rect 24618 2937 24684 2971
rect 24618 2903 24634 2937
rect 24668 2903 24684 2937
rect 24618 2869 24684 2903
rect 24618 2835 24634 2869
rect 24668 2835 24684 2869
rect 24618 2801 24684 2835
rect 24618 2767 24634 2801
rect 24668 2767 24684 2801
rect 24618 2733 24684 2767
rect 24618 2699 24634 2733
rect 24668 2699 24684 2733
rect 24618 2665 24684 2699
rect 24618 2631 24634 2665
rect 24668 2631 24684 2665
rect 24618 2597 24684 2631
rect 24618 2563 24634 2597
rect 24668 2563 24684 2597
rect 24618 2522 24684 2563
rect 24714 3481 24780 3522
rect 24714 3447 24730 3481
rect 24764 3447 24780 3481
rect 24714 3413 24780 3447
rect 24714 3379 24730 3413
rect 24764 3379 24780 3413
rect 24714 3345 24780 3379
rect 24714 3311 24730 3345
rect 24764 3311 24780 3345
rect 24714 3277 24780 3311
rect 24714 3243 24730 3277
rect 24764 3243 24780 3277
rect 24714 3209 24780 3243
rect 24714 3175 24730 3209
rect 24764 3175 24780 3209
rect 24714 3141 24780 3175
rect 24714 3107 24730 3141
rect 24764 3107 24780 3141
rect 24714 3073 24780 3107
rect 24714 3039 24730 3073
rect 24764 3039 24780 3073
rect 24714 3005 24780 3039
rect 24714 2971 24730 3005
rect 24764 2971 24780 3005
rect 24714 2937 24780 2971
rect 24714 2903 24730 2937
rect 24764 2903 24780 2937
rect 24714 2869 24780 2903
rect 24714 2835 24730 2869
rect 24764 2835 24780 2869
rect 24714 2801 24780 2835
rect 24714 2767 24730 2801
rect 24764 2767 24780 2801
rect 24714 2733 24780 2767
rect 24714 2699 24730 2733
rect 24764 2699 24780 2733
rect 24714 2665 24780 2699
rect 24714 2631 24730 2665
rect 24764 2631 24780 2665
rect 24714 2597 24780 2631
rect 24714 2563 24730 2597
rect 24764 2563 24780 2597
rect 24714 2522 24780 2563
rect 24810 3481 24872 3522
rect 24810 3447 24826 3481
rect 24860 3447 24872 3481
rect 24810 3413 24872 3447
rect 24810 3379 24826 3413
rect 24860 3379 24872 3413
rect 24810 3345 24872 3379
rect 24810 3311 24826 3345
rect 24860 3311 24872 3345
rect 24810 3277 24872 3311
rect 24810 3243 24826 3277
rect 24860 3243 24872 3277
rect 24810 3209 24872 3243
rect 24810 3175 24826 3209
rect 24860 3175 24872 3209
rect 24810 3141 24872 3175
rect 24810 3107 24826 3141
rect 24860 3107 24872 3141
rect 24810 3073 24872 3107
rect 24810 3039 24826 3073
rect 24860 3039 24872 3073
rect 24810 3005 24872 3039
rect 24810 2971 24826 3005
rect 24860 2971 24872 3005
rect 24810 2937 24872 2971
rect 24810 2903 24826 2937
rect 24860 2903 24872 2937
rect 24810 2869 24872 2903
rect 24810 2835 24826 2869
rect 24860 2835 24872 2869
rect 24810 2801 24872 2835
rect 24810 2767 24826 2801
rect 24860 2767 24872 2801
rect 24810 2733 24872 2767
rect 24810 2699 24826 2733
rect 24860 2699 24872 2733
rect 24810 2665 24872 2699
rect 24810 2631 24826 2665
rect 24860 2631 24872 2665
rect 24810 2597 24872 2631
rect 24810 2563 24826 2597
rect 24860 2563 24872 2597
rect 24810 2522 24872 2563
rect 25052 3477 25114 3518
rect 25052 3443 25064 3477
rect 25098 3443 25114 3477
rect 25052 3409 25114 3443
rect 25052 3375 25064 3409
rect 25098 3375 25114 3409
rect 25052 3341 25114 3375
rect 25052 3307 25064 3341
rect 25098 3307 25114 3341
rect 25052 3273 25114 3307
rect 25052 3239 25064 3273
rect 25098 3239 25114 3273
rect 25052 3205 25114 3239
rect 25052 3171 25064 3205
rect 25098 3171 25114 3205
rect 25052 3137 25114 3171
rect 25052 3103 25064 3137
rect 25098 3103 25114 3137
rect 25052 3069 25114 3103
rect 25052 3035 25064 3069
rect 25098 3035 25114 3069
rect 25052 3001 25114 3035
rect 25052 2967 25064 3001
rect 25098 2967 25114 3001
rect 25052 2933 25114 2967
rect 25052 2899 25064 2933
rect 25098 2899 25114 2933
rect 25052 2865 25114 2899
rect 25052 2831 25064 2865
rect 25098 2831 25114 2865
rect 25052 2797 25114 2831
rect 25052 2763 25064 2797
rect 25098 2763 25114 2797
rect 25052 2729 25114 2763
rect 25052 2695 25064 2729
rect 25098 2695 25114 2729
rect 25052 2661 25114 2695
rect 25052 2627 25064 2661
rect 25098 2627 25114 2661
rect 25052 2593 25114 2627
rect 25052 2559 25064 2593
rect 25098 2559 25114 2593
rect 25052 2518 25114 2559
rect 25144 3477 25210 3518
rect 25144 3443 25160 3477
rect 25194 3443 25210 3477
rect 25144 3409 25210 3443
rect 25144 3375 25160 3409
rect 25194 3375 25210 3409
rect 25144 3341 25210 3375
rect 25144 3307 25160 3341
rect 25194 3307 25210 3341
rect 25144 3273 25210 3307
rect 25144 3239 25160 3273
rect 25194 3239 25210 3273
rect 25144 3205 25210 3239
rect 25144 3171 25160 3205
rect 25194 3171 25210 3205
rect 25144 3137 25210 3171
rect 25144 3103 25160 3137
rect 25194 3103 25210 3137
rect 25144 3069 25210 3103
rect 25144 3035 25160 3069
rect 25194 3035 25210 3069
rect 25144 3001 25210 3035
rect 25144 2967 25160 3001
rect 25194 2967 25210 3001
rect 25144 2933 25210 2967
rect 25144 2899 25160 2933
rect 25194 2899 25210 2933
rect 25144 2865 25210 2899
rect 25144 2831 25160 2865
rect 25194 2831 25210 2865
rect 25144 2797 25210 2831
rect 25144 2763 25160 2797
rect 25194 2763 25210 2797
rect 25144 2729 25210 2763
rect 25144 2695 25160 2729
rect 25194 2695 25210 2729
rect 25144 2661 25210 2695
rect 25144 2627 25160 2661
rect 25194 2627 25210 2661
rect 25144 2593 25210 2627
rect 25144 2559 25160 2593
rect 25194 2559 25210 2593
rect 25144 2518 25210 2559
rect 25240 3477 25306 3518
rect 25240 3443 25256 3477
rect 25290 3443 25306 3477
rect 25240 3409 25306 3443
rect 25240 3375 25256 3409
rect 25290 3375 25306 3409
rect 25240 3341 25306 3375
rect 25240 3307 25256 3341
rect 25290 3307 25306 3341
rect 25240 3273 25306 3307
rect 25240 3239 25256 3273
rect 25290 3239 25306 3273
rect 25240 3205 25306 3239
rect 25240 3171 25256 3205
rect 25290 3171 25306 3205
rect 25240 3137 25306 3171
rect 25240 3103 25256 3137
rect 25290 3103 25306 3137
rect 25240 3069 25306 3103
rect 25240 3035 25256 3069
rect 25290 3035 25306 3069
rect 25240 3001 25306 3035
rect 25240 2967 25256 3001
rect 25290 2967 25306 3001
rect 25240 2933 25306 2967
rect 25240 2899 25256 2933
rect 25290 2899 25306 2933
rect 25240 2865 25306 2899
rect 25240 2831 25256 2865
rect 25290 2831 25306 2865
rect 25240 2797 25306 2831
rect 25240 2763 25256 2797
rect 25290 2763 25306 2797
rect 25240 2729 25306 2763
rect 25240 2695 25256 2729
rect 25290 2695 25306 2729
rect 25240 2661 25306 2695
rect 25240 2627 25256 2661
rect 25290 2627 25306 2661
rect 25240 2593 25306 2627
rect 25240 2559 25256 2593
rect 25290 2559 25306 2593
rect 25240 2518 25306 2559
rect 25336 3477 25402 3518
rect 25336 3443 25352 3477
rect 25386 3443 25402 3477
rect 25336 3409 25402 3443
rect 25336 3375 25352 3409
rect 25386 3375 25402 3409
rect 25336 3341 25402 3375
rect 25336 3307 25352 3341
rect 25386 3307 25402 3341
rect 25336 3273 25402 3307
rect 25336 3239 25352 3273
rect 25386 3239 25402 3273
rect 25336 3205 25402 3239
rect 25336 3171 25352 3205
rect 25386 3171 25402 3205
rect 25336 3137 25402 3171
rect 25336 3103 25352 3137
rect 25386 3103 25402 3137
rect 25336 3069 25402 3103
rect 25336 3035 25352 3069
rect 25386 3035 25402 3069
rect 25336 3001 25402 3035
rect 25336 2967 25352 3001
rect 25386 2967 25402 3001
rect 25336 2933 25402 2967
rect 25336 2899 25352 2933
rect 25386 2899 25402 2933
rect 25336 2865 25402 2899
rect 25336 2831 25352 2865
rect 25386 2831 25402 2865
rect 25336 2797 25402 2831
rect 25336 2763 25352 2797
rect 25386 2763 25402 2797
rect 25336 2729 25402 2763
rect 25336 2695 25352 2729
rect 25386 2695 25402 2729
rect 25336 2661 25402 2695
rect 25336 2627 25352 2661
rect 25386 2627 25402 2661
rect 25336 2593 25402 2627
rect 25336 2559 25352 2593
rect 25386 2559 25402 2593
rect 25336 2518 25402 2559
rect 25432 3477 25498 3518
rect 25432 3443 25448 3477
rect 25482 3443 25498 3477
rect 25432 3409 25498 3443
rect 25432 3375 25448 3409
rect 25482 3375 25498 3409
rect 25432 3341 25498 3375
rect 25432 3307 25448 3341
rect 25482 3307 25498 3341
rect 25432 3273 25498 3307
rect 25432 3239 25448 3273
rect 25482 3239 25498 3273
rect 25432 3205 25498 3239
rect 25432 3171 25448 3205
rect 25482 3171 25498 3205
rect 25432 3137 25498 3171
rect 25432 3103 25448 3137
rect 25482 3103 25498 3137
rect 25432 3069 25498 3103
rect 25432 3035 25448 3069
rect 25482 3035 25498 3069
rect 25432 3001 25498 3035
rect 25432 2967 25448 3001
rect 25482 2967 25498 3001
rect 25432 2933 25498 2967
rect 25432 2899 25448 2933
rect 25482 2899 25498 2933
rect 25432 2865 25498 2899
rect 25432 2831 25448 2865
rect 25482 2831 25498 2865
rect 25432 2797 25498 2831
rect 25432 2763 25448 2797
rect 25482 2763 25498 2797
rect 25432 2729 25498 2763
rect 25432 2695 25448 2729
rect 25482 2695 25498 2729
rect 25432 2661 25498 2695
rect 25432 2627 25448 2661
rect 25482 2627 25498 2661
rect 25432 2593 25498 2627
rect 25432 2559 25448 2593
rect 25482 2559 25498 2593
rect 25432 2518 25498 2559
rect 25528 3477 25594 3518
rect 25528 3443 25544 3477
rect 25578 3443 25594 3477
rect 25528 3409 25594 3443
rect 25528 3375 25544 3409
rect 25578 3375 25594 3409
rect 25528 3341 25594 3375
rect 25528 3307 25544 3341
rect 25578 3307 25594 3341
rect 25528 3273 25594 3307
rect 25528 3239 25544 3273
rect 25578 3239 25594 3273
rect 25528 3205 25594 3239
rect 25528 3171 25544 3205
rect 25578 3171 25594 3205
rect 25528 3137 25594 3171
rect 25528 3103 25544 3137
rect 25578 3103 25594 3137
rect 25528 3069 25594 3103
rect 25528 3035 25544 3069
rect 25578 3035 25594 3069
rect 25528 3001 25594 3035
rect 25528 2967 25544 3001
rect 25578 2967 25594 3001
rect 25528 2933 25594 2967
rect 25528 2899 25544 2933
rect 25578 2899 25594 2933
rect 25528 2865 25594 2899
rect 25528 2831 25544 2865
rect 25578 2831 25594 2865
rect 25528 2797 25594 2831
rect 25528 2763 25544 2797
rect 25578 2763 25594 2797
rect 25528 2729 25594 2763
rect 25528 2695 25544 2729
rect 25578 2695 25594 2729
rect 25528 2661 25594 2695
rect 25528 2627 25544 2661
rect 25578 2627 25594 2661
rect 25528 2593 25594 2627
rect 25528 2559 25544 2593
rect 25578 2559 25594 2593
rect 25528 2518 25594 2559
rect 25624 3477 25690 3518
rect 25624 3443 25640 3477
rect 25674 3443 25690 3477
rect 25624 3409 25690 3443
rect 25624 3375 25640 3409
rect 25674 3375 25690 3409
rect 25624 3341 25690 3375
rect 25624 3307 25640 3341
rect 25674 3307 25690 3341
rect 25624 3273 25690 3307
rect 25624 3239 25640 3273
rect 25674 3239 25690 3273
rect 25624 3205 25690 3239
rect 25624 3171 25640 3205
rect 25674 3171 25690 3205
rect 25624 3137 25690 3171
rect 25624 3103 25640 3137
rect 25674 3103 25690 3137
rect 25624 3069 25690 3103
rect 25624 3035 25640 3069
rect 25674 3035 25690 3069
rect 25624 3001 25690 3035
rect 25624 2967 25640 3001
rect 25674 2967 25690 3001
rect 25624 2933 25690 2967
rect 25624 2899 25640 2933
rect 25674 2899 25690 2933
rect 25624 2865 25690 2899
rect 25624 2831 25640 2865
rect 25674 2831 25690 2865
rect 25624 2797 25690 2831
rect 25624 2763 25640 2797
rect 25674 2763 25690 2797
rect 25624 2729 25690 2763
rect 25624 2695 25640 2729
rect 25674 2695 25690 2729
rect 25624 2661 25690 2695
rect 25624 2627 25640 2661
rect 25674 2627 25690 2661
rect 25624 2593 25690 2627
rect 25624 2559 25640 2593
rect 25674 2559 25690 2593
rect 25624 2518 25690 2559
rect 25720 3477 25786 3518
rect 25720 3443 25736 3477
rect 25770 3443 25786 3477
rect 25720 3409 25786 3443
rect 25720 3375 25736 3409
rect 25770 3375 25786 3409
rect 25720 3341 25786 3375
rect 25720 3307 25736 3341
rect 25770 3307 25786 3341
rect 25720 3273 25786 3307
rect 25720 3239 25736 3273
rect 25770 3239 25786 3273
rect 25720 3205 25786 3239
rect 25720 3171 25736 3205
rect 25770 3171 25786 3205
rect 25720 3137 25786 3171
rect 25720 3103 25736 3137
rect 25770 3103 25786 3137
rect 25720 3069 25786 3103
rect 25720 3035 25736 3069
rect 25770 3035 25786 3069
rect 25720 3001 25786 3035
rect 25720 2967 25736 3001
rect 25770 2967 25786 3001
rect 25720 2933 25786 2967
rect 25720 2899 25736 2933
rect 25770 2899 25786 2933
rect 25720 2865 25786 2899
rect 25720 2831 25736 2865
rect 25770 2831 25786 2865
rect 25720 2797 25786 2831
rect 25720 2763 25736 2797
rect 25770 2763 25786 2797
rect 25720 2729 25786 2763
rect 25720 2695 25736 2729
rect 25770 2695 25786 2729
rect 25720 2661 25786 2695
rect 25720 2627 25736 2661
rect 25770 2627 25786 2661
rect 25720 2593 25786 2627
rect 25720 2559 25736 2593
rect 25770 2559 25786 2593
rect 25720 2518 25786 2559
rect 25816 3477 25882 3518
rect 25816 3443 25832 3477
rect 25866 3443 25882 3477
rect 25816 3409 25882 3443
rect 25816 3375 25832 3409
rect 25866 3375 25882 3409
rect 25816 3341 25882 3375
rect 25816 3307 25832 3341
rect 25866 3307 25882 3341
rect 25816 3273 25882 3307
rect 25816 3239 25832 3273
rect 25866 3239 25882 3273
rect 25816 3205 25882 3239
rect 25816 3171 25832 3205
rect 25866 3171 25882 3205
rect 25816 3137 25882 3171
rect 25816 3103 25832 3137
rect 25866 3103 25882 3137
rect 25816 3069 25882 3103
rect 25816 3035 25832 3069
rect 25866 3035 25882 3069
rect 25816 3001 25882 3035
rect 25816 2967 25832 3001
rect 25866 2967 25882 3001
rect 25816 2933 25882 2967
rect 25816 2899 25832 2933
rect 25866 2899 25882 2933
rect 25816 2865 25882 2899
rect 25816 2831 25832 2865
rect 25866 2831 25882 2865
rect 25816 2797 25882 2831
rect 25816 2763 25832 2797
rect 25866 2763 25882 2797
rect 25816 2729 25882 2763
rect 25816 2695 25832 2729
rect 25866 2695 25882 2729
rect 25816 2661 25882 2695
rect 25816 2627 25832 2661
rect 25866 2627 25882 2661
rect 25816 2593 25882 2627
rect 25816 2559 25832 2593
rect 25866 2559 25882 2593
rect 25816 2518 25882 2559
rect 25912 3477 25978 3518
rect 25912 3443 25928 3477
rect 25962 3443 25978 3477
rect 25912 3409 25978 3443
rect 25912 3375 25928 3409
rect 25962 3375 25978 3409
rect 25912 3341 25978 3375
rect 25912 3307 25928 3341
rect 25962 3307 25978 3341
rect 25912 3273 25978 3307
rect 25912 3239 25928 3273
rect 25962 3239 25978 3273
rect 25912 3205 25978 3239
rect 25912 3171 25928 3205
rect 25962 3171 25978 3205
rect 25912 3137 25978 3171
rect 25912 3103 25928 3137
rect 25962 3103 25978 3137
rect 25912 3069 25978 3103
rect 25912 3035 25928 3069
rect 25962 3035 25978 3069
rect 25912 3001 25978 3035
rect 25912 2967 25928 3001
rect 25962 2967 25978 3001
rect 25912 2933 25978 2967
rect 25912 2899 25928 2933
rect 25962 2899 25978 2933
rect 25912 2865 25978 2899
rect 25912 2831 25928 2865
rect 25962 2831 25978 2865
rect 25912 2797 25978 2831
rect 25912 2763 25928 2797
rect 25962 2763 25978 2797
rect 25912 2729 25978 2763
rect 25912 2695 25928 2729
rect 25962 2695 25978 2729
rect 25912 2661 25978 2695
rect 25912 2627 25928 2661
rect 25962 2627 25978 2661
rect 25912 2593 25978 2627
rect 25912 2559 25928 2593
rect 25962 2559 25978 2593
rect 25912 2518 25978 2559
rect 26008 3477 26074 3518
rect 26008 3443 26024 3477
rect 26058 3443 26074 3477
rect 26008 3409 26074 3443
rect 26008 3375 26024 3409
rect 26058 3375 26074 3409
rect 26008 3341 26074 3375
rect 26008 3307 26024 3341
rect 26058 3307 26074 3341
rect 26008 3273 26074 3307
rect 26008 3239 26024 3273
rect 26058 3239 26074 3273
rect 26008 3205 26074 3239
rect 26008 3171 26024 3205
rect 26058 3171 26074 3205
rect 26008 3137 26074 3171
rect 26008 3103 26024 3137
rect 26058 3103 26074 3137
rect 26008 3069 26074 3103
rect 26008 3035 26024 3069
rect 26058 3035 26074 3069
rect 26008 3001 26074 3035
rect 26008 2967 26024 3001
rect 26058 2967 26074 3001
rect 26008 2933 26074 2967
rect 26008 2899 26024 2933
rect 26058 2899 26074 2933
rect 26008 2865 26074 2899
rect 26008 2831 26024 2865
rect 26058 2831 26074 2865
rect 26008 2797 26074 2831
rect 26008 2763 26024 2797
rect 26058 2763 26074 2797
rect 26008 2729 26074 2763
rect 26008 2695 26024 2729
rect 26058 2695 26074 2729
rect 26008 2661 26074 2695
rect 26008 2627 26024 2661
rect 26058 2627 26074 2661
rect 26008 2593 26074 2627
rect 26008 2559 26024 2593
rect 26058 2559 26074 2593
rect 26008 2518 26074 2559
rect 26104 3477 26170 3518
rect 26104 3443 26120 3477
rect 26154 3443 26170 3477
rect 26104 3409 26170 3443
rect 26104 3375 26120 3409
rect 26154 3375 26170 3409
rect 26104 3341 26170 3375
rect 26104 3307 26120 3341
rect 26154 3307 26170 3341
rect 26104 3273 26170 3307
rect 26104 3239 26120 3273
rect 26154 3239 26170 3273
rect 26104 3205 26170 3239
rect 26104 3171 26120 3205
rect 26154 3171 26170 3205
rect 26104 3137 26170 3171
rect 26104 3103 26120 3137
rect 26154 3103 26170 3137
rect 26104 3069 26170 3103
rect 26104 3035 26120 3069
rect 26154 3035 26170 3069
rect 26104 3001 26170 3035
rect 26104 2967 26120 3001
rect 26154 2967 26170 3001
rect 26104 2933 26170 2967
rect 26104 2899 26120 2933
rect 26154 2899 26170 2933
rect 26104 2865 26170 2899
rect 26104 2831 26120 2865
rect 26154 2831 26170 2865
rect 26104 2797 26170 2831
rect 26104 2763 26120 2797
rect 26154 2763 26170 2797
rect 26104 2729 26170 2763
rect 26104 2695 26120 2729
rect 26154 2695 26170 2729
rect 26104 2661 26170 2695
rect 26104 2627 26120 2661
rect 26154 2627 26170 2661
rect 26104 2593 26170 2627
rect 26104 2559 26120 2593
rect 26154 2559 26170 2593
rect 26104 2518 26170 2559
rect 26200 3477 26266 3518
rect 26200 3443 26216 3477
rect 26250 3443 26266 3477
rect 26200 3409 26266 3443
rect 26200 3375 26216 3409
rect 26250 3375 26266 3409
rect 26200 3341 26266 3375
rect 26200 3307 26216 3341
rect 26250 3307 26266 3341
rect 26200 3273 26266 3307
rect 26200 3239 26216 3273
rect 26250 3239 26266 3273
rect 26200 3205 26266 3239
rect 26200 3171 26216 3205
rect 26250 3171 26266 3205
rect 26200 3137 26266 3171
rect 26200 3103 26216 3137
rect 26250 3103 26266 3137
rect 26200 3069 26266 3103
rect 26200 3035 26216 3069
rect 26250 3035 26266 3069
rect 26200 3001 26266 3035
rect 26200 2967 26216 3001
rect 26250 2967 26266 3001
rect 26200 2933 26266 2967
rect 26200 2899 26216 2933
rect 26250 2899 26266 2933
rect 26200 2865 26266 2899
rect 26200 2831 26216 2865
rect 26250 2831 26266 2865
rect 26200 2797 26266 2831
rect 26200 2763 26216 2797
rect 26250 2763 26266 2797
rect 26200 2729 26266 2763
rect 26200 2695 26216 2729
rect 26250 2695 26266 2729
rect 26200 2661 26266 2695
rect 26200 2627 26216 2661
rect 26250 2627 26266 2661
rect 26200 2593 26266 2627
rect 26200 2559 26216 2593
rect 26250 2559 26266 2593
rect 26200 2518 26266 2559
rect 26296 3477 26362 3518
rect 26296 3443 26312 3477
rect 26346 3443 26362 3477
rect 26296 3409 26362 3443
rect 26296 3375 26312 3409
rect 26346 3375 26362 3409
rect 26296 3341 26362 3375
rect 26296 3307 26312 3341
rect 26346 3307 26362 3341
rect 26296 3273 26362 3307
rect 26296 3239 26312 3273
rect 26346 3239 26362 3273
rect 26296 3205 26362 3239
rect 26296 3171 26312 3205
rect 26346 3171 26362 3205
rect 26296 3137 26362 3171
rect 26296 3103 26312 3137
rect 26346 3103 26362 3137
rect 26296 3069 26362 3103
rect 26296 3035 26312 3069
rect 26346 3035 26362 3069
rect 26296 3001 26362 3035
rect 26296 2967 26312 3001
rect 26346 2967 26362 3001
rect 26296 2933 26362 2967
rect 26296 2899 26312 2933
rect 26346 2899 26362 2933
rect 26296 2865 26362 2899
rect 26296 2831 26312 2865
rect 26346 2831 26362 2865
rect 26296 2797 26362 2831
rect 26296 2763 26312 2797
rect 26346 2763 26362 2797
rect 26296 2729 26362 2763
rect 26296 2695 26312 2729
rect 26346 2695 26362 2729
rect 26296 2661 26362 2695
rect 26296 2627 26312 2661
rect 26346 2627 26362 2661
rect 26296 2593 26362 2627
rect 26296 2559 26312 2593
rect 26346 2559 26362 2593
rect 26296 2518 26362 2559
rect 26392 3477 26458 3518
rect 26392 3443 26408 3477
rect 26442 3443 26458 3477
rect 26392 3409 26458 3443
rect 26392 3375 26408 3409
rect 26442 3375 26458 3409
rect 26392 3341 26458 3375
rect 26392 3307 26408 3341
rect 26442 3307 26458 3341
rect 26392 3273 26458 3307
rect 26392 3239 26408 3273
rect 26442 3239 26458 3273
rect 26392 3205 26458 3239
rect 26392 3171 26408 3205
rect 26442 3171 26458 3205
rect 26392 3137 26458 3171
rect 26392 3103 26408 3137
rect 26442 3103 26458 3137
rect 26392 3069 26458 3103
rect 26392 3035 26408 3069
rect 26442 3035 26458 3069
rect 26392 3001 26458 3035
rect 26392 2967 26408 3001
rect 26442 2967 26458 3001
rect 26392 2933 26458 2967
rect 26392 2899 26408 2933
rect 26442 2899 26458 2933
rect 26392 2865 26458 2899
rect 26392 2831 26408 2865
rect 26442 2831 26458 2865
rect 26392 2797 26458 2831
rect 26392 2763 26408 2797
rect 26442 2763 26458 2797
rect 26392 2729 26458 2763
rect 26392 2695 26408 2729
rect 26442 2695 26458 2729
rect 26392 2661 26458 2695
rect 26392 2627 26408 2661
rect 26442 2627 26458 2661
rect 26392 2593 26458 2627
rect 26392 2559 26408 2593
rect 26442 2559 26458 2593
rect 26392 2518 26458 2559
rect 26488 3477 26550 3518
rect 26488 3443 26504 3477
rect 26538 3443 26550 3477
rect 26488 3409 26550 3443
rect 26488 3375 26504 3409
rect 26538 3375 26550 3409
rect 26488 3341 26550 3375
rect 26488 3307 26504 3341
rect 26538 3307 26550 3341
rect 26488 3273 26550 3307
rect 26488 3239 26504 3273
rect 26538 3239 26550 3273
rect 26488 3205 26550 3239
rect 26488 3171 26504 3205
rect 26538 3171 26550 3205
rect 26488 3137 26550 3171
rect 26488 3103 26504 3137
rect 26538 3103 26550 3137
rect 26488 3069 26550 3103
rect 26488 3035 26504 3069
rect 26538 3035 26550 3069
rect 26488 3001 26550 3035
rect 26488 2967 26504 3001
rect 26538 2967 26550 3001
rect 26488 2933 26550 2967
rect 26488 2899 26504 2933
rect 26538 2899 26550 2933
rect 26488 2865 26550 2899
rect 26488 2831 26504 2865
rect 26538 2831 26550 2865
rect 26488 2797 26550 2831
rect 26488 2763 26504 2797
rect 26538 2763 26550 2797
rect 26488 2729 26550 2763
rect 26488 2695 26504 2729
rect 26538 2695 26550 2729
rect 26488 2661 26550 2695
rect 26488 2627 26504 2661
rect 26538 2627 26550 2661
rect 26488 2593 26550 2627
rect 26488 2559 26504 2593
rect 26538 2559 26550 2593
rect 26488 2518 26550 2559
rect 26720 3485 26782 3526
rect 26720 3451 26732 3485
rect 26766 3451 26782 3485
rect 26720 3417 26782 3451
rect 26720 3383 26732 3417
rect 26766 3383 26782 3417
rect 26720 3349 26782 3383
rect 26720 3315 26732 3349
rect 26766 3315 26782 3349
rect 26720 3281 26782 3315
rect 26720 3247 26732 3281
rect 26766 3247 26782 3281
rect 26720 3213 26782 3247
rect 26720 3179 26732 3213
rect 26766 3179 26782 3213
rect 26720 3145 26782 3179
rect 26720 3111 26732 3145
rect 26766 3111 26782 3145
rect 26720 3077 26782 3111
rect 26720 3043 26732 3077
rect 26766 3043 26782 3077
rect 26720 3009 26782 3043
rect 26720 2975 26732 3009
rect 26766 2975 26782 3009
rect 26720 2941 26782 2975
rect 26720 2907 26732 2941
rect 26766 2907 26782 2941
rect 26720 2873 26782 2907
rect 26720 2839 26732 2873
rect 26766 2839 26782 2873
rect 26720 2805 26782 2839
rect 26720 2771 26732 2805
rect 26766 2771 26782 2805
rect 26720 2737 26782 2771
rect 26720 2703 26732 2737
rect 26766 2703 26782 2737
rect 26720 2669 26782 2703
rect 26720 2635 26732 2669
rect 26766 2635 26782 2669
rect 26720 2601 26782 2635
rect 26720 2567 26732 2601
rect 26766 2567 26782 2601
rect 26720 2526 26782 2567
rect 26812 3485 26878 3526
rect 26812 3451 26828 3485
rect 26862 3451 26878 3485
rect 26812 3417 26878 3451
rect 26812 3383 26828 3417
rect 26862 3383 26878 3417
rect 26812 3349 26878 3383
rect 26812 3315 26828 3349
rect 26862 3315 26878 3349
rect 26812 3281 26878 3315
rect 26812 3247 26828 3281
rect 26862 3247 26878 3281
rect 26812 3213 26878 3247
rect 26812 3179 26828 3213
rect 26862 3179 26878 3213
rect 26812 3145 26878 3179
rect 26812 3111 26828 3145
rect 26862 3111 26878 3145
rect 26812 3077 26878 3111
rect 26812 3043 26828 3077
rect 26862 3043 26878 3077
rect 26812 3009 26878 3043
rect 26812 2975 26828 3009
rect 26862 2975 26878 3009
rect 26812 2941 26878 2975
rect 26812 2907 26828 2941
rect 26862 2907 26878 2941
rect 26812 2873 26878 2907
rect 26812 2839 26828 2873
rect 26862 2839 26878 2873
rect 26812 2805 26878 2839
rect 26812 2771 26828 2805
rect 26862 2771 26878 2805
rect 26812 2737 26878 2771
rect 26812 2703 26828 2737
rect 26862 2703 26878 2737
rect 26812 2669 26878 2703
rect 26812 2635 26828 2669
rect 26862 2635 26878 2669
rect 26812 2601 26878 2635
rect 26812 2567 26828 2601
rect 26862 2567 26878 2601
rect 26812 2526 26878 2567
rect 26908 3485 26974 3526
rect 26908 3451 26924 3485
rect 26958 3451 26974 3485
rect 26908 3417 26974 3451
rect 26908 3383 26924 3417
rect 26958 3383 26974 3417
rect 26908 3349 26974 3383
rect 26908 3315 26924 3349
rect 26958 3315 26974 3349
rect 26908 3281 26974 3315
rect 26908 3247 26924 3281
rect 26958 3247 26974 3281
rect 26908 3213 26974 3247
rect 26908 3179 26924 3213
rect 26958 3179 26974 3213
rect 26908 3145 26974 3179
rect 26908 3111 26924 3145
rect 26958 3111 26974 3145
rect 26908 3077 26974 3111
rect 26908 3043 26924 3077
rect 26958 3043 26974 3077
rect 26908 3009 26974 3043
rect 26908 2975 26924 3009
rect 26958 2975 26974 3009
rect 26908 2941 26974 2975
rect 26908 2907 26924 2941
rect 26958 2907 26974 2941
rect 26908 2873 26974 2907
rect 26908 2839 26924 2873
rect 26958 2839 26974 2873
rect 26908 2805 26974 2839
rect 26908 2771 26924 2805
rect 26958 2771 26974 2805
rect 26908 2737 26974 2771
rect 26908 2703 26924 2737
rect 26958 2703 26974 2737
rect 26908 2669 26974 2703
rect 26908 2635 26924 2669
rect 26958 2635 26974 2669
rect 26908 2601 26974 2635
rect 26908 2567 26924 2601
rect 26958 2567 26974 2601
rect 26908 2526 26974 2567
rect 27004 3485 27070 3526
rect 27004 3451 27020 3485
rect 27054 3451 27070 3485
rect 27004 3417 27070 3451
rect 27004 3383 27020 3417
rect 27054 3383 27070 3417
rect 27004 3349 27070 3383
rect 27004 3315 27020 3349
rect 27054 3315 27070 3349
rect 27004 3281 27070 3315
rect 27004 3247 27020 3281
rect 27054 3247 27070 3281
rect 27004 3213 27070 3247
rect 27004 3179 27020 3213
rect 27054 3179 27070 3213
rect 27004 3145 27070 3179
rect 27004 3111 27020 3145
rect 27054 3111 27070 3145
rect 27004 3077 27070 3111
rect 27004 3043 27020 3077
rect 27054 3043 27070 3077
rect 27004 3009 27070 3043
rect 27004 2975 27020 3009
rect 27054 2975 27070 3009
rect 27004 2941 27070 2975
rect 27004 2907 27020 2941
rect 27054 2907 27070 2941
rect 27004 2873 27070 2907
rect 27004 2839 27020 2873
rect 27054 2839 27070 2873
rect 27004 2805 27070 2839
rect 27004 2771 27020 2805
rect 27054 2771 27070 2805
rect 27004 2737 27070 2771
rect 27004 2703 27020 2737
rect 27054 2703 27070 2737
rect 27004 2669 27070 2703
rect 27004 2635 27020 2669
rect 27054 2635 27070 2669
rect 27004 2601 27070 2635
rect 27004 2567 27020 2601
rect 27054 2567 27070 2601
rect 27004 2526 27070 2567
rect 27100 3485 27166 3526
rect 27100 3451 27116 3485
rect 27150 3451 27166 3485
rect 27100 3417 27166 3451
rect 27100 3383 27116 3417
rect 27150 3383 27166 3417
rect 27100 3349 27166 3383
rect 27100 3315 27116 3349
rect 27150 3315 27166 3349
rect 27100 3281 27166 3315
rect 27100 3247 27116 3281
rect 27150 3247 27166 3281
rect 27100 3213 27166 3247
rect 27100 3179 27116 3213
rect 27150 3179 27166 3213
rect 27100 3145 27166 3179
rect 27100 3111 27116 3145
rect 27150 3111 27166 3145
rect 27100 3077 27166 3111
rect 27100 3043 27116 3077
rect 27150 3043 27166 3077
rect 27100 3009 27166 3043
rect 27100 2975 27116 3009
rect 27150 2975 27166 3009
rect 27100 2941 27166 2975
rect 27100 2907 27116 2941
rect 27150 2907 27166 2941
rect 27100 2873 27166 2907
rect 27100 2839 27116 2873
rect 27150 2839 27166 2873
rect 27100 2805 27166 2839
rect 27100 2771 27116 2805
rect 27150 2771 27166 2805
rect 27100 2737 27166 2771
rect 27100 2703 27116 2737
rect 27150 2703 27166 2737
rect 27100 2669 27166 2703
rect 27100 2635 27116 2669
rect 27150 2635 27166 2669
rect 27100 2601 27166 2635
rect 27100 2567 27116 2601
rect 27150 2567 27166 2601
rect 27100 2526 27166 2567
rect 27196 3485 27262 3526
rect 27196 3451 27212 3485
rect 27246 3451 27262 3485
rect 27196 3417 27262 3451
rect 27196 3383 27212 3417
rect 27246 3383 27262 3417
rect 27196 3349 27262 3383
rect 27196 3315 27212 3349
rect 27246 3315 27262 3349
rect 27196 3281 27262 3315
rect 27196 3247 27212 3281
rect 27246 3247 27262 3281
rect 27196 3213 27262 3247
rect 27196 3179 27212 3213
rect 27246 3179 27262 3213
rect 27196 3145 27262 3179
rect 27196 3111 27212 3145
rect 27246 3111 27262 3145
rect 27196 3077 27262 3111
rect 27196 3043 27212 3077
rect 27246 3043 27262 3077
rect 27196 3009 27262 3043
rect 27196 2975 27212 3009
rect 27246 2975 27262 3009
rect 27196 2941 27262 2975
rect 27196 2907 27212 2941
rect 27246 2907 27262 2941
rect 27196 2873 27262 2907
rect 27196 2839 27212 2873
rect 27246 2839 27262 2873
rect 27196 2805 27262 2839
rect 27196 2771 27212 2805
rect 27246 2771 27262 2805
rect 27196 2737 27262 2771
rect 27196 2703 27212 2737
rect 27246 2703 27262 2737
rect 27196 2669 27262 2703
rect 27196 2635 27212 2669
rect 27246 2635 27262 2669
rect 27196 2601 27262 2635
rect 27196 2567 27212 2601
rect 27246 2567 27262 2601
rect 27196 2526 27262 2567
rect 27292 3485 27358 3526
rect 27292 3451 27308 3485
rect 27342 3451 27358 3485
rect 27292 3417 27358 3451
rect 27292 3383 27308 3417
rect 27342 3383 27358 3417
rect 27292 3349 27358 3383
rect 27292 3315 27308 3349
rect 27342 3315 27358 3349
rect 27292 3281 27358 3315
rect 27292 3247 27308 3281
rect 27342 3247 27358 3281
rect 27292 3213 27358 3247
rect 27292 3179 27308 3213
rect 27342 3179 27358 3213
rect 27292 3145 27358 3179
rect 27292 3111 27308 3145
rect 27342 3111 27358 3145
rect 27292 3077 27358 3111
rect 27292 3043 27308 3077
rect 27342 3043 27358 3077
rect 27292 3009 27358 3043
rect 27292 2975 27308 3009
rect 27342 2975 27358 3009
rect 27292 2941 27358 2975
rect 27292 2907 27308 2941
rect 27342 2907 27358 2941
rect 27292 2873 27358 2907
rect 27292 2839 27308 2873
rect 27342 2839 27358 2873
rect 27292 2805 27358 2839
rect 27292 2771 27308 2805
rect 27342 2771 27358 2805
rect 27292 2737 27358 2771
rect 27292 2703 27308 2737
rect 27342 2703 27358 2737
rect 27292 2669 27358 2703
rect 27292 2635 27308 2669
rect 27342 2635 27358 2669
rect 27292 2601 27358 2635
rect 27292 2567 27308 2601
rect 27342 2567 27358 2601
rect 27292 2526 27358 2567
rect 27388 3485 27454 3526
rect 27388 3451 27404 3485
rect 27438 3451 27454 3485
rect 27388 3417 27454 3451
rect 27388 3383 27404 3417
rect 27438 3383 27454 3417
rect 27388 3349 27454 3383
rect 27388 3315 27404 3349
rect 27438 3315 27454 3349
rect 27388 3281 27454 3315
rect 27388 3247 27404 3281
rect 27438 3247 27454 3281
rect 27388 3213 27454 3247
rect 27388 3179 27404 3213
rect 27438 3179 27454 3213
rect 27388 3145 27454 3179
rect 27388 3111 27404 3145
rect 27438 3111 27454 3145
rect 27388 3077 27454 3111
rect 27388 3043 27404 3077
rect 27438 3043 27454 3077
rect 27388 3009 27454 3043
rect 27388 2975 27404 3009
rect 27438 2975 27454 3009
rect 27388 2941 27454 2975
rect 27388 2907 27404 2941
rect 27438 2907 27454 2941
rect 27388 2873 27454 2907
rect 27388 2839 27404 2873
rect 27438 2839 27454 2873
rect 27388 2805 27454 2839
rect 27388 2771 27404 2805
rect 27438 2771 27454 2805
rect 27388 2737 27454 2771
rect 27388 2703 27404 2737
rect 27438 2703 27454 2737
rect 27388 2669 27454 2703
rect 27388 2635 27404 2669
rect 27438 2635 27454 2669
rect 27388 2601 27454 2635
rect 27388 2567 27404 2601
rect 27438 2567 27454 2601
rect 27388 2526 27454 2567
rect 27484 3485 27550 3526
rect 27484 3451 27500 3485
rect 27534 3451 27550 3485
rect 27484 3417 27550 3451
rect 27484 3383 27500 3417
rect 27534 3383 27550 3417
rect 27484 3349 27550 3383
rect 27484 3315 27500 3349
rect 27534 3315 27550 3349
rect 27484 3281 27550 3315
rect 27484 3247 27500 3281
rect 27534 3247 27550 3281
rect 27484 3213 27550 3247
rect 27484 3179 27500 3213
rect 27534 3179 27550 3213
rect 27484 3145 27550 3179
rect 27484 3111 27500 3145
rect 27534 3111 27550 3145
rect 27484 3077 27550 3111
rect 27484 3043 27500 3077
rect 27534 3043 27550 3077
rect 27484 3009 27550 3043
rect 27484 2975 27500 3009
rect 27534 2975 27550 3009
rect 27484 2941 27550 2975
rect 27484 2907 27500 2941
rect 27534 2907 27550 2941
rect 27484 2873 27550 2907
rect 27484 2839 27500 2873
rect 27534 2839 27550 2873
rect 27484 2805 27550 2839
rect 27484 2771 27500 2805
rect 27534 2771 27550 2805
rect 27484 2737 27550 2771
rect 27484 2703 27500 2737
rect 27534 2703 27550 2737
rect 27484 2669 27550 2703
rect 27484 2635 27500 2669
rect 27534 2635 27550 2669
rect 27484 2601 27550 2635
rect 27484 2567 27500 2601
rect 27534 2567 27550 2601
rect 27484 2526 27550 2567
rect 27580 3485 27646 3526
rect 27580 3451 27596 3485
rect 27630 3451 27646 3485
rect 27580 3417 27646 3451
rect 27580 3383 27596 3417
rect 27630 3383 27646 3417
rect 27580 3349 27646 3383
rect 27580 3315 27596 3349
rect 27630 3315 27646 3349
rect 27580 3281 27646 3315
rect 27580 3247 27596 3281
rect 27630 3247 27646 3281
rect 27580 3213 27646 3247
rect 27580 3179 27596 3213
rect 27630 3179 27646 3213
rect 27580 3145 27646 3179
rect 27580 3111 27596 3145
rect 27630 3111 27646 3145
rect 27580 3077 27646 3111
rect 27580 3043 27596 3077
rect 27630 3043 27646 3077
rect 27580 3009 27646 3043
rect 27580 2975 27596 3009
rect 27630 2975 27646 3009
rect 27580 2941 27646 2975
rect 27580 2907 27596 2941
rect 27630 2907 27646 2941
rect 27580 2873 27646 2907
rect 27580 2839 27596 2873
rect 27630 2839 27646 2873
rect 27580 2805 27646 2839
rect 27580 2771 27596 2805
rect 27630 2771 27646 2805
rect 27580 2737 27646 2771
rect 27580 2703 27596 2737
rect 27630 2703 27646 2737
rect 27580 2669 27646 2703
rect 27580 2635 27596 2669
rect 27630 2635 27646 2669
rect 27580 2601 27646 2635
rect 27580 2567 27596 2601
rect 27630 2567 27646 2601
rect 27580 2526 27646 2567
rect 27676 3485 27742 3526
rect 27676 3451 27692 3485
rect 27726 3451 27742 3485
rect 27676 3417 27742 3451
rect 27676 3383 27692 3417
rect 27726 3383 27742 3417
rect 27676 3349 27742 3383
rect 27676 3315 27692 3349
rect 27726 3315 27742 3349
rect 27676 3281 27742 3315
rect 27676 3247 27692 3281
rect 27726 3247 27742 3281
rect 27676 3213 27742 3247
rect 27676 3179 27692 3213
rect 27726 3179 27742 3213
rect 27676 3145 27742 3179
rect 27676 3111 27692 3145
rect 27726 3111 27742 3145
rect 27676 3077 27742 3111
rect 27676 3043 27692 3077
rect 27726 3043 27742 3077
rect 27676 3009 27742 3043
rect 27676 2975 27692 3009
rect 27726 2975 27742 3009
rect 27676 2941 27742 2975
rect 27676 2907 27692 2941
rect 27726 2907 27742 2941
rect 27676 2873 27742 2907
rect 27676 2839 27692 2873
rect 27726 2839 27742 2873
rect 27676 2805 27742 2839
rect 27676 2771 27692 2805
rect 27726 2771 27742 2805
rect 27676 2737 27742 2771
rect 27676 2703 27692 2737
rect 27726 2703 27742 2737
rect 27676 2669 27742 2703
rect 27676 2635 27692 2669
rect 27726 2635 27742 2669
rect 27676 2601 27742 2635
rect 27676 2567 27692 2601
rect 27726 2567 27742 2601
rect 27676 2526 27742 2567
rect 27772 3485 27838 3526
rect 27772 3451 27788 3485
rect 27822 3451 27838 3485
rect 27772 3417 27838 3451
rect 27772 3383 27788 3417
rect 27822 3383 27838 3417
rect 27772 3349 27838 3383
rect 27772 3315 27788 3349
rect 27822 3315 27838 3349
rect 27772 3281 27838 3315
rect 27772 3247 27788 3281
rect 27822 3247 27838 3281
rect 27772 3213 27838 3247
rect 27772 3179 27788 3213
rect 27822 3179 27838 3213
rect 27772 3145 27838 3179
rect 27772 3111 27788 3145
rect 27822 3111 27838 3145
rect 27772 3077 27838 3111
rect 27772 3043 27788 3077
rect 27822 3043 27838 3077
rect 27772 3009 27838 3043
rect 27772 2975 27788 3009
rect 27822 2975 27838 3009
rect 27772 2941 27838 2975
rect 27772 2907 27788 2941
rect 27822 2907 27838 2941
rect 27772 2873 27838 2907
rect 27772 2839 27788 2873
rect 27822 2839 27838 2873
rect 27772 2805 27838 2839
rect 27772 2771 27788 2805
rect 27822 2771 27838 2805
rect 27772 2737 27838 2771
rect 27772 2703 27788 2737
rect 27822 2703 27838 2737
rect 27772 2669 27838 2703
rect 27772 2635 27788 2669
rect 27822 2635 27838 2669
rect 27772 2601 27838 2635
rect 27772 2567 27788 2601
rect 27822 2567 27838 2601
rect 27772 2526 27838 2567
rect 27868 3485 27934 3526
rect 27868 3451 27884 3485
rect 27918 3451 27934 3485
rect 27868 3417 27934 3451
rect 27868 3383 27884 3417
rect 27918 3383 27934 3417
rect 27868 3349 27934 3383
rect 27868 3315 27884 3349
rect 27918 3315 27934 3349
rect 27868 3281 27934 3315
rect 27868 3247 27884 3281
rect 27918 3247 27934 3281
rect 27868 3213 27934 3247
rect 27868 3179 27884 3213
rect 27918 3179 27934 3213
rect 27868 3145 27934 3179
rect 27868 3111 27884 3145
rect 27918 3111 27934 3145
rect 27868 3077 27934 3111
rect 27868 3043 27884 3077
rect 27918 3043 27934 3077
rect 27868 3009 27934 3043
rect 27868 2975 27884 3009
rect 27918 2975 27934 3009
rect 27868 2941 27934 2975
rect 27868 2907 27884 2941
rect 27918 2907 27934 2941
rect 27868 2873 27934 2907
rect 27868 2839 27884 2873
rect 27918 2839 27934 2873
rect 27868 2805 27934 2839
rect 27868 2771 27884 2805
rect 27918 2771 27934 2805
rect 27868 2737 27934 2771
rect 27868 2703 27884 2737
rect 27918 2703 27934 2737
rect 27868 2669 27934 2703
rect 27868 2635 27884 2669
rect 27918 2635 27934 2669
rect 27868 2601 27934 2635
rect 27868 2567 27884 2601
rect 27918 2567 27934 2601
rect 27868 2526 27934 2567
rect 27964 3485 28030 3526
rect 27964 3451 27980 3485
rect 28014 3451 28030 3485
rect 27964 3417 28030 3451
rect 27964 3383 27980 3417
rect 28014 3383 28030 3417
rect 27964 3349 28030 3383
rect 27964 3315 27980 3349
rect 28014 3315 28030 3349
rect 27964 3281 28030 3315
rect 27964 3247 27980 3281
rect 28014 3247 28030 3281
rect 27964 3213 28030 3247
rect 27964 3179 27980 3213
rect 28014 3179 28030 3213
rect 27964 3145 28030 3179
rect 27964 3111 27980 3145
rect 28014 3111 28030 3145
rect 27964 3077 28030 3111
rect 27964 3043 27980 3077
rect 28014 3043 28030 3077
rect 27964 3009 28030 3043
rect 27964 2975 27980 3009
rect 28014 2975 28030 3009
rect 27964 2941 28030 2975
rect 27964 2907 27980 2941
rect 28014 2907 28030 2941
rect 27964 2873 28030 2907
rect 27964 2839 27980 2873
rect 28014 2839 28030 2873
rect 27964 2805 28030 2839
rect 27964 2771 27980 2805
rect 28014 2771 28030 2805
rect 27964 2737 28030 2771
rect 27964 2703 27980 2737
rect 28014 2703 28030 2737
rect 27964 2669 28030 2703
rect 27964 2635 27980 2669
rect 28014 2635 28030 2669
rect 27964 2601 28030 2635
rect 27964 2567 27980 2601
rect 28014 2567 28030 2601
rect 27964 2526 28030 2567
rect 28060 3485 28126 3526
rect 28060 3451 28076 3485
rect 28110 3451 28126 3485
rect 28060 3417 28126 3451
rect 28060 3383 28076 3417
rect 28110 3383 28126 3417
rect 28060 3349 28126 3383
rect 28060 3315 28076 3349
rect 28110 3315 28126 3349
rect 28060 3281 28126 3315
rect 28060 3247 28076 3281
rect 28110 3247 28126 3281
rect 28060 3213 28126 3247
rect 28060 3179 28076 3213
rect 28110 3179 28126 3213
rect 28060 3145 28126 3179
rect 28060 3111 28076 3145
rect 28110 3111 28126 3145
rect 28060 3077 28126 3111
rect 28060 3043 28076 3077
rect 28110 3043 28126 3077
rect 28060 3009 28126 3043
rect 28060 2975 28076 3009
rect 28110 2975 28126 3009
rect 28060 2941 28126 2975
rect 28060 2907 28076 2941
rect 28110 2907 28126 2941
rect 28060 2873 28126 2907
rect 28060 2839 28076 2873
rect 28110 2839 28126 2873
rect 28060 2805 28126 2839
rect 28060 2771 28076 2805
rect 28110 2771 28126 2805
rect 28060 2737 28126 2771
rect 28060 2703 28076 2737
rect 28110 2703 28126 2737
rect 28060 2669 28126 2703
rect 28060 2635 28076 2669
rect 28110 2635 28126 2669
rect 28060 2601 28126 2635
rect 28060 2567 28076 2601
rect 28110 2567 28126 2601
rect 28060 2526 28126 2567
rect 28156 3485 28222 3526
rect 28156 3451 28172 3485
rect 28206 3451 28222 3485
rect 28156 3417 28222 3451
rect 28156 3383 28172 3417
rect 28206 3383 28222 3417
rect 28156 3349 28222 3383
rect 28156 3315 28172 3349
rect 28206 3315 28222 3349
rect 28156 3281 28222 3315
rect 28156 3247 28172 3281
rect 28206 3247 28222 3281
rect 28156 3213 28222 3247
rect 28156 3179 28172 3213
rect 28206 3179 28222 3213
rect 28156 3145 28222 3179
rect 28156 3111 28172 3145
rect 28206 3111 28222 3145
rect 28156 3077 28222 3111
rect 28156 3043 28172 3077
rect 28206 3043 28222 3077
rect 28156 3009 28222 3043
rect 28156 2975 28172 3009
rect 28206 2975 28222 3009
rect 28156 2941 28222 2975
rect 28156 2907 28172 2941
rect 28206 2907 28222 2941
rect 28156 2873 28222 2907
rect 28156 2839 28172 2873
rect 28206 2839 28222 2873
rect 28156 2805 28222 2839
rect 28156 2771 28172 2805
rect 28206 2771 28222 2805
rect 28156 2737 28222 2771
rect 28156 2703 28172 2737
rect 28206 2703 28222 2737
rect 28156 2669 28222 2703
rect 28156 2635 28172 2669
rect 28206 2635 28222 2669
rect 28156 2601 28222 2635
rect 28156 2567 28172 2601
rect 28206 2567 28222 2601
rect 28156 2526 28222 2567
rect 28252 3485 28318 3526
rect 28252 3451 28268 3485
rect 28302 3451 28318 3485
rect 28252 3417 28318 3451
rect 28252 3383 28268 3417
rect 28302 3383 28318 3417
rect 28252 3349 28318 3383
rect 28252 3315 28268 3349
rect 28302 3315 28318 3349
rect 28252 3281 28318 3315
rect 28252 3247 28268 3281
rect 28302 3247 28318 3281
rect 28252 3213 28318 3247
rect 28252 3179 28268 3213
rect 28302 3179 28318 3213
rect 28252 3145 28318 3179
rect 28252 3111 28268 3145
rect 28302 3111 28318 3145
rect 28252 3077 28318 3111
rect 28252 3043 28268 3077
rect 28302 3043 28318 3077
rect 28252 3009 28318 3043
rect 28252 2975 28268 3009
rect 28302 2975 28318 3009
rect 28252 2941 28318 2975
rect 28252 2907 28268 2941
rect 28302 2907 28318 2941
rect 28252 2873 28318 2907
rect 28252 2839 28268 2873
rect 28302 2839 28318 2873
rect 28252 2805 28318 2839
rect 28252 2771 28268 2805
rect 28302 2771 28318 2805
rect 28252 2737 28318 2771
rect 28252 2703 28268 2737
rect 28302 2703 28318 2737
rect 28252 2669 28318 2703
rect 28252 2635 28268 2669
rect 28302 2635 28318 2669
rect 28252 2601 28318 2635
rect 28252 2567 28268 2601
rect 28302 2567 28318 2601
rect 28252 2526 28318 2567
rect 28348 3485 28414 3526
rect 28348 3451 28364 3485
rect 28398 3451 28414 3485
rect 28348 3417 28414 3451
rect 28348 3383 28364 3417
rect 28398 3383 28414 3417
rect 28348 3349 28414 3383
rect 28348 3315 28364 3349
rect 28398 3315 28414 3349
rect 28348 3281 28414 3315
rect 28348 3247 28364 3281
rect 28398 3247 28414 3281
rect 28348 3213 28414 3247
rect 28348 3179 28364 3213
rect 28398 3179 28414 3213
rect 28348 3145 28414 3179
rect 28348 3111 28364 3145
rect 28398 3111 28414 3145
rect 28348 3077 28414 3111
rect 28348 3043 28364 3077
rect 28398 3043 28414 3077
rect 28348 3009 28414 3043
rect 28348 2975 28364 3009
rect 28398 2975 28414 3009
rect 28348 2941 28414 2975
rect 28348 2907 28364 2941
rect 28398 2907 28414 2941
rect 28348 2873 28414 2907
rect 28348 2839 28364 2873
rect 28398 2839 28414 2873
rect 28348 2805 28414 2839
rect 28348 2771 28364 2805
rect 28398 2771 28414 2805
rect 28348 2737 28414 2771
rect 28348 2703 28364 2737
rect 28398 2703 28414 2737
rect 28348 2669 28414 2703
rect 28348 2635 28364 2669
rect 28398 2635 28414 2669
rect 28348 2601 28414 2635
rect 28348 2567 28364 2601
rect 28398 2567 28414 2601
rect 28348 2526 28414 2567
rect 28444 3485 28510 3526
rect 28444 3451 28460 3485
rect 28494 3451 28510 3485
rect 28444 3417 28510 3451
rect 28444 3383 28460 3417
rect 28494 3383 28510 3417
rect 28444 3349 28510 3383
rect 28444 3315 28460 3349
rect 28494 3315 28510 3349
rect 28444 3281 28510 3315
rect 28444 3247 28460 3281
rect 28494 3247 28510 3281
rect 28444 3213 28510 3247
rect 28444 3179 28460 3213
rect 28494 3179 28510 3213
rect 28444 3145 28510 3179
rect 28444 3111 28460 3145
rect 28494 3111 28510 3145
rect 28444 3077 28510 3111
rect 28444 3043 28460 3077
rect 28494 3043 28510 3077
rect 28444 3009 28510 3043
rect 28444 2975 28460 3009
rect 28494 2975 28510 3009
rect 28444 2941 28510 2975
rect 28444 2907 28460 2941
rect 28494 2907 28510 2941
rect 28444 2873 28510 2907
rect 28444 2839 28460 2873
rect 28494 2839 28510 2873
rect 28444 2805 28510 2839
rect 28444 2771 28460 2805
rect 28494 2771 28510 2805
rect 28444 2737 28510 2771
rect 28444 2703 28460 2737
rect 28494 2703 28510 2737
rect 28444 2669 28510 2703
rect 28444 2635 28460 2669
rect 28494 2635 28510 2669
rect 28444 2601 28510 2635
rect 28444 2567 28460 2601
rect 28494 2567 28510 2601
rect 28444 2526 28510 2567
rect 28540 3485 28606 3526
rect 28540 3451 28556 3485
rect 28590 3451 28606 3485
rect 28540 3417 28606 3451
rect 28540 3383 28556 3417
rect 28590 3383 28606 3417
rect 28540 3349 28606 3383
rect 28540 3315 28556 3349
rect 28590 3315 28606 3349
rect 28540 3281 28606 3315
rect 28540 3247 28556 3281
rect 28590 3247 28606 3281
rect 28540 3213 28606 3247
rect 28540 3179 28556 3213
rect 28590 3179 28606 3213
rect 28540 3145 28606 3179
rect 28540 3111 28556 3145
rect 28590 3111 28606 3145
rect 28540 3077 28606 3111
rect 28540 3043 28556 3077
rect 28590 3043 28606 3077
rect 28540 3009 28606 3043
rect 28540 2975 28556 3009
rect 28590 2975 28606 3009
rect 28540 2941 28606 2975
rect 28540 2907 28556 2941
rect 28590 2907 28606 2941
rect 28540 2873 28606 2907
rect 28540 2839 28556 2873
rect 28590 2839 28606 2873
rect 28540 2805 28606 2839
rect 28540 2771 28556 2805
rect 28590 2771 28606 2805
rect 28540 2737 28606 2771
rect 28540 2703 28556 2737
rect 28590 2703 28606 2737
rect 28540 2669 28606 2703
rect 28540 2635 28556 2669
rect 28590 2635 28606 2669
rect 28540 2601 28606 2635
rect 28540 2567 28556 2601
rect 28590 2567 28606 2601
rect 28540 2526 28606 2567
rect 28636 3485 28698 3526
rect 28636 3451 28652 3485
rect 28686 3451 28698 3485
rect 28636 3417 28698 3451
rect 28636 3383 28652 3417
rect 28686 3383 28698 3417
rect 28636 3349 28698 3383
rect 28636 3315 28652 3349
rect 28686 3315 28698 3349
rect 28636 3281 28698 3315
rect 28636 3247 28652 3281
rect 28686 3247 28698 3281
rect 28636 3213 28698 3247
rect 28636 3179 28652 3213
rect 28686 3179 28698 3213
rect 28636 3145 28698 3179
rect 28636 3111 28652 3145
rect 28686 3111 28698 3145
rect 28636 3077 28698 3111
rect 28636 3043 28652 3077
rect 28686 3043 28698 3077
rect 28636 3009 28698 3043
rect 28636 2975 28652 3009
rect 28686 2975 28698 3009
rect 28636 2941 28698 2975
rect 28636 2907 28652 2941
rect 28686 2907 28698 2941
rect 28636 2873 28698 2907
rect 28636 2839 28652 2873
rect 28686 2839 28698 2873
rect 28636 2805 28698 2839
rect 28636 2771 28652 2805
rect 28686 2771 28698 2805
rect 28636 2737 28698 2771
rect 28636 2703 28652 2737
rect 28686 2703 28698 2737
rect 28636 2669 28698 2703
rect 28636 2635 28652 2669
rect 28686 2635 28698 2669
rect 28636 2601 28698 2635
rect 28636 2567 28652 2601
rect 28686 2567 28698 2601
rect 28636 2526 28698 2567
rect 14080 2439 14096 2473
rect 14130 2439 14142 2473
rect 14080 2405 14142 2439
rect 14080 2371 14096 2405
rect 14130 2371 14142 2405
rect 14080 2337 14142 2371
rect 14080 2303 14096 2337
rect 14130 2303 14142 2337
rect 14080 2269 14142 2303
rect 14080 2235 14096 2269
rect 14130 2235 14142 2269
rect 14080 2201 14142 2235
rect 14080 2167 14096 2201
rect 14130 2167 14142 2201
rect 14080 2133 14142 2167
rect 14080 2099 14096 2133
rect 14130 2099 14142 2133
rect 14080 2065 14142 2099
rect 14488 2261 14546 2276
rect 14488 2227 14500 2261
rect 14534 2227 14546 2261
rect 14488 2193 14546 2227
rect 14488 2159 14500 2193
rect 14534 2159 14546 2193
rect 14488 2125 14546 2159
rect 14488 2091 14500 2125
rect 14534 2091 14546 2125
rect 14488 2076 14546 2091
rect 14646 2261 14704 2276
rect 14646 2227 14658 2261
rect 14692 2227 14704 2261
rect 14646 2193 14704 2227
rect 14646 2159 14658 2193
rect 14692 2159 14704 2193
rect 14646 2125 14704 2159
rect 14646 2091 14658 2125
rect 14692 2091 14704 2125
rect 14646 2076 14704 2091
rect 14080 2031 14096 2065
rect 14130 2031 14142 2065
rect 14080 1997 14142 2031
rect 14080 1963 14096 1997
rect 14130 1963 14142 1997
rect 14080 1929 14142 1963
rect 14080 1895 14096 1929
rect 14130 1895 14142 1929
rect 14080 1861 14142 1895
rect 14080 1827 14096 1861
rect 14130 1827 14142 1861
rect 14080 1786 14142 1827
rect 146 1227 208 1268
rect 146 1193 158 1227
rect 192 1193 208 1227
rect 146 1159 208 1193
rect 146 1125 158 1159
rect 192 1125 208 1159
rect 146 1091 208 1125
rect -1698 1025 -1640 1066
rect -1698 991 -1686 1025
rect -1652 991 -1640 1025
rect -1698 957 -1640 991
rect -1698 923 -1686 957
rect -1652 923 -1640 957
rect -1698 889 -1640 923
rect -1698 855 -1686 889
rect -1652 855 -1640 889
rect -1698 821 -1640 855
rect -1698 787 -1686 821
rect -1652 787 -1640 821
rect -1698 753 -1640 787
rect -1698 719 -1686 753
rect -1652 719 -1640 753
rect -1698 685 -1640 719
rect -1698 651 -1686 685
rect -1652 651 -1640 685
rect -1698 617 -1640 651
rect -1698 583 -1686 617
rect -1652 583 -1640 617
rect -1698 549 -1640 583
rect -1698 515 -1686 549
rect -1652 515 -1640 549
rect -1698 481 -1640 515
rect -1698 447 -1686 481
rect -1652 447 -1640 481
rect -1698 413 -1640 447
rect -1698 379 -1686 413
rect -1652 379 -1640 413
rect -1698 345 -1640 379
rect -1698 311 -1686 345
rect -1652 311 -1640 345
rect -1698 277 -1640 311
rect -1698 243 -1686 277
rect -1652 243 -1640 277
rect -1698 209 -1640 243
rect -1698 175 -1686 209
rect -1652 175 -1640 209
rect -1698 141 -1640 175
rect -1698 107 -1686 141
rect -1652 107 -1640 141
rect -1698 66 -1640 107
rect -1600 1025 -1542 1066
rect -1600 991 -1588 1025
rect -1554 991 -1542 1025
rect -1600 957 -1542 991
rect -1600 923 -1588 957
rect -1554 923 -1542 957
rect -1600 889 -1542 923
rect -1600 855 -1588 889
rect -1554 855 -1542 889
rect -1600 821 -1542 855
rect -1600 787 -1588 821
rect -1554 787 -1542 821
rect -1600 753 -1542 787
rect -1600 719 -1588 753
rect -1554 719 -1542 753
rect -1600 685 -1542 719
rect -1600 651 -1588 685
rect -1554 651 -1542 685
rect -1600 617 -1542 651
rect -1600 583 -1588 617
rect -1554 583 -1542 617
rect -1600 549 -1542 583
rect -1600 515 -1588 549
rect -1554 515 -1542 549
rect -1600 481 -1542 515
rect -1600 447 -1588 481
rect -1554 447 -1542 481
rect -1600 413 -1542 447
rect -1600 379 -1588 413
rect -1554 379 -1542 413
rect -1600 345 -1542 379
rect -1600 311 -1588 345
rect -1554 311 -1542 345
rect -1600 277 -1542 311
rect -1600 243 -1588 277
rect -1554 243 -1542 277
rect -1600 209 -1542 243
rect -1600 175 -1588 209
rect -1554 175 -1542 209
rect -1600 141 -1542 175
rect -1600 107 -1588 141
rect -1554 107 -1542 141
rect -1600 66 -1542 107
rect -1502 1025 -1444 1066
rect -1502 991 -1490 1025
rect -1456 991 -1444 1025
rect -1502 957 -1444 991
rect -1502 923 -1490 957
rect -1456 923 -1444 957
rect -1502 889 -1444 923
rect -1502 855 -1490 889
rect -1456 855 -1444 889
rect -1502 821 -1444 855
rect -1502 787 -1490 821
rect -1456 787 -1444 821
rect -1502 753 -1444 787
rect -1502 719 -1490 753
rect -1456 719 -1444 753
rect -1502 685 -1444 719
rect -1502 651 -1490 685
rect -1456 651 -1444 685
rect -1502 617 -1444 651
rect -1502 583 -1490 617
rect -1456 583 -1444 617
rect -1502 549 -1444 583
rect -1502 515 -1490 549
rect -1456 515 -1444 549
rect -1502 481 -1444 515
rect -1502 447 -1490 481
rect -1456 447 -1444 481
rect -1502 413 -1444 447
rect -1502 379 -1490 413
rect -1456 379 -1444 413
rect -1502 345 -1444 379
rect -1502 311 -1490 345
rect -1456 311 -1444 345
rect -1502 277 -1444 311
rect -1502 243 -1490 277
rect -1456 243 -1444 277
rect -1502 209 -1444 243
rect -1502 175 -1490 209
rect -1456 175 -1444 209
rect -1502 141 -1444 175
rect -1502 107 -1490 141
rect -1456 107 -1444 141
rect -1502 66 -1444 107
rect -1404 1025 -1346 1066
rect -1404 991 -1392 1025
rect -1358 991 -1346 1025
rect -1404 957 -1346 991
rect -1404 923 -1392 957
rect -1358 923 -1346 957
rect -1404 889 -1346 923
rect -1404 855 -1392 889
rect -1358 855 -1346 889
rect -1404 821 -1346 855
rect -1404 787 -1392 821
rect -1358 787 -1346 821
rect -1404 753 -1346 787
rect -1404 719 -1392 753
rect -1358 719 -1346 753
rect -1404 685 -1346 719
rect -1404 651 -1392 685
rect -1358 651 -1346 685
rect -1404 617 -1346 651
rect -1404 583 -1392 617
rect -1358 583 -1346 617
rect -1404 549 -1346 583
rect -1404 515 -1392 549
rect -1358 515 -1346 549
rect -1404 481 -1346 515
rect -1404 447 -1392 481
rect -1358 447 -1346 481
rect -1404 413 -1346 447
rect -1404 379 -1392 413
rect -1358 379 -1346 413
rect -1404 345 -1346 379
rect -1404 311 -1392 345
rect -1358 311 -1346 345
rect -1404 277 -1346 311
rect -1404 243 -1392 277
rect -1358 243 -1346 277
rect -1404 209 -1346 243
rect -1404 175 -1392 209
rect -1358 175 -1346 209
rect -1404 141 -1346 175
rect -1404 107 -1392 141
rect -1358 107 -1346 141
rect -1404 66 -1346 107
rect -1306 1025 -1248 1066
rect -1306 991 -1294 1025
rect -1260 991 -1248 1025
rect -1306 957 -1248 991
rect -1306 923 -1294 957
rect -1260 923 -1248 957
rect -1306 889 -1248 923
rect -1306 855 -1294 889
rect -1260 855 -1248 889
rect -1306 821 -1248 855
rect -1306 787 -1294 821
rect -1260 787 -1248 821
rect -1306 753 -1248 787
rect -1306 719 -1294 753
rect -1260 719 -1248 753
rect -1306 685 -1248 719
rect -1306 651 -1294 685
rect -1260 651 -1248 685
rect -1306 617 -1248 651
rect -1306 583 -1294 617
rect -1260 583 -1248 617
rect -1306 549 -1248 583
rect -1306 515 -1294 549
rect -1260 515 -1248 549
rect -1306 481 -1248 515
rect -1306 447 -1294 481
rect -1260 447 -1248 481
rect -1306 413 -1248 447
rect -1306 379 -1294 413
rect -1260 379 -1248 413
rect -1306 345 -1248 379
rect -1306 311 -1294 345
rect -1260 311 -1248 345
rect -1306 277 -1248 311
rect -1306 243 -1294 277
rect -1260 243 -1248 277
rect -1306 209 -1248 243
rect -1306 175 -1294 209
rect -1260 175 -1248 209
rect -1306 141 -1248 175
rect -1306 107 -1294 141
rect -1260 107 -1248 141
rect -1306 66 -1248 107
rect -1208 1025 -1150 1066
rect -1208 991 -1196 1025
rect -1162 991 -1150 1025
rect -1208 957 -1150 991
rect -1208 923 -1196 957
rect -1162 923 -1150 957
rect -1208 889 -1150 923
rect -1208 855 -1196 889
rect -1162 855 -1150 889
rect -1208 821 -1150 855
rect -1208 787 -1196 821
rect -1162 787 -1150 821
rect -1208 753 -1150 787
rect -1208 719 -1196 753
rect -1162 719 -1150 753
rect -1208 685 -1150 719
rect -1208 651 -1196 685
rect -1162 651 -1150 685
rect -1208 617 -1150 651
rect -1208 583 -1196 617
rect -1162 583 -1150 617
rect -1208 549 -1150 583
rect -1208 515 -1196 549
rect -1162 515 -1150 549
rect -1208 481 -1150 515
rect -1208 447 -1196 481
rect -1162 447 -1150 481
rect -1208 413 -1150 447
rect -1208 379 -1196 413
rect -1162 379 -1150 413
rect -1208 345 -1150 379
rect -1208 311 -1196 345
rect -1162 311 -1150 345
rect -1208 277 -1150 311
rect -1208 243 -1196 277
rect -1162 243 -1150 277
rect -1208 209 -1150 243
rect -1208 175 -1196 209
rect -1162 175 -1150 209
rect -1208 141 -1150 175
rect -1208 107 -1196 141
rect -1162 107 -1150 141
rect -1208 66 -1150 107
rect -1110 1025 -1052 1066
rect -1110 991 -1098 1025
rect -1064 991 -1052 1025
rect -1110 957 -1052 991
rect -1110 923 -1098 957
rect -1064 923 -1052 957
rect -1110 889 -1052 923
rect -1110 855 -1098 889
rect -1064 855 -1052 889
rect -1110 821 -1052 855
rect -1110 787 -1098 821
rect -1064 787 -1052 821
rect -1110 753 -1052 787
rect -1110 719 -1098 753
rect -1064 719 -1052 753
rect -1110 685 -1052 719
rect -1110 651 -1098 685
rect -1064 651 -1052 685
rect -1110 617 -1052 651
rect -1110 583 -1098 617
rect -1064 583 -1052 617
rect -1110 549 -1052 583
rect -1110 515 -1098 549
rect -1064 515 -1052 549
rect -1110 481 -1052 515
rect -1110 447 -1098 481
rect -1064 447 -1052 481
rect -1110 413 -1052 447
rect -1110 379 -1098 413
rect -1064 379 -1052 413
rect -1110 345 -1052 379
rect -1110 311 -1098 345
rect -1064 311 -1052 345
rect -1110 277 -1052 311
rect -1110 243 -1098 277
rect -1064 243 -1052 277
rect -1110 209 -1052 243
rect -1110 175 -1098 209
rect -1064 175 -1052 209
rect -1110 141 -1052 175
rect -1110 107 -1098 141
rect -1064 107 -1052 141
rect -1110 66 -1052 107
rect -1012 1025 -954 1066
rect -1012 991 -1000 1025
rect -966 991 -954 1025
rect -1012 957 -954 991
rect -1012 923 -1000 957
rect -966 923 -954 957
rect -1012 889 -954 923
rect -1012 855 -1000 889
rect -966 855 -954 889
rect -1012 821 -954 855
rect -1012 787 -1000 821
rect -966 787 -954 821
rect -1012 753 -954 787
rect -1012 719 -1000 753
rect -966 719 -954 753
rect -1012 685 -954 719
rect -1012 651 -1000 685
rect -966 651 -954 685
rect -1012 617 -954 651
rect -1012 583 -1000 617
rect -966 583 -954 617
rect -1012 549 -954 583
rect -1012 515 -1000 549
rect -966 515 -954 549
rect -1012 481 -954 515
rect -1012 447 -1000 481
rect -966 447 -954 481
rect -1012 413 -954 447
rect -1012 379 -1000 413
rect -966 379 -954 413
rect -1012 345 -954 379
rect -1012 311 -1000 345
rect -966 311 -954 345
rect -1012 277 -954 311
rect -1012 243 -1000 277
rect -966 243 -954 277
rect -1012 209 -954 243
rect -1012 175 -1000 209
rect -966 175 -954 209
rect -1012 141 -954 175
rect -1012 107 -1000 141
rect -966 107 -954 141
rect -1012 66 -954 107
rect -914 1025 -856 1066
rect -914 991 -902 1025
rect -868 991 -856 1025
rect -914 957 -856 991
rect -914 923 -902 957
rect -868 923 -856 957
rect -914 889 -856 923
rect -914 855 -902 889
rect -868 855 -856 889
rect -914 821 -856 855
rect -914 787 -902 821
rect -868 787 -856 821
rect -914 753 -856 787
rect -914 719 -902 753
rect -868 719 -856 753
rect -914 685 -856 719
rect -914 651 -902 685
rect -868 651 -856 685
rect -914 617 -856 651
rect -914 583 -902 617
rect -868 583 -856 617
rect -914 549 -856 583
rect -914 515 -902 549
rect -868 515 -856 549
rect -914 481 -856 515
rect -914 447 -902 481
rect -868 447 -856 481
rect -914 413 -856 447
rect -914 379 -902 413
rect -868 379 -856 413
rect -914 345 -856 379
rect -914 311 -902 345
rect -868 311 -856 345
rect -914 277 -856 311
rect -914 243 -902 277
rect -868 243 -856 277
rect 146 1057 158 1091
rect 192 1057 208 1091
rect 146 1023 208 1057
rect 146 989 158 1023
rect 192 989 208 1023
rect 146 955 208 989
rect 146 921 158 955
rect 192 921 208 955
rect 146 887 208 921
rect 146 853 158 887
rect 192 853 208 887
rect 146 819 208 853
rect 146 785 158 819
rect 192 785 208 819
rect 146 751 208 785
rect 146 717 158 751
rect 192 717 208 751
rect 146 683 208 717
rect 146 649 158 683
rect 192 649 208 683
rect 146 615 208 649
rect 146 581 158 615
rect 192 581 208 615
rect 146 547 208 581
rect 146 513 158 547
rect 192 513 208 547
rect 146 479 208 513
rect 146 445 158 479
rect 192 445 208 479
rect 146 411 208 445
rect 146 377 158 411
rect 192 377 208 411
rect 146 343 208 377
rect 146 309 158 343
rect 192 309 208 343
rect 146 268 208 309
rect 238 1227 304 1268
rect 238 1193 254 1227
rect 288 1193 304 1227
rect 238 1159 304 1193
rect 238 1125 254 1159
rect 288 1125 304 1159
rect 238 1091 304 1125
rect 238 1057 254 1091
rect 288 1057 304 1091
rect 238 1023 304 1057
rect 238 989 254 1023
rect 288 989 304 1023
rect 238 955 304 989
rect 238 921 254 955
rect 288 921 304 955
rect 238 887 304 921
rect 238 853 254 887
rect 288 853 304 887
rect 238 819 304 853
rect 238 785 254 819
rect 288 785 304 819
rect 238 751 304 785
rect 238 717 254 751
rect 288 717 304 751
rect 238 683 304 717
rect 238 649 254 683
rect 288 649 304 683
rect 238 615 304 649
rect 238 581 254 615
rect 288 581 304 615
rect 238 547 304 581
rect 238 513 254 547
rect 288 513 304 547
rect 238 479 304 513
rect 238 445 254 479
rect 288 445 304 479
rect 238 411 304 445
rect 238 377 254 411
rect 288 377 304 411
rect 238 343 304 377
rect 238 309 254 343
rect 288 309 304 343
rect 238 268 304 309
rect 334 1227 400 1268
rect 334 1193 350 1227
rect 384 1193 400 1227
rect 334 1159 400 1193
rect 334 1125 350 1159
rect 384 1125 400 1159
rect 334 1091 400 1125
rect 334 1057 350 1091
rect 384 1057 400 1091
rect 334 1023 400 1057
rect 334 989 350 1023
rect 384 989 400 1023
rect 334 955 400 989
rect 334 921 350 955
rect 384 921 400 955
rect 334 887 400 921
rect 334 853 350 887
rect 384 853 400 887
rect 334 819 400 853
rect 334 785 350 819
rect 384 785 400 819
rect 334 751 400 785
rect 334 717 350 751
rect 384 717 400 751
rect 334 683 400 717
rect 334 649 350 683
rect 384 649 400 683
rect 334 615 400 649
rect 334 581 350 615
rect 384 581 400 615
rect 334 547 400 581
rect 334 513 350 547
rect 384 513 400 547
rect 334 479 400 513
rect 334 445 350 479
rect 384 445 400 479
rect 334 411 400 445
rect 334 377 350 411
rect 384 377 400 411
rect 334 343 400 377
rect 334 309 350 343
rect 384 309 400 343
rect 334 268 400 309
rect 430 1227 496 1268
rect 430 1193 446 1227
rect 480 1193 496 1227
rect 430 1159 496 1193
rect 430 1125 446 1159
rect 480 1125 496 1159
rect 430 1091 496 1125
rect 430 1057 446 1091
rect 480 1057 496 1091
rect 430 1023 496 1057
rect 430 989 446 1023
rect 480 989 496 1023
rect 430 955 496 989
rect 430 921 446 955
rect 480 921 496 955
rect 430 887 496 921
rect 430 853 446 887
rect 480 853 496 887
rect 430 819 496 853
rect 430 785 446 819
rect 480 785 496 819
rect 430 751 496 785
rect 430 717 446 751
rect 480 717 496 751
rect 430 683 496 717
rect 430 649 446 683
rect 480 649 496 683
rect 430 615 496 649
rect 430 581 446 615
rect 480 581 496 615
rect 430 547 496 581
rect 430 513 446 547
rect 480 513 496 547
rect 430 479 496 513
rect 430 445 446 479
rect 480 445 496 479
rect 430 411 496 445
rect 430 377 446 411
rect 480 377 496 411
rect 430 343 496 377
rect 430 309 446 343
rect 480 309 496 343
rect 430 268 496 309
rect 526 1227 592 1268
rect 526 1193 542 1227
rect 576 1193 592 1227
rect 526 1159 592 1193
rect 526 1125 542 1159
rect 576 1125 592 1159
rect 526 1091 592 1125
rect 526 1057 542 1091
rect 576 1057 592 1091
rect 526 1023 592 1057
rect 526 989 542 1023
rect 576 989 592 1023
rect 526 955 592 989
rect 526 921 542 955
rect 576 921 592 955
rect 526 887 592 921
rect 526 853 542 887
rect 576 853 592 887
rect 526 819 592 853
rect 526 785 542 819
rect 576 785 592 819
rect 526 751 592 785
rect 526 717 542 751
rect 576 717 592 751
rect 526 683 592 717
rect 526 649 542 683
rect 576 649 592 683
rect 526 615 592 649
rect 526 581 542 615
rect 576 581 592 615
rect 526 547 592 581
rect 526 513 542 547
rect 576 513 592 547
rect 526 479 592 513
rect 526 445 542 479
rect 576 445 592 479
rect 526 411 592 445
rect 526 377 542 411
rect 576 377 592 411
rect 526 343 592 377
rect 526 309 542 343
rect 576 309 592 343
rect 526 268 592 309
rect 622 1227 688 1268
rect 622 1193 638 1227
rect 672 1193 688 1227
rect 622 1159 688 1193
rect 622 1125 638 1159
rect 672 1125 688 1159
rect 622 1091 688 1125
rect 622 1057 638 1091
rect 672 1057 688 1091
rect 622 1023 688 1057
rect 622 989 638 1023
rect 672 989 688 1023
rect 622 955 688 989
rect 622 921 638 955
rect 672 921 688 955
rect 622 887 688 921
rect 622 853 638 887
rect 672 853 688 887
rect 622 819 688 853
rect 622 785 638 819
rect 672 785 688 819
rect 622 751 688 785
rect 622 717 638 751
rect 672 717 688 751
rect 622 683 688 717
rect 622 649 638 683
rect 672 649 688 683
rect 622 615 688 649
rect 622 581 638 615
rect 672 581 688 615
rect 622 547 688 581
rect 622 513 638 547
rect 672 513 688 547
rect 622 479 688 513
rect 622 445 638 479
rect 672 445 688 479
rect 622 411 688 445
rect 622 377 638 411
rect 672 377 688 411
rect 622 343 688 377
rect 622 309 638 343
rect 672 309 688 343
rect 622 268 688 309
rect 718 1227 784 1268
rect 718 1193 734 1227
rect 768 1193 784 1227
rect 718 1159 784 1193
rect 718 1125 734 1159
rect 768 1125 784 1159
rect 718 1091 784 1125
rect 718 1057 734 1091
rect 768 1057 784 1091
rect 718 1023 784 1057
rect 718 989 734 1023
rect 768 989 784 1023
rect 718 955 784 989
rect 718 921 734 955
rect 768 921 784 955
rect 718 887 784 921
rect 718 853 734 887
rect 768 853 784 887
rect 718 819 784 853
rect 718 785 734 819
rect 768 785 784 819
rect 718 751 784 785
rect 718 717 734 751
rect 768 717 784 751
rect 718 683 784 717
rect 718 649 734 683
rect 768 649 784 683
rect 718 615 784 649
rect 718 581 734 615
rect 768 581 784 615
rect 718 547 784 581
rect 718 513 734 547
rect 768 513 784 547
rect 718 479 784 513
rect 718 445 734 479
rect 768 445 784 479
rect 718 411 784 445
rect 718 377 734 411
rect 768 377 784 411
rect 718 343 784 377
rect 718 309 734 343
rect 768 309 784 343
rect 718 268 784 309
rect 814 1227 880 1268
rect 814 1193 830 1227
rect 864 1193 880 1227
rect 814 1159 880 1193
rect 814 1125 830 1159
rect 864 1125 880 1159
rect 814 1091 880 1125
rect 814 1057 830 1091
rect 864 1057 880 1091
rect 814 1023 880 1057
rect 814 989 830 1023
rect 864 989 880 1023
rect 814 955 880 989
rect 814 921 830 955
rect 864 921 880 955
rect 814 887 880 921
rect 814 853 830 887
rect 864 853 880 887
rect 814 819 880 853
rect 814 785 830 819
rect 864 785 880 819
rect 814 751 880 785
rect 814 717 830 751
rect 864 717 880 751
rect 814 683 880 717
rect 814 649 830 683
rect 864 649 880 683
rect 814 615 880 649
rect 814 581 830 615
rect 864 581 880 615
rect 814 547 880 581
rect 814 513 830 547
rect 864 513 880 547
rect 814 479 880 513
rect 814 445 830 479
rect 864 445 880 479
rect 814 411 880 445
rect 814 377 830 411
rect 864 377 880 411
rect 814 343 880 377
rect 814 309 830 343
rect 864 309 880 343
rect 814 268 880 309
rect 910 1227 976 1268
rect 910 1193 926 1227
rect 960 1193 976 1227
rect 910 1159 976 1193
rect 910 1125 926 1159
rect 960 1125 976 1159
rect 910 1091 976 1125
rect 910 1057 926 1091
rect 960 1057 976 1091
rect 910 1023 976 1057
rect 910 989 926 1023
rect 960 989 976 1023
rect 910 955 976 989
rect 910 921 926 955
rect 960 921 976 955
rect 910 887 976 921
rect 910 853 926 887
rect 960 853 976 887
rect 910 819 976 853
rect 910 785 926 819
rect 960 785 976 819
rect 910 751 976 785
rect 910 717 926 751
rect 960 717 976 751
rect 910 683 976 717
rect 910 649 926 683
rect 960 649 976 683
rect 910 615 976 649
rect 910 581 926 615
rect 960 581 976 615
rect 910 547 976 581
rect 910 513 926 547
rect 960 513 976 547
rect 910 479 976 513
rect 910 445 926 479
rect 960 445 976 479
rect 910 411 976 445
rect 910 377 926 411
rect 960 377 976 411
rect 910 343 976 377
rect 910 309 926 343
rect 960 309 976 343
rect 910 268 976 309
rect 1006 1227 1072 1268
rect 1006 1193 1022 1227
rect 1056 1193 1072 1227
rect 1006 1159 1072 1193
rect 1006 1125 1022 1159
rect 1056 1125 1072 1159
rect 1006 1091 1072 1125
rect 1006 1057 1022 1091
rect 1056 1057 1072 1091
rect 1006 1023 1072 1057
rect 1006 989 1022 1023
rect 1056 989 1072 1023
rect 1006 955 1072 989
rect 1006 921 1022 955
rect 1056 921 1072 955
rect 1006 887 1072 921
rect 1006 853 1022 887
rect 1056 853 1072 887
rect 1006 819 1072 853
rect 1006 785 1022 819
rect 1056 785 1072 819
rect 1006 751 1072 785
rect 1006 717 1022 751
rect 1056 717 1072 751
rect 1006 683 1072 717
rect 1006 649 1022 683
rect 1056 649 1072 683
rect 1006 615 1072 649
rect 1006 581 1022 615
rect 1056 581 1072 615
rect 1006 547 1072 581
rect 1006 513 1022 547
rect 1056 513 1072 547
rect 1006 479 1072 513
rect 1006 445 1022 479
rect 1056 445 1072 479
rect 1006 411 1072 445
rect 1006 377 1022 411
rect 1056 377 1072 411
rect 1006 343 1072 377
rect 1006 309 1022 343
rect 1056 309 1072 343
rect 1006 268 1072 309
rect 1102 1227 1168 1268
rect 1102 1193 1118 1227
rect 1152 1193 1168 1227
rect 1102 1159 1168 1193
rect 1102 1125 1118 1159
rect 1152 1125 1168 1159
rect 1102 1091 1168 1125
rect 1102 1057 1118 1091
rect 1152 1057 1168 1091
rect 1102 1023 1168 1057
rect 1102 989 1118 1023
rect 1152 989 1168 1023
rect 1102 955 1168 989
rect 1102 921 1118 955
rect 1152 921 1168 955
rect 1102 887 1168 921
rect 1102 853 1118 887
rect 1152 853 1168 887
rect 1102 819 1168 853
rect 1102 785 1118 819
rect 1152 785 1168 819
rect 1102 751 1168 785
rect 1102 717 1118 751
rect 1152 717 1168 751
rect 1102 683 1168 717
rect 1102 649 1118 683
rect 1152 649 1168 683
rect 1102 615 1168 649
rect 1102 581 1118 615
rect 1152 581 1168 615
rect 1102 547 1168 581
rect 1102 513 1118 547
rect 1152 513 1168 547
rect 1102 479 1168 513
rect 1102 445 1118 479
rect 1152 445 1168 479
rect 1102 411 1168 445
rect 1102 377 1118 411
rect 1152 377 1168 411
rect 1102 343 1168 377
rect 1102 309 1118 343
rect 1152 309 1168 343
rect 1102 268 1168 309
rect 1198 1227 1264 1268
rect 1198 1193 1214 1227
rect 1248 1193 1264 1227
rect 1198 1159 1264 1193
rect 1198 1125 1214 1159
rect 1248 1125 1264 1159
rect 1198 1091 1264 1125
rect 1198 1057 1214 1091
rect 1248 1057 1264 1091
rect 1198 1023 1264 1057
rect 1198 989 1214 1023
rect 1248 989 1264 1023
rect 1198 955 1264 989
rect 1198 921 1214 955
rect 1248 921 1264 955
rect 1198 887 1264 921
rect 1198 853 1214 887
rect 1248 853 1264 887
rect 1198 819 1264 853
rect 1198 785 1214 819
rect 1248 785 1264 819
rect 1198 751 1264 785
rect 1198 717 1214 751
rect 1248 717 1264 751
rect 1198 683 1264 717
rect 1198 649 1214 683
rect 1248 649 1264 683
rect 1198 615 1264 649
rect 1198 581 1214 615
rect 1248 581 1264 615
rect 1198 547 1264 581
rect 1198 513 1214 547
rect 1248 513 1264 547
rect 1198 479 1264 513
rect 1198 445 1214 479
rect 1248 445 1264 479
rect 1198 411 1264 445
rect 1198 377 1214 411
rect 1248 377 1264 411
rect 1198 343 1264 377
rect 1198 309 1214 343
rect 1248 309 1264 343
rect 1198 268 1264 309
rect 1294 1227 1356 1268
rect 1294 1193 1310 1227
rect 1344 1193 1356 1227
rect 1294 1159 1356 1193
rect 1294 1125 1310 1159
rect 1344 1125 1356 1159
rect 1294 1091 1356 1125
rect 1294 1057 1310 1091
rect 1344 1057 1356 1091
rect 1294 1023 1356 1057
rect 1294 989 1310 1023
rect 1344 989 1356 1023
rect 1294 955 1356 989
rect 1294 921 1310 955
rect 1344 921 1356 955
rect 1294 887 1356 921
rect 1294 853 1310 887
rect 1344 853 1356 887
rect 1294 819 1356 853
rect 1294 785 1310 819
rect 1344 785 1356 819
rect 1294 751 1356 785
rect 1294 717 1310 751
rect 1344 717 1356 751
rect 1294 683 1356 717
rect 1294 649 1310 683
rect 1344 649 1356 683
rect 1294 615 1356 649
rect 1294 581 1310 615
rect 1344 581 1356 615
rect 1294 547 1356 581
rect 1294 513 1310 547
rect 1344 513 1356 547
rect 1294 479 1356 513
rect 1294 445 1310 479
rect 1344 445 1356 479
rect 1294 411 1356 445
rect 1294 377 1310 411
rect 1344 377 1356 411
rect 1294 343 1356 377
rect 1294 309 1310 343
rect 1344 309 1356 343
rect 1294 268 1356 309
rect 1914 1227 1976 1268
rect 1914 1193 1926 1227
rect 1960 1193 1976 1227
rect 1914 1159 1976 1193
rect 1914 1125 1926 1159
rect 1960 1125 1976 1159
rect 1914 1091 1976 1125
rect 1914 1057 1926 1091
rect 1960 1057 1976 1091
rect 1914 1023 1976 1057
rect 1914 989 1926 1023
rect 1960 989 1976 1023
rect 1914 955 1976 989
rect 1914 921 1926 955
rect 1960 921 1976 955
rect 1914 887 1976 921
rect 1914 853 1926 887
rect 1960 853 1976 887
rect 1914 819 1976 853
rect 1914 785 1926 819
rect 1960 785 1976 819
rect 1914 751 1976 785
rect 1914 717 1926 751
rect 1960 717 1976 751
rect 1914 683 1976 717
rect 1914 649 1926 683
rect 1960 649 1976 683
rect 1914 615 1976 649
rect 1914 581 1926 615
rect 1960 581 1976 615
rect 1914 547 1976 581
rect 1914 513 1926 547
rect 1960 513 1976 547
rect 1914 479 1976 513
rect 1914 445 1926 479
rect 1960 445 1976 479
rect 1914 411 1976 445
rect 1914 377 1926 411
rect 1960 377 1976 411
rect 1914 343 1976 377
rect 1914 309 1926 343
rect 1960 309 1976 343
rect 1914 268 1976 309
rect 2006 1227 2072 1268
rect 2006 1193 2022 1227
rect 2056 1193 2072 1227
rect 2006 1159 2072 1193
rect 2006 1125 2022 1159
rect 2056 1125 2072 1159
rect 2006 1091 2072 1125
rect 2006 1057 2022 1091
rect 2056 1057 2072 1091
rect 2006 1023 2072 1057
rect 2006 989 2022 1023
rect 2056 989 2072 1023
rect 2006 955 2072 989
rect 2006 921 2022 955
rect 2056 921 2072 955
rect 2006 887 2072 921
rect 2006 853 2022 887
rect 2056 853 2072 887
rect 2006 819 2072 853
rect 2006 785 2022 819
rect 2056 785 2072 819
rect 2006 751 2072 785
rect 2006 717 2022 751
rect 2056 717 2072 751
rect 2006 683 2072 717
rect 2006 649 2022 683
rect 2056 649 2072 683
rect 2006 615 2072 649
rect 2006 581 2022 615
rect 2056 581 2072 615
rect 2006 547 2072 581
rect 2006 513 2022 547
rect 2056 513 2072 547
rect 2006 479 2072 513
rect 2006 445 2022 479
rect 2056 445 2072 479
rect 2006 411 2072 445
rect 2006 377 2022 411
rect 2056 377 2072 411
rect 2006 343 2072 377
rect 2006 309 2022 343
rect 2056 309 2072 343
rect 2006 268 2072 309
rect 2102 1227 2168 1268
rect 2102 1193 2118 1227
rect 2152 1193 2168 1227
rect 2102 1159 2168 1193
rect 2102 1125 2118 1159
rect 2152 1125 2168 1159
rect 2102 1091 2168 1125
rect 2102 1057 2118 1091
rect 2152 1057 2168 1091
rect 2102 1023 2168 1057
rect 2102 989 2118 1023
rect 2152 989 2168 1023
rect 2102 955 2168 989
rect 2102 921 2118 955
rect 2152 921 2168 955
rect 2102 887 2168 921
rect 2102 853 2118 887
rect 2152 853 2168 887
rect 2102 819 2168 853
rect 2102 785 2118 819
rect 2152 785 2168 819
rect 2102 751 2168 785
rect 2102 717 2118 751
rect 2152 717 2168 751
rect 2102 683 2168 717
rect 2102 649 2118 683
rect 2152 649 2168 683
rect 2102 615 2168 649
rect 2102 581 2118 615
rect 2152 581 2168 615
rect 2102 547 2168 581
rect 2102 513 2118 547
rect 2152 513 2168 547
rect 2102 479 2168 513
rect 2102 445 2118 479
rect 2152 445 2168 479
rect 2102 411 2168 445
rect 2102 377 2118 411
rect 2152 377 2168 411
rect 2102 343 2168 377
rect 2102 309 2118 343
rect 2152 309 2168 343
rect 2102 268 2168 309
rect 2198 1227 2264 1268
rect 2198 1193 2214 1227
rect 2248 1193 2264 1227
rect 2198 1159 2264 1193
rect 2198 1125 2214 1159
rect 2248 1125 2264 1159
rect 2198 1091 2264 1125
rect 2198 1057 2214 1091
rect 2248 1057 2264 1091
rect 2198 1023 2264 1057
rect 2198 989 2214 1023
rect 2248 989 2264 1023
rect 2198 955 2264 989
rect 2198 921 2214 955
rect 2248 921 2264 955
rect 2198 887 2264 921
rect 2198 853 2214 887
rect 2248 853 2264 887
rect 2198 819 2264 853
rect 2198 785 2214 819
rect 2248 785 2264 819
rect 2198 751 2264 785
rect 2198 717 2214 751
rect 2248 717 2264 751
rect 2198 683 2264 717
rect 2198 649 2214 683
rect 2248 649 2264 683
rect 2198 615 2264 649
rect 2198 581 2214 615
rect 2248 581 2264 615
rect 2198 547 2264 581
rect 2198 513 2214 547
rect 2248 513 2264 547
rect 2198 479 2264 513
rect 2198 445 2214 479
rect 2248 445 2264 479
rect 2198 411 2264 445
rect 2198 377 2214 411
rect 2248 377 2264 411
rect 2198 343 2264 377
rect 2198 309 2214 343
rect 2248 309 2264 343
rect 2198 268 2264 309
rect 2294 1227 2360 1268
rect 2294 1193 2310 1227
rect 2344 1193 2360 1227
rect 2294 1159 2360 1193
rect 2294 1125 2310 1159
rect 2344 1125 2360 1159
rect 2294 1091 2360 1125
rect 2294 1057 2310 1091
rect 2344 1057 2360 1091
rect 2294 1023 2360 1057
rect 2294 989 2310 1023
rect 2344 989 2360 1023
rect 2294 955 2360 989
rect 2294 921 2310 955
rect 2344 921 2360 955
rect 2294 887 2360 921
rect 2294 853 2310 887
rect 2344 853 2360 887
rect 2294 819 2360 853
rect 2294 785 2310 819
rect 2344 785 2360 819
rect 2294 751 2360 785
rect 2294 717 2310 751
rect 2344 717 2360 751
rect 2294 683 2360 717
rect 2294 649 2310 683
rect 2344 649 2360 683
rect 2294 615 2360 649
rect 2294 581 2310 615
rect 2344 581 2360 615
rect 2294 547 2360 581
rect 2294 513 2310 547
rect 2344 513 2360 547
rect 2294 479 2360 513
rect 2294 445 2310 479
rect 2344 445 2360 479
rect 2294 411 2360 445
rect 2294 377 2310 411
rect 2344 377 2360 411
rect 2294 343 2360 377
rect 2294 309 2310 343
rect 2344 309 2360 343
rect 2294 268 2360 309
rect 2390 1227 2456 1268
rect 2390 1193 2406 1227
rect 2440 1193 2456 1227
rect 2390 1159 2456 1193
rect 2390 1125 2406 1159
rect 2440 1125 2456 1159
rect 2390 1091 2456 1125
rect 2390 1057 2406 1091
rect 2440 1057 2456 1091
rect 2390 1023 2456 1057
rect 2390 989 2406 1023
rect 2440 989 2456 1023
rect 2390 955 2456 989
rect 2390 921 2406 955
rect 2440 921 2456 955
rect 2390 887 2456 921
rect 2390 853 2406 887
rect 2440 853 2456 887
rect 2390 819 2456 853
rect 2390 785 2406 819
rect 2440 785 2456 819
rect 2390 751 2456 785
rect 2390 717 2406 751
rect 2440 717 2456 751
rect 2390 683 2456 717
rect 2390 649 2406 683
rect 2440 649 2456 683
rect 2390 615 2456 649
rect 2390 581 2406 615
rect 2440 581 2456 615
rect 2390 547 2456 581
rect 2390 513 2406 547
rect 2440 513 2456 547
rect 2390 479 2456 513
rect 2390 445 2406 479
rect 2440 445 2456 479
rect 2390 411 2456 445
rect 2390 377 2406 411
rect 2440 377 2456 411
rect 2390 343 2456 377
rect 2390 309 2406 343
rect 2440 309 2456 343
rect 2390 268 2456 309
rect 2486 1227 2552 1268
rect 2486 1193 2502 1227
rect 2536 1193 2552 1227
rect 2486 1159 2552 1193
rect 2486 1125 2502 1159
rect 2536 1125 2552 1159
rect 2486 1091 2552 1125
rect 2486 1057 2502 1091
rect 2536 1057 2552 1091
rect 2486 1023 2552 1057
rect 2486 989 2502 1023
rect 2536 989 2552 1023
rect 2486 955 2552 989
rect 2486 921 2502 955
rect 2536 921 2552 955
rect 2486 887 2552 921
rect 2486 853 2502 887
rect 2536 853 2552 887
rect 2486 819 2552 853
rect 2486 785 2502 819
rect 2536 785 2552 819
rect 2486 751 2552 785
rect 2486 717 2502 751
rect 2536 717 2552 751
rect 2486 683 2552 717
rect 2486 649 2502 683
rect 2536 649 2552 683
rect 2486 615 2552 649
rect 2486 581 2502 615
rect 2536 581 2552 615
rect 2486 547 2552 581
rect 2486 513 2502 547
rect 2536 513 2552 547
rect 2486 479 2552 513
rect 2486 445 2502 479
rect 2536 445 2552 479
rect 2486 411 2552 445
rect 2486 377 2502 411
rect 2536 377 2552 411
rect 2486 343 2552 377
rect 2486 309 2502 343
rect 2536 309 2552 343
rect 2486 268 2552 309
rect 2582 1227 2648 1268
rect 2582 1193 2598 1227
rect 2632 1193 2648 1227
rect 2582 1159 2648 1193
rect 2582 1125 2598 1159
rect 2632 1125 2648 1159
rect 2582 1091 2648 1125
rect 2582 1057 2598 1091
rect 2632 1057 2648 1091
rect 2582 1023 2648 1057
rect 2582 989 2598 1023
rect 2632 989 2648 1023
rect 2582 955 2648 989
rect 2582 921 2598 955
rect 2632 921 2648 955
rect 2582 887 2648 921
rect 2582 853 2598 887
rect 2632 853 2648 887
rect 2582 819 2648 853
rect 2582 785 2598 819
rect 2632 785 2648 819
rect 2582 751 2648 785
rect 2582 717 2598 751
rect 2632 717 2648 751
rect 2582 683 2648 717
rect 2582 649 2598 683
rect 2632 649 2648 683
rect 2582 615 2648 649
rect 2582 581 2598 615
rect 2632 581 2648 615
rect 2582 547 2648 581
rect 2582 513 2598 547
rect 2632 513 2648 547
rect 2582 479 2648 513
rect 2582 445 2598 479
rect 2632 445 2648 479
rect 2582 411 2648 445
rect 2582 377 2598 411
rect 2632 377 2648 411
rect 2582 343 2648 377
rect 2582 309 2598 343
rect 2632 309 2648 343
rect 2582 268 2648 309
rect 2678 1227 2744 1268
rect 2678 1193 2694 1227
rect 2728 1193 2744 1227
rect 2678 1159 2744 1193
rect 2678 1125 2694 1159
rect 2728 1125 2744 1159
rect 2678 1091 2744 1125
rect 2678 1057 2694 1091
rect 2728 1057 2744 1091
rect 2678 1023 2744 1057
rect 2678 989 2694 1023
rect 2728 989 2744 1023
rect 2678 955 2744 989
rect 2678 921 2694 955
rect 2728 921 2744 955
rect 2678 887 2744 921
rect 2678 853 2694 887
rect 2728 853 2744 887
rect 2678 819 2744 853
rect 2678 785 2694 819
rect 2728 785 2744 819
rect 2678 751 2744 785
rect 2678 717 2694 751
rect 2728 717 2744 751
rect 2678 683 2744 717
rect 2678 649 2694 683
rect 2728 649 2744 683
rect 2678 615 2744 649
rect 2678 581 2694 615
rect 2728 581 2744 615
rect 2678 547 2744 581
rect 2678 513 2694 547
rect 2728 513 2744 547
rect 2678 479 2744 513
rect 2678 445 2694 479
rect 2728 445 2744 479
rect 2678 411 2744 445
rect 2678 377 2694 411
rect 2728 377 2744 411
rect 2678 343 2744 377
rect 2678 309 2694 343
rect 2728 309 2744 343
rect 2678 268 2744 309
rect 2774 1227 2840 1268
rect 2774 1193 2790 1227
rect 2824 1193 2840 1227
rect 2774 1159 2840 1193
rect 2774 1125 2790 1159
rect 2824 1125 2840 1159
rect 2774 1091 2840 1125
rect 2774 1057 2790 1091
rect 2824 1057 2840 1091
rect 2774 1023 2840 1057
rect 2774 989 2790 1023
rect 2824 989 2840 1023
rect 2774 955 2840 989
rect 2774 921 2790 955
rect 2824 921 2840 955
rect 2774 887 2840 921
rect 2774 853 2790 887
rect 2824 853 2840 887
rect 2774 819 2840 853
rect 2774 785 2790 819
rect 2824 785 2840 819
rect 2774 751 2840 785
rect 2774 717 2790 751
rect 2824 717 2840 751
rect 2774 683 2840 717
rect 2774 649 2790 683
rect 2824 649 2840 683
rect 2774 615 2840 649
rect 2774 581 2790 615
rect 2824 581 2840 615
rect 2774 547 2840 581
rect 2774 513 2790 547
rect 2824 513 2840 547
rect 2774 479 2840 513
rect 2774 445 2790 479
rect 2824 445 2840 479
rect 2774 411 2840 445
rect 2774 377 2790 411
rect 2824 377 2840 411
rect 2774 343 2840 377
rect 2774 309 2790 343
rect 2824 309 2840 343
rect 2774 268 2840 309
rect 2870 1227 2936 1268
rect 2870 1193 2886 1227
rect 2920 1193 2936 1227
rect 2870 1159 2936 1193
rect 2870 1125 2886 1159
rect 2920 1125 2936 1159
rect 2870 1091 2936 1125
rect 2870 1057 2886 1091
rect 2920 1057 2936 1091
rect 2870 1023 2936 1057
rect 2870 989 2886 1023
rect 2920 989 2936 1023
rect 2870 955 2936 989
rect 2870 921 2886 955
rect 2920 921 2936 955
rect 2870 887 2936 921
rect 2870 853 2886 887
rect 2920 853 2936 887
rect 2870 819 2936 853
rect 2870 785 2886 819
rect 2920 785 2936 819
rect 2870 751 2936 785
rect 2870 717 2886 751
rect 2920 717 2936 751
rect 2870 683 2936 717
rect 2870 649 2886 683
rect 2920 649 2936 683
rect 2870 615 2936 649
rect 2870 581 2886 615
rect 2920 581 2936 615
rect 2870 547 2936 581
rect 2870 513 2886 547
rect 2920 513 2936 547
rect 2870 479 2936 513
rect 2870 445 2886 479
rect 2920 445 2936 479
rect 2870 411 2936 445
rect 2870 377 2886 411
rect 2920 377 2936 411
rect 2870 343 2936 377
rect 2870 309 2886 343
rect 2920 309 2936 343
rect 2870 268 2936 309
rect 2966 1227 3028 1268
rect 2966 1193 2982 1227
rect 3016 1193 3028 1227
rect 2966 1159 3028 1193
rect 2966 1125 2982 1159
rect 3016 1125 3028 1159
rect 2966 1091 3028 1125
rect 2966 1057 2982 1091
rect 3016 1057 3028 1091
rect 2966 1023 3028 1057
rect 2966 989 2982 1023
rect 3016 989 3028 1023
rect 2966 955 3028 989
rect 2966 921 2982 955
rect 3016 921 3028 955
rect 2966 887 3028 921
rect 2966 853 2982 887
rect 3016 853 3028 887
rect 2966 819 3028 853
rect 2966 785 2982 819
rect 3016 785 3028 819
rect 2966 751 3028 785
rect 2966 717 2982 751
rect 3016 717 3028 751
rect 2966 683 3028 717
rect 2966 649 2982 683
rect 3016 649 3028 683
rect 2966 615 3028 649
rect 2966 581 2982 615
rect 3016 581 3028 615
rect 2966 547 3028 581
rect 2966 513 2982 547
rect 3016 513 3028 547
rect 2966 479 3028 513
rect 2966 445 2982 479
rect 3016 445 3028 479
rect 2966 411 3028 445
rect 2966 377 2982 411
rect 3016 377 3028 411
rect 2966 343 3028 377
rect 2966 309 2982 343
rect 3016 309 3028 343
rect 2966 268 3028 309
rect 3102 1211 3164 1252
rect 3102 1177 3114 1211
rect 3148 1177 3164 1211
rect 3102 1143 3164 1177
rect 3102 1109 3114 1143
rect 3148 1109 3164 1143
rect 3102 1075 3164 1109
rect 3102 1041 3114 1075
rect 3148 1041 3164 1075
rect 3102 1007 3164 1041
rect 3102 973 3114 1007
rect 3148 973 3164 1007
rect 3102 939 3164 973
rect 3102 905 3114 939
rect 3148 905 3164 939
rect 3102 871 3164 905
rect 3102 837 3114 871
rect 3148 837 3164 871
rect 3102 803 3164 837
rect 3102 769 3114 803
rect 3148 769 3164 803
rect 3102 735 3164 769
rect 3102 701 3114 735
rect 3148 701 3164 735
rect 3102 667 3164 701
rect 3102 633 3114 667
rect 3148 633 3164 667
rect 3102 599 3164 633
rect 3102 565 3114 599
rect 3148 565 3164 599
rect 3102 531 3164 565
rect 3102 497 3114 531
rect 3148 497 3164 531
rect 3102 463 3164 497
rect 3102 429 3114 463
rect 3148 429 3164 463
rect 3102 395 3164 429
rect 3102 361 3114 395
rect 3148 361 3164 395
rect 3102 327 3164 361
rect 3102 293 3114 327
rect 3148 293 3164 327
rect -914 209 -856 243
rect -914 175 -902 209
rect -868 175 -856 209
rect -914 141 -856 175
rect 3102 252 3164 293
rect 3194 1211 3260 1252
rect 3194 1177 3210 1211
rect 3244 1177 3260 1211
rect 3194 1143 3260 1177
rect 3194 1109 3210 1143
rect 3244 1109 3260 1143
rect 3194 1075 3260 1109
rect 3194 1041 3210 1075
rect 3244 1041 3260 1075
rect 3194 1007 3260 1041
rect 3194 973 3210 1007
rect 3244 973 3260 1007
rect 3194 939 3260 973
rect 3194 905 3210 939
rect 3244 905 3260 939
rect 3194 871 3260 905
rect 3194 837 3210 871
rect 3244 837 3260 871
rect 3194 803 3260 837
rect 3194 769 3210 803
rect 3244 769 3260 803
rect 3194 735 3260 769
rect 3194 701 3210 735
rect 3244 701 3260 735
rect 3194 667 3260 701
rect 3194 633 3210 667
rect 3244 633 3260 667
rect 3194 599 3260 633
rect 3194 565 3210 599
rect 3244 565 3260 599
rect 3194 531 3260 565
rect 3194 497 3210 531
rect 3244 497 3260 531
rect 3194 463 3260 497
rect 3194 429 3210 463
rect 3244 429 3260 463
rect 3194 395 3260 429
rect 3194 361 3210 395
rect 3244 361 3260 395
rect 3194 327 3260 361
rect 3194 293 3210 327
rect 3244 293 3260 327
rect 3194 252 3260 293
rect 3290 1211 3356 1252
rect 3290 1177 3306 1211
rect 3340 1177 3356 1211
rect 3290 1143 3356 1177
rect 3290 1109 3306 1143
rect 3340 1109 3356 1143
rect 3290 1075 3356 1109
rect 3290 1041 3306 1075
rect 3340 1041 3356 1075
rect 3290 1007 3356 1041
rect 3290 973 3306 1007
rect 3340 973 3356 1007
rect 3290 939 3356 973
rect 3290 905 3306 939
rect 3340 905 3356 939
rect 3290 871 3356 905
rect 3290 837 3306 871
rect 3340 837 3356 871
rect 3290 803 3356 837
rect 3290 769 3306 803
rect 3340 769 3356 803
rect 3290 735 3356 769
rect 3290 701 3306 735
rect 3340 701 3356 735
rect 3290 667 3356 701
rect 3290 633 3306 667
rect 3340 633 3356 667
rect 3290 599 3356 633
rect 3290 565 3306 599
rect 3340 565 3356 599
rect 3290 531 3356 565
rect 3290 497 3306 531
rect 3340 497 3356 531
rect 3290 463 3356 497
rect 3290 429 3306 463
rect 3340 429 3356 463
rect 3290 395 3356 429
rect 3290 361 3306 395
rect 3340 361 3356 395
rect 3290 327 3356 361
rect 3290 293 3306 327
rect 3340 293 3356 327
rect 3290 252 3356 293
rect 3386 1211 3452 1252
rect 3386 1177 3402 1211
rect 3436 1177 3452 1211
rect 3386 1143 3452 1177
rect 3386 1109 3402 1143
rect 3436 1109 3452 1143
rect 3386 1075 3452 1109
rect 3386 1041 3402 1075
rect 3436 1041 3452 1075
rect 3386 1007 3452 1041
rect 3386 973 3402 1007
rect 3436 973 3452 1007
rect 3386 939 3452 973
rect 3386 905 3402 939
rect 3436 905 3452 939
rect 3386 871 3452 905
rect 3386 837 3402 871
rect 3436 837 3452 871
rect 3386 803 3452 837
rect 3386 769 3402 803
rect 3436 769 3452 803
rect 3386 735 3452 769
rect 3386 701 3402 735
rect 3436 701 3452 735
rect 3386 667 3452 701
rect 3386 633 3402 667
rect 3436 633 3452 667
rect 3386 599 3452 633
rect 3386 565 3402 599
rect 3436 565 3452 599
rect 3386 531 3452 565
rect 3386 497 3402 531
rect 3436 497 3452 531
rect 3386 463 3452 497
rect 3386 429 3402 463
rect 3436 429 3452 463
rect 3386 395 3452 429
rect 3386 361 3402 395
rect 3436 361 3452 395
rect 3386 327 3452 361
rect 3386 293 3402 327
rect 3436 293 3452 327
rect 3386 252 3452 293
rect 3482 1211 3548 1252
rect 3482 1177 3498 1211
rect 3532 1177 3548 1211
rect 3482 1143 3548 1177
rect 3482 1109 3498 1143
rect 3532 1109 3548 1143
rect 3482 1075 3548 1109
rect 3482 1041 3498 1075
rect 3532 1041 3548 1075
rect 3482 1007 3548 1041
rect 3482 973 3498 1007
rect 3532 973 3548 1007
rect 3482 939 3548 973
rect 3482 905 3498 939
rect 3532 905 3548 939
rect 3482 871 3548 905
rect 3482 837 3498 871
rect 3532 837 3548 871
rect 3482 803 3548 837
rect 3482 769 3498 803
rect 3532 769 3548 803
rect 3482 735 3548 769
rect 3482 701 3498 735
rect 3532 701 3548 735
rect 3482 667 3548 701
rect 3482 633 3498 667
rect 3532 633 3548 667
rect 3482 599 3548 633
rect 3482 565 3498 599
rect 3532 565 3548 599
rect 3482 531 3548 565
rect 3482 497 3498 531
rect 3532 497 3548 531
rect 3482 463 3548 497
rect 3482 429 3498 463
rect 3532 429 3548 463
rect 3482 395 3548 429
rect 3482 361 3498 395
rect 3532 361 3548 395
rect 3482 327 3548 361
rect 3482 293 3498 327
rect 3532 293 3548 327
rect 3482 252 3548 293
rect 3578 1211 3644 1252
rect 3578 1177 3594 1211
rect 3628 1177 3644 1211
rect 3578 1143 3644 1177
rect 3578 1109 3594 1143
rect 3628 1109 3644 1143
rect 3578 1075 3644 1109
rect 3578 1041 3594 1075
rect 3628 1041 3644 1075
rect 3578 1007 3644 1041
rect 3578 973 3594 1007
rect 3628 973 3644 1007
rect 3578 939 3644 973
rect 3578 905 3594 939
rect 3628 905 3644 939
rect 3578 871 3644 905
rect 3578 837 3594 871
rect 3628 837 3644 871
rect 3578 803 3644 837
rect 3578 769 3594 803
rect 3628 769 3644 803
rect 3578 735 3644 769
rect 3578 701 3594 735
rect 3628 701 3644 735
rect 3578 667 3644 701
rect 3578 633 3594 667
rect 3628 633 3644 667
rect 3578 599 3644 633
rect 3578 565 3594 599
rect 3628 565 3644 599
rect 3578 531 3644 565
rect 3578 497 3594 531
rect 3628 497 3644 531
rect 3578 463 3644 497
rect 3578 429 3594 463
rect 3628 429 3644 463
rect 3578 395 3644 429
rect 3578 361 3594 395
rect 3628 361 3644 395
rect 3578 327 3644 361
rect 3578 293 3594 327
rect 3628 293 3644 327
rect 3578 252 3644 293
rect 3674 1211 3740 1252
rect 3674 1177 3690 1211
rect 3724 1177 3740 1211
rect 3674 1143 3740 1177
rect 3674 1109 3690 1143
rect 3724 1109 3740 1143
rect 3674 1075 3740 1109
rect 3674 1041 3690 1075
rect 3724 1041 3740 1075
rect 3674 1007 3740 1041
rect 3674 973 3690 1007
rect 3724 973 3740 1007
rect 3674 939 3740 973
rect 3674 905 3690 939
rect 3724 905 3740 939
rect 3674 871 3740 905
rect 3674 837 3690 871
rect 3724 837 3740 871
rect 3674 803 3740 837
rect 3674 769 3690 803
rect 3724 769 3740 803
rect 3674 735 3740 769
rect 3674 701 3690 735
rect 3724 701 3740 735
rect 3674 667 3740 701
rect 3674 633 3690 667
rect 3724 633 3740 667
rect 3674 599 3740 633
rect 3674 565 3690 599
rect 3724 565 3740 599
rect 3674 531 3740 565
rect 3674 497 3690 531
rect 3724 497 3740 531
rect 3674 463 3740 497
rect 3674 429 3690 463
rect 3724 429 3740 463
rect 3674 395 3740 429
rect 3674 361 3690 395
rect 3724 361 3740 395
rect 3674 327 3740 361
rect 3674 293 3690 327
rect 3724 293 3740 327
rect 3674 252 3740 293
rect 3770 1211 3836 1252
rect 3770 1177 3786 1211
rect 3820 1177 3836 1211
rect 3770 1143 3836 1177
rect 3770 1109 3786 1143
rect 3820 1109 3836 1143
rect 3770 1075 3836 1109
rect 3770 1041 3786 1075
rect 3820 1041 3836 1075
rect 3770 1007 3836 1041
rect 3770 973 3786 1007
rect 3820 973 3836 1007
rect 3770 939 3836 973
rect 3770 905 3786 939
rect 3820 905 3836 939
rect 3770 871 3836 905
rect 3770 837 3786 871
rect 3820 837 3836 871
rect 3770 803 3836 837
rect 3770 769 3786 803
rect 3820 769 3836 803
rect 3770 735 3836 769
rect 3770 701 3786 735
rect 3820 701 3836 735
rect 3770 667 3836 701
rect 3770 633 3786 667
rect 3820 633 3836 667
rect 3770 599 3836 633
rect 3770 565 3786 599
rect 3820 565 3836 599
rect 3770 531 3836 565
rect 3770 497 3786 531
rect 3820 497 3836 531
rect 3770 463 3836 497
rect 3770 429 3786 463
rect 3820 429 3836 463
rect 3770 395 3836 429
rect 3770 361 3786 395
rect 3820 361 3836 395
rect 3770 327 3836 361
rect 3770 293 3786 327
rect 3820 293 3836 327
rect 3770 252 3836 293
rect 3866 1211 3932 1252
rect 3866 1177 3882 1211
rect 3916 1177 3932 1211
rect 3866 1143 3932 1177
rect 3866 1109 3882 1143
rect 3916 1109 3932 1143
rect 3866 1075 3932 1109
rect 3866 1041 3882 1075
rect 3916 1041 3932 1075
rect 3866 1007 3932 1041
rect 3866 973 3882 1007
rect 3916 973 3932 1007
rect 3866 939 3932 973
rect 3866 905 3882 939
rect 3916 905 3932 939
rect 3866 871 3932 905
rect 3866 837 3882 871
rect 3916 837 3932 871
rect 3866 803 3932 837
rect 3866 769 3882 803
rect 3916 769 3932 803
rect 3866 735 3932 769
rect 3866 701 3882 735
rect 3916 701 3932 735
rect 3866 667 3932 701
rect 3866 633 3882 667
rect 3916 633 3932 667
rect 3866 599 3932 633
rect 3866 565 3882 599
rect 3916 565 3932 599
rect 3866 531 3932 565
rect 3866 497 3882 531
rect 3916 497 3932 531
rect 3866 463 3932 497
rect 3866 429 3882 463
rect 3916 429 3932 463
rect 3866 395 3932 429
rect 3866 361 3882 395
rect 3916 361 3932 395
rect 3866 327 3932 361
rect 3866 293 3882 327
rect 3916 293 3932 327
rect 3866 252 3932 293
rect 3962 1211 4028 1252
rect 3962 1177 3978 1211
rect 4012 1177 4028 1211
rect 3962 1143 4028 1177
rect 3962 1109 3978 1143
rect 4012 1109 4028 1143
rect 3962 1075 4028 1109
rect 3962 1041 3978 1075
rect 4012 1041 4028 1075
rect 3962 1007 4028 1041
rect 3962 973 3978 1007
rect 4012 973 4028 1007
rect 3962 939 4028 973
rect 3962 905 3978 939
rect 4012 905 4028 939
rect 3962 871 4028 905
rect 3962 837 3978 871
rect 4012 837 4028 871
rect 3962 803 4028 837
rect 3962 769 3978 803
rect 4012 769 4028 803
rect 3962 735 4028 769
rect 3962 701 3978 735
rect 4012 701 4028 735
rect 3962 667 4028 701
rect 3962 633 3978 667
rect 4012 633 4028 667
rect 3962 599 4028 633
rect 3962 565 3978 599
rect 4012 565 4028 599
rect 3962 531 4028 565
rect 3962 497 3978 531
rect 4012 497 4028 531
rect 3962 463 4028 497
rect 3962 429 3978 463
rect 4012 429 4028 463
rect 3962 395 4028 429
rect 3962 361 3978 395
rect 4012 361 4028 395
rect 3962 327 4028 361
rect 3962 293 3978 327
rect 4012 293 4028 327
rect 3962 252 4028 293
rect 4058 1211 4124 1252
rect 4058 1177 4074 1211
rect 4108 1177 4124 1211
rect 4058 1143 4124 1177
rect 4058 1109 4074 1143
rect 4108 1109 4124 1143
rect 4058 1075 4124 1109
rect 4058 1041 4074 1075
rect 4108 1041 4124 1075
rect 4058 1007 4124 1041
rect 4058 973 4074 1007
rect 4108 973 4124 1007
rect 4058 939 4124 973
rect 4058 905 4074 939
rect 4108 905 4124 939
rect 4058 871 4124 905
rect 4058 837 4074 871
rect 4108 837 4124 871
rect 4058 803 4124 837
rect 4058 769 4074 803
rect 4108 769 4124 803
rect 4058 735 4124 769
rect 4058 701 4074 735
rect 4108 701 4124 735
rect 4058 667 4124 701
rect 4058 633 4074 667
rect 4108 633 4124 667
rect 4058 599 4124 633
rect 4058 565 4074 599
rect 4108 565 4124 599
rect 4058 531 4124 565
rect 4058 497 4074 531
rect 4108 497 4124 531
rect 4058 463 4124 497
rect 4058 429 4074 463
rect 4108 429 4124 463
rect 4058 395 4124 429
rect 4058 361 4074 395
rect 4108 361 4124 395
rect 4058 327 4124 361
rect 4058 293 4074 327
rect 4108 293 4124 327
rect 4058 252 4124 293
rect 4154 1211 4220 1252
rect 4154 1177 4170 1211
rect 4204 1177 4220 1211
rect 4154 1143 4220 1177
rect 4154 1109 4170 1143
rect 4204 1109 4220 1143
rect 4154 1075 4220 1109
rect 4154 1041 4170 1075
rect 4204 1041 4220 1075
rect 4154 1007 4220 1041
rect 4154 973 4170 1007
rect 4204 973 4220 1007
rect 4154 939 4220 973
rect 4154 905 4170 939
rect 4204 905 4220 939
rect 4154 871 4220 905
rect 4154 837 4170 871
rect 4204 837 4220 871
rect 4154 803 4220 837
rect 4154 769 4170 803
rect 4204 769 4220 803
rect 4154 735 4220 769
rect 4154 701 4170 735
rect 4204 701 4220 735
rect 4154 667 4220 701
rect 4154 633 4170 667
rect 4204 633 4220 667
rect 4154 599 4220 633
rect 4154 565 4170 599
rect 4204 565 4220 599
rect 4154 531 4220 565
rect 4154 497 4170 531
rect 4204 497 4220 531
rect 4154 463 4220 497
rect 4154 429 4170 463
rect 4204 429 4220 463
rect 4154 395 4220 429
rect 4154 361 4170 395
rect 4204 361 4220 395
rect 4154 327 4220 361
rect 4154 293 4170 327
rect 4204 293 4220 327
rect 4154 252 4220 293
rect 4250 1211 4312 1252
rect 4250 1177 4266 1211
rect 4300 1177 4312 1211
rect 4250 1143 4312 1177
rect 4250 1109 4266 1143
rect 4300 1109 4312 1143
rect 4250 1075 4312 1109
rect 4250 1041 4266 1075
rect 4300 1041 4312 1075
rect 4250 1007 4312 1041
rect 4250 973 4266 1007
rect 4300 973 4312 1007
rect 4250 939 4312 973
rect 4250 905 4266 939
rect 4300 905 4312 939
rect 4250 871 4312 905
rect 4250 837 4266 871
rect 4300 837 4312 871
rect 4250 803 4312 837
rect 4250 769 4266 803
rect 4300 769 4312 803
rect 4250 735 4312 769
rect 4250 701 4266 735
rect 4300 701 4312 735
rect 4250 667 4312 701
rect 4250 633 4266 667
rect 4300 633 4312 667
rect 4250 599 4312 633
rect 4250 565 4266 599
rect 4300 565 4312 599
rect 4250 531 4312 565
rect 4250 497 4266 531
rect 4300 497 4312 531
rect 4250 463 4312 497
rect 4250 429 4266 463
rect 4300 429 4312 463
rect 4250 395 4312 429
rect 4250 361 4266 395
rect 4300 361 4312 395
rect 4250 327 4312 361
rect 4250 293 4266 327
rect 4300 293 4312 327
rect 4250 252 4312 293
rect 4870 1211 4932 1252
rect 4870 1177 4882 1211
rect 4916 1177 4932 1211
rect 4870 1143 4932 1177
rect 4870 1109 4882 1143
rect 4916 1109 4932 1143
rect 4870 1075 4932 1109
rect 4870 1041 4882 1075
rect 4916 1041 4932 1075
rect 4870 1007 4932 1041
rect 4870 973 4882 1007
rect 4916 973 4932 1007
rect 4870 939 4932 973
rect 4870 905 4882 939
rect 4916 905 4932 939
rect 4870 871 4932 905
rect 4870 837 4882 871
rect 4916 837 4932 871
rect 4870 803 4932 837
rect 4870 769 4882 803
rect 4916 769 4932 803
rect 4870 735 4932 769
rect 4870 701 4882 735
rect 4916 701 4932 735
rect 4870 667 4932 701
rect 4870 633 4882 667
rect 4916 633 4932 667
rect 4870 599 4932 633
rect 4870 565 4882 599
rect 4916 565 4932 599
rect 4870 531 4932 565
rect 4870 497 4882 531
rect 4916 497 4932 531
rect 4870 463 4932 497
rect 4870 429 4882 463
rect 4916 429 4932 463
rect 4870 395 4932 429
rect 4870 361 4882 395
rect 4916 361 4932 395
rect 4870 327 4932 361
rect 4870 293 4882 327
rect 4916 293 4932 327
rect 4870 252 4932 293
rect 4962 1211 5028 1252
rect 4962 1177 4978 1211
rect 5012 1177 5028 1211
rect 4962 1143 5028 1177
rect 4962 1109 4978 1143
rect 5012 1109 5028 1143
rect 4962 1075 5028 1109
rect 4962 1041 4978 1075
rect 5012 1041 5028 1075
rect 4962 1007 5028 1041
rect 4962 973 4978 1007
rect 5012 973 5028 1007
rect 4962 939 5028 973
rect 4962 905 4978 939
rect 5012 905 5028 939
rect 4962 871 5028 905
rect 4962 837 4978 871
rect 5012 837 5028 871
rect 4962 803 5028 837
rect 4962 769 4978 803
rect 5012 769 5028 803
rect 4962 735 5028 769
rect 4962 701 4978 735
rect 5012 701 5028 735
rect 4962 667 5028 701
rect 4962 633 4978 667
rect 5012 633 5028 667
rect 4962 599 5028 633
rect 4962 565 4978 599
rect 5012 565 5028 599
rect 4962 531 5028 565
rect 4962 497 4978 531
rect 5012 497 5028 531
rect 4962 463 5028 497
rect 4962 429 4978 463
rect 5012 429 5028 463
rect 4962 395 5028 429
rect 4962 361 4978 395
rect 5012 361 5028 395
rect 4962 327 5028 361
rect 4962 293 4978 327
rect 5012 293 5028 327
rect 4962 252 5028 293
rect 5058 1211 5124 1252
rect 5058 1177 5074 1211
rect 5108 1177 5124 1211
rect 5058 1143 5124 1177
rect 5058 1109 5074 1143
rect 5108 1109 5124 1143
rect 5058 1075 5124 1109
rect 5058 1041 5074 1075
rect 5108 1041 5124 1075
rect 5058 1007 5124 1041
rect 5058 973 5074 1007
rect 5108 973 5124 1007
rect 5058 939 5124 973
rect 5058 905 5074 939
rect 5108 905 5124 939
rect 5058 871 5124 905
rect 5058 837 5074 871
rect 5108 837 5124 871
rect 5058 803 5124 837
rect 5058 769 5074 803
rect 5108 769 5124 803
rect 5058 735 5124 769
rect 5058 701 5074 735
rect 5108 701 5124 735
rect 5058 667 5124 701
rect 5058 633 5074 667
rect 5108 633 5124 667
rect 5058 599 5124 633
rect 5058 565 5074 599
rect 5108 565 5124 599
rect 5058 531 5124 565
rect 5058 497 5074 531
rect 5108 497 5124 531
rect 5058 463 5124 497
rect 5058 429 5074 463
rect 5108 429 5124 463
rect 5058 395 5124 429
rect 5058 361 5074 395
rect 5108 361 5124 395
rect 5058 327 5124 361
rect 5058 293 5074 327
rect 5108 293 5124 327
rect 5058 252 5124 293
rect 5154 1211 5220 1252
rect 5154 1177 5170 1211
rect 5204 1177 5220 1211
rect 5154 1143 5220 1177
rect 5154 1109 5170 1143
rect 5204 1109 5220 1143
rect 5154 1075 5220 1109
rect 5154 1041 5170 1075
rect 5204 1041 5220 1075
rect 5154 1007 5220 1041
rect 5154 973 5170 1007
rect 5204 973 5220 1007
rect 5154 939 5220 973
rect 5154 905 5170 939
rect 5204 905 5220 939
rect 5154 871 5220 905
rect 5154 837 5170 871
rect 5204 837 5220 871
rect 5154 803 5220 837
rect 5154 769 5170 803
rect 5204 769 5220 803
rect 5154 735 5220 769
rect 5154 701 5170 735
rect 5204 701 5220 735
rect 5154 667 5220 701
rect 5154 633 5170 667
rect 5204 633 5220 667
rect 5154 599 5220 633
rect 5154 565 5170 599
rect 5204 565 5220 599
rect 5154 531 5220 565
rect 5154 497 5170 531
rect 5204 497 5220 531
rect 5154 463 5220 497
rect 5154 429 5170 463
rect 5204 429 5220 463
rect 5154 395 5220 429
rect 5154 361 5170 395
rect 5204 361 5220 395
rect 5154 327 5220 361
rect 5154 293 5170 327
rect 5204 293 5220 327
rect 5154 252 5220 293
rect 5250 1211 5316 1252
rect 5250 1177 5266 1211
rect 5300 1177 5316 1211
rect 5250 1143 5316 1177
rect 5250 1109 5266 1143
rect 5300 1109 5316 1143
rect 5250 1075 5316 1109
rect 5250 1041 5266 1075
rect 5300 1041 5316 1075
rect 5250 1007 5316 1041
rect 5250 973 5266 1007
rect 5300 973 5316 1007
rect 5250 939 5316 973
rect 5250 905 5266 939
rect 5300 905 5316 939
rect 5250 871 5316 905
rect 5250 837 5266 871
rect 5300 837 5316 871
rect 5250 803 5316 837
rect 5250 769 5266 803
rect 5300 769 5316 803
rect 5250 735 5316 769
rect 5250 701 5266 735
rect 5300 701 5316 735
rect 5250 667 5316 701
rect 5250 633 5266 667
rect 5300 633 5316 667
rect 5250 599 5316 633
rect 5250 565 5266 599
rect 5300 565 5316 599
rect 5250 531 5316 565
rect 5250 497 5266 531
rect 5300 497 5316 531
rect 5250 463 5316 497
rect 5250 429 5266 463
rect 5300 429 5316 463
rect 5250 395 5316 429
rect 5250 361 5266 395
rect 5300 361 5316 395
rect 5250 327 5316 361
rect 5250 293 5266 327
rect 5300 293 5316 327
rect 5250 252 5316 293
rect 5346 1211 5412 1252
rect 5346 1177 5362 1211
rect 5396 1177 5412 1211
rect 5346 1143 5412 1177
rect 5346 1109 5362 1143
rect 5396 1109 5412 1143
rect 5346 1075 5412 1109
rect 5346 1041 5362 1075
rect 5396 1041 5412 1075
rect 5346 1007 5412 1041
rect 5346 973 5362 1007
rect 5396 973 5412 1007
rect 5346 939 5412 973
rect 5346 905 5362 939
rect 5396 905 5412 939
rect 5346 871 5412 905
rect 5346 837 5362 871
rect 5396 837 5412 871
rect 5346 803 5412 837
rect 5346 769 5362 803
rect 5396 769 5412 803
rect 5346 735 5412 769
rect 5346 701 5362 735
rect 5396 701 5412 735
rect 5346 667 5412 701
rect 5346 633 5362 667
rect 5396 633 5412 667
rect 5346 599 5412 633
rect 5346 565 5362 599
rect 5396 565 5412 599
rect 5346 531 5412 565
rect 5346 497 5362 531
rect 5396 497 5412 531
rect 5346 463 5412 497
rect 5346 429 5362 463
rect 5396 429 5412 463
rect 5346 395 5412 429
rect 5346 361 5362 395
rect 5396 361 5412 395
rect 5346 327 5412 361
rect 5346 293 5362 327
rect 5396 293 5412 327
rect 5346 252 5412 293
rect 5442 1211 5508 1252
rect 5442 1177 5458 1211
rect 5492 1177 5508 1211
rect 5442 1143 5508 1177
rect 5442 1109 5458 1143
rect 5492 1109 5508 1143
rect 5442 1075 5508 1109
rect 5442 1041 5458 1075
rect 5492 1041 5508 1075
rect 5442 1007 5508 1041
rect 5442 973 5458 1007
rect 5492 973 5508 1007
rect 5442 939 5508 973
rect 5442 905 5458 939
rect 5492 905 5508 939
rect 5442 871 5508 905
rect 5442 837 5458 871
rect 5492 837 5508 871
rect 5442 803 5508 837
rect 5442 769 5458 803
rect 5492 769 5508 803
rect 5442 735 5508 769
rect 5442 701 5458 735
rect 5492 701 5508 735
rect 5442 667 5508 701
rect 5442 633 5458 667
rect 5492 633 5508 667
rect 5442 599 5508 633
rect 5442 565 5458 599
rect 5492 565 5508 599
rect 5442 531 5508 565
rect 5442 497 5458 531
rect 5492 497 5508 531
rect 5442 463 5508 497
rect 5442 429 5458 463
rect 5492 429 5508 463
rect 5442 395 5508 429
rect 5442 361 5458 395
rect 5492 361 5508 395
rect 5442 327 5508 361
rect 5442 293 5458 327
rect 5492 293 5508 327
rect 5442 252 5508 293
rect 5538 1211 5604 1252
rect 5538 1177 5554 1211
rect 5588 1177 5604 1211
rect 5538 1143 5604 1177
rect 5538 1109 5554 1143
rect 5588 1109 5604 1143
rect 5538 1075 5604 1109
rect 5538 1041 5554 1075
rect 5588 1041 5604 1075
rect 5538 1007 5604 1041
rect 5538 973 5554 1007
rect 5588 973 5604 1007
rect 5538 939 5604 973
rect 5538 905 5554 939
rect 5588 905 5604 939
rect 5538 871 5604 905
rect 5538 837 5554 871
rect 5588 837 5604 871
rect 5538 803 5604 837
rect 5538 769 5554 803
rect 5588 769 5604 803
rect 5538 735 5604 769
rect 5538 701 5554 735
rect 5588 701 5604 735
rect 5538 667 5604 701
rect 5538 633 5554 667
rect 5588 633 5604 667
rect 5538 599 5604 633
rect 5538 565 5554 599
rect 5588 565 5604 599
rect 5538 531 5604 565
rect 5538 497 5554 531
rect 5588 497 5604 531
rect 5538 463 5604 497
rect 5538 429 5554 463
rect 5588 429 5604 463
rect 5538 395 5604 429
rect 5538 361 5554 395
rect 5588 361 5604 395
rect 5538 327 5604 361
rect 5538 293 5554 327
rect 5588 293 5604 327
rect 5538 252 5604 293
rect 5634 1211 5700 1252
rect 5634 1177 5650 1211
rect 5684 1177 5700 1211
rect 5634 1143 5700 1177
rect 5634 1109 5650 1143
rect 5684 1109 5700 1143
rect 5634 1075 5700 1109
rect 5634 1041 5650 1075
rect 5684 1041 5700 1075
rect 5634 1007 5700 1041
rect 5634 973 5650 1007
rect 5684 973 5700 1007
rect 5634 939 5700 973
rect 5634 905 5650 939
rect 5684 905 5700 939
rect 5634 871 5700 905
rect 5634 837 5650 871
rect 5684 837 5700 871
rect 5634 803 5700 837
rect 5634 769 5650 803
rect 5684 769 5700 803
rect 5634 735 5700 769
rect 5634 701 5650 735
rect 5684 701 5700 735
rect 5634 667 5700 701
rect 5634 633 5650 667
rect 5684 633 5700 667
rect 5634 599 5700 633
rect 5634 565 5650 599
rect 5684 565 5700 599
rect 5634 531 5700 565
rect 5634 497 5650 531
rect 5684 497 5700 531
rect 5634 463 5700 497
rect 5634 429 5650 463
rect 5684 429 5700 463
rect 5634 395 5700 429
rect 5634 361 5650 395
rect 5684 361 5700 395
rect 5634 327 5700 361
rect 5634 293 5650 327
rect 5684 293 5700 327
rect 5634 252 5700 293
rect 5730 1211 5796 1252
rect 5730 1177 5746 1211
rect 5780 1177 5796 1211
rect 5730 1143 5796 1177
rect 5730 1109 5746 1143
rect 5780 1109 5796 1143
rect 5730 1075 5796 1109
rect 5730 1041 5746 1075
rect 5780 1041 5796 1075
rect 5730 1007 5796 1041
rect 5730 973 5746 1007
rect 5780 973 5796 1007
rect 5730 939 5796 973
rect 5730 905 5746 939
rect 5780 905 5796 939
rect 5730 871 5796 905
rect 5730 837 5746 871
rect 5780 837 5796 871
rect 5730 803 5796 837
rect 5730 769 5746 803
rect 5780 769 5796 803
rect 5730 735 5796 769
rect 5730 701 5746 735
rect 5780 701 5796 735
rect 5730 667 5796 701
rect 5730 633 5746 667
rect 5780 633 5796 667
rect 5730 599 5796 633
rect 5730 565 5746 599
rect 5780 565 5796 599
rect 5730 531 5796 565
rect 5730 497 5746 531
rect 5780 497 5796 531
rect 5730 463 5796 497
rect 5730 429 5746 463
rect 5780 429 5796 463
rect 5730 395 5796 429
rect 5730 361 5746 395
rect 5780 361 5796 395
rect 5730 327 5796 361
rect 5730 293 5746 327
rect 5780 293 5796 327
rect 5730 252 5796 293
rect 5826 1211 5892 1252
rect 5826 1177 5842 1211
rect 5876 1177 5892 1211
rect 5826 1143 5892 1177
rect 5826 1109 5842 1143
rect 5876 1109 5892 1143
rect 5826 1075 5892 1109
rect 5826 1041 5842 1075
rect 5876 1041 5892 1075
rect 5826 1007 5892 1041
rect 5826 973 5842 1007
rect 5876 973 5892 1007
rect 5826 939 5892 973
rect 5826 905 5842 939
rect 5876 905 5892 939
rect 5826 871 5892 905
rect 5826 837 5842 871
rect 5876 837 5892 871
rect 5826 803 5892 837
rect 5826 769 5842 803
rect 5876 769 5892 803
rect 5826 735 5892 769
rect 5826 701 5842 735
rect 5876 701 5892 735
rect 5826 667 5892 701
rect 5826 633 5842 667
rect 5876 633 5892 667
rect 5826 599 5892 633
rect 5826 565 5842 599
rect 5876 565 5892 599
rect 5826 531 5892 565
rect 5826 497 5842 531
rect 5876 497 5892 531
rect 5826 463 5892 497
rect 5826 429 5842 463
rect 5876 429 5892 463
rect 5826 395 5892 429
rect 5826 361 5842 395
rect 5876 361 5892 395
rect 5826 327 5892 361
rect 5826 293 5842 327
rect 5876 293 5892 327
rect 5826 252 5892 293
rect 5922 1211 5984 1252
rect 5922 1177 5938 1211
rect 5972 1177 5984 1211
rect 5922 1143 5984 1177
rect 5922 1109 5938 1143
rect 5972 1109 5984 1143
rect 5922 1075 5984 1109
rect 5922 1041 5938 1075
rect 5972 1041 5984 1075
rect 5922 1007 5984 1041
rect 5922 973 5938 1007
rect 5972 973 5984 1007
rect 5922 939 5984 973
rect 5922 905 5938 939
rect 5972 905 5984 939
rect 5922 871 5984 905
rect 5922 837 5938 871
rect 5972 837 5984 871
rect 5922 803 5984 837
rect 5922 769 5938 803
rect 5972 769 5984 803
rect 5922 735 5984 769
rect 5922 701 5938 735
rect 5972 701 5984 735
rect 5922 667 5984 701
rect 5922 633 5938 667
rect 5972 633 5984 667
rect 5922 599 5984 633
rect 5922 565 5938 599
rect 5972 565 5984 599
rect 5922 531 5984 565
rect 5922 497 5938 531
rect 5972 497 5984 531
rect 5922 463 5984 497
rect 5922 429 5938 463
rect 5972 429 5984 463
rect 5922 395 5984 429
rect 5922 361 5938 395
rect 5972 361 5984 395
rect 5922 327 5984 361
rect 5922 293 5938 327
rect 5972 293 5984 327
rect 5922 252 5984 293
rect 6132 1211 6194 1252
rect 6132 1177 6144 1211
rect 6178 1177 6194 1211
rect 6132 1143 6194 1177
rect 6132 1109 6144 1143
rect 6178 1109 6194 1143
rect 6132 1075 6194 1109
rect 6132 1041 6144 1075
rect 6178 1041 6194 1075
rect 6132 1007 6194 1041
rect 6132 973 6144 1007
rect 6178 973 6194 1007
rect 6132 939 6194 973
rect 6132 905 6144 939
rect 6178 905 6194 939
rect 6132 871 6194 905
rect 6132 837 6144 871
rect 6178 837 6194 871
rect 6132 803 6194 837
rect 6132 769 6144 803
rect 6178 769 6194 803
rect 6132 735 6194 769
rect 6132 701 6144 735
rect 6178 701 6194 735
rect 6132 667 6194 701
rect 6132 633 6144 667
rect 6178 633 6194 667
rect 6132 599 6194 633
rect 6132 565 6144 599
rect 6178 565 6194 599
rect 6132 531 6194 565
rect 6132 497 6144 531
rect 6178 497 6194 531
rect 6132 463 6194 497
rect 6132 429 6144 463
rect 6178 429 6194 463
rect 6132 395 6194 429
rect 6132 361 6144 395
rect 6178 361 6194 395
rect 6132 327 6194 361
rect 6132 293 6144 327
rect 6178 293 6194 327
rect 6132 252 6194 293
rect 6224 1211 6290 1252
rect 6224 1177 6240 1211
rect 6274 1177 6290 1211
rect 6224 1143 6290 1177
rect 6224 1109 6240 1143
rect 6274 1109 6290 1143
rect 6224 1075 6290 1109
rect 6224 1041 6240 1075
rect 6274 1041 6290 1075
rect 6224 1007 6290 1041
rect 6224 973 6240 1007
rect 6274 973 6290 1007
rect 6224 939 6290 973
rect 6224 905 6240 939
rect 6274 905 6290 939
rect 6224 871 6290 905
rect 6224 837 6240 871
rect 6274 837 6290 871
rect 6224 803 6290 837
rect 6224 769 6240 803
rect 6274 769 6290 803
rect 6224 735 6290 769
rect 6224 701 6240 735
rect 6274 701 6290 735
rect 6224 667 6290 701
rect 6224 633 6240 667
rect 6274 633 6290 667
rect 6224 599 6290 633
rect 6224 565 6240 599
rect 6274 565 6290 599
rect 6224 531 6290 565
rect 6224 497 6240 531
rect 6274 497 6290 531
rect 6224 463 6290 497
rect 6224 429 6240 463
rect 6274 429 6290 463
rect 6224 395 6290 429
rect 6224 361 6240 395
rect 6274 361 6290 395
rect 6224 327 6290 361
rect 6224 293 6240 327
rect 6274 293 6290 327
rect 6224 252 6290 293
rect 6320 1211 6386 1252
rect 6320 1177 6336 1211
rect 6370 1177 6386 1211
rect 6320 1143 6386 1177
rect 6320 1109 6336 1143
rect 6370 1109 6386 1143
rect 6320 1075 6386 1109
rect 6320 1041 6336 1075
rect 6370 1041 6386 1075
rect 6320 1007 6386 1041
rect 6320 973 6336 1007
rect 6370 973 6386 1007
rect 6320 939 6386 973
rect 6320 905 6336 939
rect 6370 905 6386 939
rect 6320 871 6386 905
rect 6320 837 6336 871
rect 6370 837 6386 871
rect 6320 803 6386 837
rect 6320 769 6336 803
rect 6370 769 6386 803
rect 6320 735 6386 769
rect 6320 701 6336 735
rect 6370 701 6386 735
rect 6320 667 6386 701
rect 6320 633 6336 667
rect 6370 633 6386 667
rect 6320 599 6386 633
rect 6320 565 6336 599
rect 6370 565 6386 599
rect 6320 531 6386 565
rect 6320 497 6336 531
rect 6370 497 6386 531
rect 6320 463 6386 497
rect 6320 429 6336 463
rect 6370 429 6386 463
rect 6320 395 6386 429
rect 6320 361 6336 395
rect 6370 361 6386 395
rect 6320 327 6386 361
rect 6320 293 6336 327
rect 6370 293 6386 327
rect 6320 252 6386 293
rect 6416 1211 6482 1252
rect 6416 1177 6432 1211
rect 6466 1177 6482 1211
rect 6416 1143 6482 1177
rect 6416 1109 6432 1143
rect 6466 1109 6482 1143
rect 6416 1075 6482 1109
rect 6416 1041 6432 1075
rect 6466 1041 6482 1075
rect 6416 1007 6482 1041
rect 6416 973 6432 1007
rect 6466 973 6482 1007
rect 6416 939 6482 973
rect 6416 905 6432 939
rect 6466 905 6482 939
rect 6416 871 6482 905
rect 6416 837 6432 871
rect 6466 837 6482 871
rect 6416 803 6482 837
rect 6416 769 6432 803
rect 6466 769 6482 803
rect 6416 735 6482 769
rect 6416 701 6432 735
rect 6466 701 6482 735
rect 6416 667 6482 701
rect 6416 633 6432 667
rect 6466 633 6482 667
rect 6416 599 6482 633
rect 6416 565 6432 599
rect 6466 565 6482 599
rect 6416 531 6482 565
rect 6416 497 6432 531
rect 6466 497 6482 531
rect 6416 463 6482 497
rect 6416 429 6432 463
rect 6466 429 6482 463
rect 6416 395 6482 429
rect 6416 361 6432 395
rect 6466 361 6482 395
rect 6416 327 6482 361
rect 6416 293 6432 327
rect 6466 293 6482 327
rect 6416 252 6482 293
rect 6512 1211 6578 1252
rect 6512 1177 6528 1211
rect 6562 1177 6578 1211
rect 6512 1143 6578 1177
rect 6512 1109 6528 1143
rect 6562 1109 6578 1143
rect 6512 1075 6578 1109
rect 6512 1041 6528 1075
rect 6562 1041 6578 1075
rect 6512 1007 6578 1041
rect 6512 973 6528 1007
rect 6562 973 6578 1007
rect 6512 939 6578 973
rect 6512 905 6528 939
rect 6562 905 6578 939
rect 6512 871 6578 905
rect 6512 837 6528 871
rect 6562 837 6578 871
rect 6512 803 6578 837
rect 6512 769 6528 803
rect 6562 769 6578 803
rect 6512 735 6578 769
rect 6512 701 6528 735
rect 6562 701 6578 735
rect 6512 667 6578 701
rect 6512 633 6528 667
rect 6562 633 6578 667
rect 6512 599 6578 633
rect 6512 565 6528 599
rect 6562 565 6578 599
rect 6512 531 6578 565
rect 6512 497 6528 531
rect 6562 497 6578 531
rect 6512 463 6578 497
rect 6512 429 6528 463
rect 6562 429 6578 463
rect 6512 395 6578 429
rect 6512 361 6528 395
rect 6562 361 6578 395
rect 6512 327 6578 361
rect 6512 293 6528 327
rect 6562 293 6578 327
rect 6512 252 6578 293
rect 6608 1211 6674 1252
rect 6608 1177 6624 1211
rect 6658 1177 6674 1211
rect 6608 1143 6674 1177
rect 6608 1109 6624 1143
rect 6658 1109 6674 1143
rect 6608 1075 6674 1109
rect 6608 1041 6624 1075
rect 6658 1041 6674 1075
rect 6608 1007 6674 1041
rect 6608 973 6624 1007
rect 6658 973 6674 1007
rect 6608 939 6674 973
rect 6608 905 6624 939
rect 6658 905 6674 939
rect 6608 871 6674 905
rect 6608 837 6624 871
rect 6658 837 6674 871
rect 6608 803 6674 837
rect 6608 769 6624 803
rect 6658 769 6674 803
rect 6608 735 6674 769
rect 6608 701 6624 735
rect 6658 701 6674 735
rect 6608 667 6674 701
rect 6608 633 6624 667
rect 6658 633 6674 667
rect 6608 599 6674 633
rect 6608 565 6624 599
rect 6658 565 6674 599
rect 6608 531 6674 565
rect 6608 497 6624 531
rect 6658 497 6674 531
rect 6608 463 6674 497
rect 6608 429 6624 463
rect 6658 429 6674 463
rect 6608 395 6674 429
rect 6608 361 6624 395
rect 6658 361 6674 395
rect 6608 327 6674 361
rect 6608 293 6624 327
rect 6658 293 6674 327
rect 6608 252 6674 293
rect 6704 1211 6770 1252
rect 6704 1177 6720 1211
rect 6754 1177 6770 1211
rect 6704 1143 6770 1177
rect 6704 1109 6720 1143
rect 6754 1109 6770 1143
rect 6704 1075 6770 1109
rect 6704 1041 6720 1075
rect 6754 1041 6770 1075
rect 6704 1007 6770 1041
rect 6704 973 6720 1007
rect 6754 973 6770 1007
rect 6704 939 6770 973
rect 6704 905 6720 939
rect 6754 905 6770 939
rect 6704 871 6770 905
rect 6704 837 6720 871
rect 6754 837 6770 871
rect 6704 803 6770 837
rect 6704 769 6720 803
rect 6754 769 6770 803
rect 6704 735 6770 769
rect 6704 701 6720 735
rect 6754 701 6770 735
rect 6704 667 6770 701
rect 6704 633 6720 667
rect 6754 633 6770 667
rect 6704 599 6770 633
rect 6704 565 6720 599
rect 6754 565 6770 599
rect 6704 531 6770 565
rect 6704 497 6720 531
rect 6754 497 6770 531
rect 6704 463 6770 497
rect 6704 429 6720 463
rect 6754 429 6770 463
rect 6704 395 6770 429
rect 6704 361 6720 395
rect 6754 361 6770 395
rect 6704 327 6770 361
rect 6704 293 6720 327
rect 6754 293 6770 327
rect 6704 252 6770 293
rect 6800 1211 6866 1252
rect 6800 1177 6816 1211
rect 6850 1177 6866 1211
rect 6800 1143 6866 1177
rect 6800 1109 6816 1143
rect 6850 1109 6866 1143
rect 6800 1075 6866 1109
rect 6800 1041 6816 1075
rect 6850 1041 6866 1075
rect 6800 1007 6866 1041
rect 6800 973 6816 1007
rect 6850 973 6866 1007
rect 6800 939 6866 973
rect 6800 905 6816 939
rect 6850 905 6866 939
rect 6800 871 6866 905
rect 6800 837 6816 871
rect 6850 837 6866 871
rect 6800 803 6866 837
rect 6800 769 6816 803
rect 6850 769 6866 803
rect 6800 735 6866 769
rect 6800 701 6816 735
rect 6850 701 6866 735
rect 6800 667 6866 701
rect 6800 633 6816 667
rect 6850 633 6866 667
rect 6800 599 6866 633
rect 6800 565 6816 599
rect 6850 565 6866 599
rect 6800 531 6866 565
rect 6800 497 6816 531
rect 6850 497 6866 531
rect 6800 463 6866 497
rect 6800 429 6816 463
rect 6850 429 6866 463
rect 6800 395 6866 429
rect 6800 361 6816 395
rect 6850 361 6866 395
rect 6800 327 6866 361
rect 6800 293 6816 327
rect 6850 293 6866 327
rect 6800 252 6866 293
rect 6896 1211 6962 1252
rect 6896 1177 6912 1211
rect 6946 1177 6962 1211
rect 6896 1143 6962 1177
rect 6896 1109 6912 1143
rect 6946 1109 6962 1143
rect 6896 1075 6962 1109
rect 6896 1041 6912 1075
rect 6946 1041 6962 1075
rect 6896 1007 6962 1041
rect 6896 973 6912 1007
rect 6946 973 6962 1007
rect 6896 939 6962 973
rect 6896 905 6912 939
rect 6946 905 6962 939
rect 6896 871 6962 905
rect 6896 837 6912 871
rect 6946 837 6962 871
rect 6896 803 6962 837
rect 6896 769 6912 803
rect 6946 769 6962 803
rect 6896 735 6962 769
rect 6896 701 6912 735
rect 6946 701 6962 735
rect 6896 667 6962 701
rect 6896 633 6912 667
rect 6946 633 6962 667
rect 6896 599 6962 633
rect 6896 565 6912 599
rect 6946 565 6962 599
rect 6896 531 6962 565
rect 6896 497 6912 531
rect 6946 497 6962 531
rect 6896 463 6962 497
rect 6896 429 6912 463
rect 6946 429 6962 463
rect 6896 395 6962 429
rect 6896 361 6912 395
rect 6946 361 6962 395
rect 6896 327 6962 361
rect 6896 293 6912 327
rect 6946 293 6962 327
rect 6896 252 6962 293
rect 6992 1211 7058 1252
rect 6992 1177 7008 1211
rect 7042 1177 7058 1211
rect 6992 1143 7058 1177
rect 6992 1109 7008 1143
rect 7042 1109 7058 1143
rect 6992 1075 7058 1109
rect 6992 1041 7008 1075
rect 7042 1041 7058 1075
rect 6992 1007 7058 1041
rect 6992 973 7008 1007
rect 7042 973 7058 1007
rect 6992 939 7058 973
rect 6992 905 7008 939
rect 7042 905 7058 939
rect 6992 871 7058 905
rect 6992 837 7008 871
rect 7042 837 7058 871
rect 6992 803 7058 837
rect 6992 769 7008 803
rect 7042 769 7058 803
rect 6992 735 7058 769
rect 6992 701 7008 735
rect 7042 701 7058 735
rect 6992 667 7058 701
rect 6992 633 7008 667
rect 7042 633 7058 667
rect 6992 599 7058 633
rect 6992 565 7008 599
rect 7042 565 7058 599
rect 6992 531 7058 565
rect 6992 497 7008 531
rect 7042 497 7058 531
rect 6992 463 7058 497
rect 6992 429 7008 463
rect 7042 429 7058 463
rect 6992 395 7058 429
rect 6992 361 7008 395
rect 7042 361 7058 395
rect 6992 327 7058 361
rect 6992 293 7008 327
rect 7042 293 7058 327
rect 6992 252 7058 293
rect 7088 1211 7154 1252
rect 7088 1177 7104 1211
rect 7138 1177 7154 1211
rect 7088 1143 7154 1177
rect 7088 1109 7104 1143
rect 7138 1109 7154 1143
rect 7088 1075 7154 1109
rect 7088 1041 7104 1075
rect 7138 1041 7154 1075
rect 7088 1007 7154 1041
rect 7088 973 7104 1007
rect 7138 973 7154 1007
rect 7088 939 7154 973
rect 7088 905 7104 939
rect 7138 905 7154 939
rect 7088 871 7154 905
rect 7088 837 7104 871
rect 7138 837 7154 871
rect 7088 803 7154 837
rect 7088 769 7104 803
rect 7138 769 7154 803
rect 7088 735 7154 769
rect 7088 701 7104 735
rect 7138 701 7154 735
rect 7088 667 7154 701
rect 7088 633 7104 667
rect 7138 633 7154 667
rect 7088 599 7154 633
rect 7088 565 7104 599
rect 7138 565 7154 599
rect 7088 531 7154 565
rect 7088 497 7104 531
rect 7138 497 7154 531
rect 7088 463 7154 497
rect 7088 429 7104 463
rect 7138 429 7154 463
rect 7088 395 7154 429
rect 7088 361 7104 395
rect 7138 361 7154 395
rect 7088 327 7154 361
rect 7088 293 7104 327
rect 7138 293 7154 327
rect 7088 252 7154 293
rect 7184 1211 7250 1252
rect 7184 1177 7200 1211
rect 7234 1177 7250 1211
rect 7184 1143 7250 1177
rect 7184 1109 7200 1143
rect 7234 1109 7250 1143
rect 7184 1075 7250 1109
rect 7184 1041 7200 1075
rect 7234 1041 7250 1075
rect 7184 1007 7250 1041
rect 7184 973 7200 1007
rect 7234 973 7250 1007
rect 7184 939 7250 973
rect 7184 905 7200 939
rect 7234 905 7250 939
rect 7184 871 7250 905
rect 7184 837 7200 871
rect 7234 837 7250 871
rect 7184 803 7250 837
rect 7184 769 7200 803
rect 7234 769 7250 803
rect 7184 735 7250 769
rect 7184 701 7200 735
rect 7234 701 7250 735
rect 7184 667 7250 701
rect 7184 633 7200 667
rect 7234 633 7250 667
rect 7184 599 7250 633
rect 7184 565 7200 599
rect 7234 565 7250 599
rect 7184 531 7250 565
rect 7184 497 7200 531
rect 7234 497 7250 531
rect 7184 463 7250 497
rect 7184 429 7200 463
rect 7234 429 7250 463
rect 7184 395 7250 429
rect 7184 361 7200 395
rect 7234 361 7250 395
rect 7184 327 7250 361
rect 7184 293 7200 327
rect 7234 293 7250 327
rect 7184 252 7250 293
rect 7280 1211 7342 1252
rect 7280 1177 7296 1211
rect 7330 1177 7342 1211
rect 7280 1143 7342 1177
rect 7280 1109 7296 1143
rect 7330 1109 7342 1143
rect 7280 1075 7342 1109
rect 7280 1041 7296 1075
rect 7330 1041 7342 1075
rect 7280 1007 7342 1041
rect 7280 973 7296 1007
rect 7330 973 7342 1007
rect 7280 939 7342 973
rect 7280 905 7296 939
rect 7330 905 7342 939
rect 7280 871 7342 905
rect 7280 837 7296 871
rect 7330 837 7342 871
rect 7280 803 7342 837
rect 7280 769 7296 803
rect 7330 769 7342 803
rect 7280 735 7342 769
rect 7280 701 7296 735
rect 7330 701 7342 735
rect 7280 667 7342 701
rect 7280 633 7296 667
rect 7330 633 7342 667
rect 7280 599 7342 633
rect 7280 565 7296 599
rect 7330 565 7342 599
rect 7280 531 7342 565
rect 7280 497 7296 531
rect 7330 497 7342 531
rect 7280 463 7342 497
rect 7280 429 7296 463
rect 7330 429 7342 463
rect 7280 395 7342 429
rect 7280 361 7296 395
rect 7330 361 7342 395
rect 7280 327 7342 361
rect 7280 293 7296 327
rect 7330 293 7342 327
rect 7280 252 7342 293
rect 7900 1211 7962 1252
rect 7900 1177 7912 1211
rect 7946 1177 7962 1211
rect 7900 1143 7962 1177
rect 7900 1109 7912 1143
rect 7946 1109 7962 1143
rect 7900 1075 7962 1109
rect 7900 1041 7912 1075
rect 7946 1041 7962 1075
rect 7900 1007 7962 1041
rect 7900 973 7912 1007
rect 7946 973 7962 1007
rect 7900 939 7962 973
rect 7900 905 7912 939
rect 7946 905 7962 939
rect 7900 871 7962 905
rect 7900 837 7912 871
rect 7946 837 7962 871
rect 7900 803 7962 837
rect 7900 769 7912 803
rect 7946 769 7962 803
rect 7900 735 7962 769
rect 7900 701 7912 735
rect 7946 701 7962 735
rect 7900 667 7962 701
rect 7900 633 7912 667
rect 7946 633 7962 667
rect 7900 599 7962 633
rect 7900 565 7912 599
rect 7946 565 7962 599
rect 7900 531 7962 565
rect 7900 497 7912 531
rect 7946 497 7962 531
rect 7900 463 7962 497
rect 7900 429 7912 463
rect 7946 429 7962 463
rect 7900 395 7962 429
rect 7900 361 7912 395
rect 7946 361 7962 395
rect 7900 327 7962 361
rect 7900 293 7912 327
rect 7946 293 7962 327
rect 7900 252 7962 293
rect 7992 1211 8058 1252
rect 7992 1177 8008 1211
rect 8042 1177 8058 1211
rect 7992 1143 8058 1177
rect 7992 1109 8008 1143
rect 8042 1109 8058 1143
rect 7992 1075 8058 1109
rect 7992 1041 8008 1075
rect 8042 1041 8058 1075
rect 7992 1007 8058 1041
rect 7992 973 8008 1007
rect 8042 973 8058 1007
rect 7992 939 8058 973
rect 7992 905 8008 939
rect 8042 905 8058 939
rect 7992 871 8058 905
rect 7992 837 8008 871
rect 8042 837 8058 871
rect 7992 803 8058 837
rect 7992 769 8008 803
rect 8042 769 8058 803
rect 7992 735 8058 769
rect 7992 701 8008 735
rect 8042 701 8058 735
rect 7992 667 8058 701
rect 7992 633 8008 667
rect 8042 633 8058 667
rect 7992 599 8058 633
rect 7992 565 8008 599
rect 8042 565 8058 599
rect 7992 531 8058 565
rect 7992 497 8008 531
rect 8042 497 8058 531
rect 7992 463 8058 497
rect 7992 429 8008 463
rect 8042 429 8058 463
rect 7992 395 8058 429
rect 7992 361 8008 395
rect 8042 361 8058 395
rect 7992 327 8058 361
rect 7992 293 8008 327
rect 8042 293 8058 327
rect 7992 252 8058 293
rect 8088 1211 8154 1252
rect 8088 1177 8104 1211
rect 8138 1177 8154 1211
rect 8088 1143 8154 1177
rect 8088 1109 8104 1143
rect 8138 1109 8154 1143
rect 8088 1075 8154 1109
rect 8088 1041 8104 1075
rect 8138 1041 8154 1075
rect 8088 1007 8154 1041
rect 8088 973 8104 1007
rect 8138 973 8154 1007
rect 8088 939 8154 973
rect 8088 905 8104 939
rect 8138 905 8154 939
rect 8088 871 8154 905
rect 8088 837 8104 871
rect 8138 837 8154 871
rect 8088 803 8154 837
rect 8088 769 8104 803
rect 8138 769 8154 803
rect 8088 735 8154 769
rect 8088 701 8104 735
rect 8138 701 8154 735
rect 8088 667 8154 701
rect 8088 633 8104 667
rect 8138 633 8154 667
rect 8088 599 8154 633
rect 8088 565 8104 599
rect 8138 565 8154 599
rect 8088 531 8154 565
rect 8088 497 8104 531
rect 8138 497 8154 531
rect 8088 463 8154 497
rect 8088 429 8104 463
rect 8138 429 8154 463
rect 8088 395 8154 429
rect 8088 361 8104 395
rect 8138 361 8154 395
rect 8088 327 8154 361
rect 8088 293 8104 327
rect 8138 293 8154 327
rect 8088 252 8154 293
rect 8184 1211 8250 1252
rect 8184 1177 8200 1211
rect 8234 1177 8250 1211
rect 8184 1143 8250 1177
rect 8184 1109 8200 1143
rect 8234 1109 8250 1143
rect 8184 1075 8250 1109
rect 8184 1041 8200 1075
rect 8234 1041 8250 1075
rect 8184 1007 8250 1041
rect 8184 973 8200 1007
rect 8234 973 8250 1007
rect 8184 939 8250 973
rect 8184 905 8200 939
rect 8234 905 8250 939
rect 8184 871 8250 905
rect 8184 837 8200 871
rect 8234 837 8250 871
rect 8184 803 8250 837
rect 8184 769 8200 803
rect 8234 769 8250 803
rect 8184 735 8250 769
rect 8184 701 8200 735
rect 8234 701 8250 735
rect 8184 667 8250 701
rect 8184 633 8200 667
rect 8234 633 8250 667
rect 8184 599 8250 633
rect 8184 565 8200 599
rect 8234 565 8250 599
rect 8184 531 8250 565
rect 8184 497 8200 531
rect 8234 497 8250 531
rect 8184 463 8250 497
rect 8184 429 8200 463
rect 8234 429 8250 463
rect 8184 395 8250 429
rect 8184 361 8200 395
rect 8234 361 8250 395
rect 8184 327 8250 361
rect 8184 293 8200 327
rect 8234 293 8250 327
rect 8184 252 8250 293
rect 8280 1211 8346 1252
rect 8280 1177 8296 1211
rect 8330 1177 8346 1211
rect 8280 1143 8346 1177
rect 8280 1109 8296 1143
rect 8330 1109 8346 1143
rect 8280 1075 8346 1109
rect 8280 1041 8296 1075
rect 8330 1041 8346 1075
rect 8280 1007 8346 1041
rect 8280 973 8296 1007
rect 8330 973 8346 1007
rect 8280 939 8346 973
rect 8280 905 8296 939
rect 8330 905 8346 939
rect 8280 871 8346 905
rect 8280 837 8296 871
rect 8330 837 8346 871
rect 8280 803 8346 837
rect 8280 769 8296 803
rect 8330 769 8346 803
rect 8280 735 8346 769
rect 8280 701 8296 735
rect 8330 701 8346 735
rect 8280 667 8346 701
rect 8280 633 8296 667
rect 8330 633 8346 667
rect 8280 599 8346 633
rect 8280 565 8296 599
rect 8330 565 8346 599
rect 8280 531 8346 565
rect 8280 497 8296 531
rect 8330 497 8346 531
rect 8280 463 8346 497
rect 8280 429 8296 463
rect 8330 429 8346 463
rect 8280 395 8346 429
rect 8280 361 8296 395
rect 8330 361 8346 395
rect 8280 327 8346 361
rect 8280 293 8296 327
rect 8330 293 8346 327
rect 8280 252 8346 293
rect 8376 1211 8442 1252
rect 8376 1177 8392 1211
rect 8426 1177 8442 1211
rect 8376 1143 8442 1177
rect 8376 1109 8392 1143
rect 8426 1109 8442 1143
rect 8376 1075 8442 1109
rect 8376 1041 8392 1075
rect 8426 1041 8442 1075
rect 8376 1007 8442 1041
rect 8376 973 8392 1007
rect 8426 973 8442 1007
rect 8376 939 8442 973
rect 8376 905 8392 939
rect 8426 905 8442 939
rect 8376 871 8442 905
rect 8376 837 8392 871
rect 8426 837 8442 871
rect 8376 803 8442 837
rect 8376 769 8392 803
rect 8426 769 8442 803
rect 8376 735 8442 769
rect 8376 701 8392 735
rect 8426 701 8442 735
rect 8376 667 8442 701
rect 8376 633 8392 667
rect 8426 633 8442 667
rect 8376 599 8442 633
rect 8376 565 8392 599
rect 8426 565 8442 599
rect 8376 531 8442 565
rect 8376 497 8392 531
rect 8426 497 8442 531
rect 8376 463 8442 497
rect 8376 429 8392 463
rect 8426 429 8442 463
rect 8376 395 8442 429
rect 8376 361 8392 395
rect 8426 361 8442 395
rect 8376 327 8442 361
rect 8376 293 8392 327
rect 8426 293 8442 327
rect 8376 252 8442 293
rect 8472 1211 8538 1252
rect 8472 1177 8488 1211
rect 8522 1177 8538 1211
rect 8472 1143 8538 1177
rect 8472 1109 8488 1143
rect 8522 1109 8538 1143
rect 8472 1075 8538 1109
rect 8472 1041 8488 1075
rect 8522 1041 8538 1075
rect 8472 1007 8538 1041
rect 8472 973 8488 1007
rect 8522 973 8538 1007
rect 8472 939 8538 973
rect 8472 905 8488 939
rect 8522 905 8538 939
rect 8472 871 8538 905
rect 8472 837 8488 871
rect 8522 837 8538 871
rect 8472 803 8538 837
rect 8472 769 8488 803
rect 8522 769 8538 803
rect 8472 735 8538 769
rect 8472 701 8488 735
rect 8522 701 8538 735
rect 8472 667 8538 701
rect 8472 633 8488 667
rect 8522 633 8538 667
rect 8472 599 8538 633
rect 8472 565 8488 599
rect 8522 565 8538 599
rect 8472 531 8538 565
rect 8472 497 8488 531
rect 8522 497 8538 531
rect 8472 463 8538 497
rect 8472 429 8488 463
rect 8522 429 8538 463
rect 8472 395 8538 429
rect 8472 361 8488 395
rect 8522 361 8538 395
rect 8472 327 8538 361
rect 8472 293 8488 327
rect 8522 293 8538 327
rect 8472 252 8538 293
rect 8568 1211 8634 1252
rect 8568 1177 8584 1211
rect 8618 1177 8634 1211
rect 8568 1143 8634 1177
rect 8568 1109 8584 1143
rect 8618 1109 8634 1143
rect 8568 1075 8634 1109
rect 8568 1041 8584 1075
rect 8618 1041 8634 1075
rect 8568 1007 8634 1041
rect 8568 973 8584 1007
rect 8618 973 8634 1007
rect 8568 939 8634 973
rect 8568 905 8584 939
rect 8618 905 8634 939
rect 8568 871 8634 905
rect 8568 837 8584 871
rect 8618 837 8634 871
rect 8568 803 8634 837
rect 8568 769 8584 803
rect 8618 769 8634 803
rect 8568 735 8634 769
rect 8568 701 8584 735
rect 8618 701 8634 735
rect 8568 667 8634 701
rect 8568 633 8584 667
rect 8618 633 8634 667
rect 8568 599 8634 633
rect 8568 565 8584 599
rect 8618 565 8634 599
rect 8568 531 8634 565
rect 8568 497 8584 531
rect 8618 497 8634 531
rect 8568 463 8634 497
rect 8568 429 8584 463
rect 8618 429 8634 463
rect 8568 395 8634 429
rect 8568 361 8584 395
rect 8618 361 8634 395
rect 8568 327 8634 361
rect 8568 293 8584 327
rect 8618 293 8634 327
rect 8568 252 8634 293
rect 8664 1211 8730 1252
rect 8664 1177 8680 1211
rect 8714 1177 8730 1211
rect 8664 1143 8730 1177
rect 8664 1109 8680 1143
rect 8714 1109 8730 1143
rect 8664 1075 8730 1109
rect 8664 1041 8680 1075
rect 8714 1041 8730 1075
rect 8664 1007 8730 1041
rect 8664 973 8680 1007
rect 8714 973 8730 1007
rect 8664 939 8730 973
rect 8664 905 8680 939
rect 8714 905 8730 939
rect 8664 871 8730 905
rect 8664 837 8680 871
rect 8714 837 8730 871
rect 8664 803 8730 837
rect 8664 769 8680 803
rect 8714 769 8730 803
rect 8664 735 8730 769
rect 8664 701 8680 735
rect 8714 701 8730 735
rect 8664 667 8730 701
rect 8664 633 8680 667
rect 8714 633 8730 667
rect 8664 599 8730 633
rect 8664 565 8680 599
rect 8714 565 8730 599
rect 8664 531 8730 565
rect 8664 497 8680 531
rect 8714 497 8730 531
rect 8664 463 8730 497
rect 8664 429 8680 463
rect 8714 429 8730 463
rect 8664 395 8730 429
rect 8664 361 8680 395
rect 8714 361 8730 395
rect 8664 327 8730 361
rect 8664 293 8680 327
rect 8714 293 8730 327
rect 8664 252 8730 293
rect 8760 1211 8826 1252
rect 8760 1177 8776 1211
rect 8810 1177 8826 1211
rect 8760 1143 8826 1177
rect 8760 1109 8776 1143
rect 8810 1109 8826 1143
rect 8760 1075 8826 1109
rect 8760 1041 8776 1075
rect 8810 1041 8826 1075
rect 8760 1007 8826 1041
rect 8760 973 8776 1007
rect 8810 973 8826 1007
rect 8760 939 8826 973
rect 8760 905 8776 939
rect 8810 905 8826 939
rect 8760 871 8826 905
rect 8760 837 8776 871
rect 8810 837 8826 871
rect 8760 803 8826 837
rect 8760 769 8776 803
rect 8810 769 8826 803
rect 8760 735 8826 769
rect 8760 701 8776 735
rect 8810 701 8826 735
rect 8760 667 8826 701
rect 8760 633 8776 667
rect 8810 633 8826 667
rect 8760 599 8826 633
rect 8760 565 8776 599
rect 8810 565 8826 599
rect 8760 531 8826 565
rect 8760 497 8776 531
rect 8810 497 8826 531
rect 8760 463 8826 497
rect 8760 429 8776 463
rect 8810 429 8826 463
rect 8760 395 8826 429
rect 8760 361 8776 395
rect 8810 361 8826 395
rect 8760 327 8826 361
rect 8760 293 8776 327
rect 8810 293 8826 327
rect 8760 252 8826 293
rect 8856 1211 8922 1252
rect 8856 1177 8872 1211
rect 8906 1177 8922 1211
rect 8856 1143 8922 1177
rect 8856 1109 8872 1143
rect 8906 1109 8922 1143
rect 8856 1075 8922 1109
rect 8856 1041 8872 1075
rect 8906 1041 8922 1075
rect 8856 1007 8922 1041
rect 8856 973 8872 1007
rect 8906 973 8922 1007
rect 8856 939 8922 973
rect 8856 905 8872 939
rect 8906 905 8922 939
rect 8856 871 8922 905
rect 8856 837 8872 871
rect 8906 837 8922 871
rect 8856 803 8922 837
rect 8856 769 8872 803
rect 8906 769 8922 803
rect 8856 735 8922 769
rect 8856 701 8872 735
rect 8906 701 8922 735
rect 8856 667 8922 701
rect 8856 633 8872 667
rect 8906 633 8922 667
rect 8856 599 8922 633
rect 8856 565 8872 599
rect 8906 565 8922 599
rect 8856 531 8922 565
rect 8856 497 8872 531
rect 8906 497 8922 531
rect 8856 463 8922 497
rect 8856 429 8872 463
rect 8906 429 8922 463
rect 8856 395 8922 429
rect 8856 361 8872 395
rect 8906 361 8922 395
rect 8856 327 8922 361
rect 8856 293 8872 327
rect 8906 293 8922 327
rect 8856 252 8922 293
rect 8952 1211 9014 1252
rect 8952 1177 8968 1211
rect 9002 1177 9014 1211
rect 8952 1143 9014 1177
rect 8952 1109 8968 1143
rect 9002 1109 9014 1143
rect 8952 1075 9014 1109
rect 8952 1041 8968 1075
rect 9002 1041 9014 1075
rect 8952 1007 9014 1041
rect 8952 973 8968 1007
rect 9002 973 9014 1007
rect 8952 939 9014 973
rect 8952 905 8968 939
rect 9002 905 9014 939
rect 8952 871 9014 905
rect 8952 837 8968 871
rect 9002 837 9014 871
rect 8952 803 9014 837
rect 8952 769 8968 803
rect 9002 769 9014 803
rect 8952 735 9014 769
rect 8952 701 8968 735
rect 9002 701 9014 735
rect 8952 667 9014 701
rect 8952 633 8968 667
rect 9002 633 9014 667
rect 8952 599 9014 633
rect 8952 565 8968 599
rect 9002 565 9014 599
rect 8952 531 9014 565
rect 8952 497 8968 531
rect 9002 497 9014 531
rect 8952 463 9014 497
rect 8952 429 8968 463
rect 9002 429 9014 463
rect 8952 395 9014 429
rect 8952 361 8968 395
rect 9002 361 9014 395
rect 8952 327 9014 361
rect 8952 293 8968 327
rect 9002 293 9014 327
rect 8952 252 9014 293
rect 9220 1209 9282 1250
rect 9220 1175 9232 1209
rect 9266 1175 9282 1209
rect 9220 1141 9282 1175
rect 9220 1107 9232 1141
rect 9266 1107 9282 1141
rect 9220 1073 9282 1107
rect 9220 1039 9232 1073
rect 9266 1039 9282 1073
rect 9220 1005 9282 1039
rect 9220 971 9232 1005
rect 9266 971 9282 1005
rect 9220 937 9282 971
rect 9220 903 9232 937
rect 9266 903 9282 937
rect 9220 869 9282 903
rect 9220 835 9232 869
rect 9266 835 9282 869
rect 9220 801 9282 835
rect 9220 767 9232 801
rect 9266 767 9282 801
rect 9220 733 9282 767
rect 9220 699 9232 733
rect 9266 699 9282 733
rect 9220 665 9282 699
rect 9220 631 9232 665
rect 9266 631 9282 665
rect 9220 597 9282 631
rect 9220 563 9232 597
rect 9266 563 9282 597
rect 9220 529 9282 563
rect 9220 495 9232 529
rect 9266 495 9282 529
rect 9220 461 9282 495
rect 9220 427 9232 461
rect 9266 427 9282 461
rect 9220 393 9282 427
rect 9220 359 9232 393
rect 9266 359 9282 393
rect 9220 325 9282 359
rect 9220 291 9232 325
rect 9266 291 9282 325
rect -914 107 -902 141
rect -868 107 -856 141
rect -914 66 -856 107
rect 9220 250 9282 291
rect 9312 1209 9378 1250
rect 9312 1175 9328 1209
rect 9362 1175 9378 1209
rect 9312 1141 9378 1175
rect 9312 1107 9328 1141
rect 9362 1107 9378 1141
rect 9312 1073 9378 1107
rect 9312 1039 9328 1073
rect 9362 1039 9378 1073
rect 9312 1005 9378 1039
rect 9312 971 9328 1005
rect 9362 971 9378 1005
rect 9312 937 9378 971
rect 9312 903 9328 937
rect 9362 903 9378 937
rect 9312 869 9378 903
rect 9312 835 9328 869
rect 9362 835 9378 869
rect 9312 801 9378 835
rect 9312 767 9328 801
rect 9362 767 9378 801
rect 9312 733 9378 767
rect 9312 699 9328 733
rect 9362 699 9378 733
rect 9312 665 9378 699
rect 9312 631 9328 665
rect 9362 631 9378 665
rect 9312 597 9378 631
rect 9312 563 9328 597
rect 9362 563 9378 597
rect 9312 529 9378 563
rect 9312 495 9328 529
rect 9362 495 9378 529
rect 9312 461 9378 495
rect 9312 427 9328 461
rect 9362 427 9378 461
rect 9312 393 9378 427
rect 9312 359 9328 393
rect 9362 359 9378 393
rect 9312 325 9378 359
rect 9312 291 9328 325
rect 9362 291 9378 325
rect 9312 250 9378 291
rect 9408 1209 9474 1250
rect 9408 1175 9424 1209
rect 9458 1175 9474 1209
rect 9408 1141 9474 1175
rect 9408 1107 9424 1141
rect 9458 1107 9474 1141
rect 9408 1073 9474 1107
rect 9408 1039 9424 1073
rect 9458 1039 9474 1073
rect 9408 1005 9474 1039
rect 9408 971 9424 1005
rect 9458 971 9474 1005
rect 9408 937 9474 971
rect 9408 903 9424 937
rect 9458 903 9474 937
rect 9408 869 9474 903
rect 9408 835 9424 869
rect 9458 835 9474 869
rect 9408 801 9474 835
rect 9408 767 9424 801
rect 9458 767 9474 801
rect 9408 733 9474 767
rect 9408 699 9424 733
rect 9458 699 9474 733
rect 9408 665 9474 699
rect 9408 631 9424 665
rect 9458 631 9474 665
rect 9408 597 9474 631
rect 9408 563 9424 597
rect 9458 563 9474 597
rect 9408 529 9474 563
rect 9408 495 9424 529
rect 9458 495 9474 529
rect 9408 461 9474 495
rect 9408 427 9424 461
rect 9458 427 9474 461
rect 9408 393 9474 427
rect 9408 359 9424 393
rect 9458 359 9474 393
rect 9408 325 9474 359
rect 9408 291 9424 325
rect 9458 291 9474 325
rect 9408 250 9474 291
rect 9504 1209 9570 1250
rect 9504 1175 9520 1209
rect 9554 1175 9570 1209
rect 9504 1141 9570 1175
rect 9504 1107 9520 1141
rect 9554 1107 9570 1141
rect 9504 1073 9570 1107
rect 9504 1039 9520 1073
rect 9554 1039 9570 1073
rect 9504 1005 9570 1039
rect 9504 971 9520 1005
rect 9554 971 9570 1005
rect 9504 937 9570 971
rect 9504 903 9520 937
rect 9554 903 9570 937
rect 9504 869 9570 903
rect 9504 835 9520 869
rect 9554 835 9570 869
rect 9504 801 9570 835
rect 9504 767 9520 801
rect 9554 767 9570 801
rect 9504 733 9570 767
rect 9504 699 9520 733
rect 9554 699 9570 733
rect 9504 665 9570 699
rect 9504 631 9520 665
rect 9554 631 9570 665
rect 9504 597 9570 631
rect 9504 563 9520 597
rect 9554 563 9570 597
rect 9504 529 9570 563
rect 9504 495 9520 529
rect 9554 495 9570 529
rect 9504 461 9570 495
rect 9504 427 9520 461
rect 9554 427 9570 461
rect 9504 393 9570 427
rect 9504 359 9520 393
rect 9554 359 9570 393
rect 9504 325 9570 359
rect 9504 291 9520 325
rect 9554 291 9570 325
rect 9504 250 9570 291
rect 9600 1209 9666 1250
rect 9600 1175 9616 1209
rect 9650 1175 9666 1209
rect 9600 1141 9666 1175
rect 9600 1107 9616 1141
rect 9650 1107 9666 1141
rect 9600 1073 9666 1107
rect 9600 1039 9616 1073
rect 9650 1039 9666 1073
rect 9600 1005 9666 1039
rect 9600 971 9616 1005
rect 9650 971 9666 1005
rect 9600 937 9666 971
rect 9600 903 9616 937
rect 9650 903 9666 937
rect 9600 869 9666 903
rect 9600 835 9616 869
rect 9650 835 9666 869
rect 9600 801 9666 835
rect 9600 767 9616 801
rect 9650 767 9666 801
rect 9600 733 9666 767
rect 9600 699 9616 733
rect 9650 699 9666 733
rect 9600 665 9666 699
rect 9600 631 9616 665
rect 9650 631 9666 665
rect 9600 597 9666 631
rect 9600 563 9616 597
rect 9650 563 9666 597
rect 9600 529 9666 563
rect 9600 495 9616 529
rect 9650 495 9666 529
rect 9600 461 9666 495
rect 9600 427 9616 461
rect 9650 427 9666 461
rect 9600 393 9666 427
rect 9600 359 9616 393
rect 9650 359 9666 393
rect 9600 325 9666 359
rect 9600 291 9616 325
rect 9650 291 9666 325
rect 9600 250 9666 291
rect 9696 1209 9762 1250
rect 9696 1175 9712 1209
rect 9746 1175 9762 1209
rect 9696 1141 9762 1175
rect 9696 1107 9712 1141
rect 9746 1107 9762 1141
rect 9696 1073 9762 1107
rect 9696 1039 9712 1073
rect 9746 1039 9762 1073
rect 9696 1005 9762 1039
rect 9696 971 9712 1005
rect 9746 971 9762 1005
rect 9696 937 9762 971
rect 9696 903 9712 937
rect 9746 903 9762 937
rect 9696 869 9762 903
rect 9696 835 9712 869
rect 9746 835 9762 869
rect 9696 801 9762 835
rect 9696 767 9712 801
rect 9746 767 9762 801
rect 9696 733 9762 767
rect 9696 699 9712 733
rect 9746 699 9762 733
rect 9696 665 9762 699
rect 9696 631 9712 665
rect 9746 631 9762 665
rect 9696 597 9762 631
rect 9696 563 9712 597
rect 9746 563 9762 597
rect 9696 529 9762 563
rect 9696 495 9712 529
rect 9746 495 9762 529
rect 9696 461 9762 495
rect 9696 427 9712 461
rect 9746 427 9762 461
rect 9696 393 9762 427
rect 9696 359 9712 393
rect 9746 359 9762 393
rect 9696 325 9762 359
rect 9696 291 9712 325
rect 9746 291 9762 325
rect 9696 250 9762 291
rect 9792 1209 9858 1250
rect 9792 1175 9808 1209
rect 9842 1175 9858 1209
rect 9792 1141 9858 1175
rect 9792 1107 9808 1141
rect 9842 1107 9858 1141
rect 9792 1073 9858 1107
rect 9792 1039 9808 1073
rect 9842 1039 9858 1073
rect 9792 1005 9858 1039
rect 9792 971 9808 1005
rect 9842 971 9858 1005
rect 9792 937 9858 971
rect 9792 903 9808 937
rect 9842 903 9858 937
rect 9792 869 9858 903
rect 9792 835 9808 869
rect 9842 835 9858 869
rect 9792 801 9858 835
rect 9792 767 9808 801
rect 9842 767 9858 801
rect 9792 733 9858 767
rect 9792 699 9808 733
rect 9842 699 9858 733
rect 9792 665 9858 699
rect 9792 631 9808 665
rect 9842 631 9858 665
rect 9792 597 9858 631
rect 9792 563 9808 597
rect 9842 563 9858 597
rect 9792 529 9858 563
rect 9792 495 9808 529
rect 9842 495 9858 529
rect 9792 461 9858 495
rect 9792 427 9808 461
rect 9842 427 9858 461
rect 9792 393 9858 427
rect 9792 359 9808 393
rect 9842 359 9858 393
rect 9792 325 9858 359
rect 9792 291 9808 325
rect 9842 291 9858 325
rect 9792 250 9858 291
rect 9888 1209 9954 1250
rect 9888 1175 9904 1209
rect 9938 1175 9954 1209
rect 9888 1141 9954 1175
rect 9888 1107 9904 1141
rect 9938 1107 9954 1141
rect 9888 1073 9954 1107
rect 9888 1039 9904 1073
rect 9938 1039 9954 1073
rect 9888 1005 9954 1039
rect 9888 971 9904 1005
rect 9938 971 9954 1005
rect 9888 937 9954 971
rect 9888 903 9904 937
rect 9938 903 9954 937
rect 9888 869 9954 903
rect 9888 835 9904 869
rect 9938 835 9954 869
rect 9888 801 9954 835
rect 9888 767 9904 801
rect 9938 767 9954 801
rect 9888 733 9954 767
rect 9888 699 9904 733
rect 9938 699 9954 733
rect 9888 665 9954 699
rect 9888 631 9904 665
rect 9938 631 9954 665
rect 9888 597 9954 631
rect 9888 563 9904 597
rect 9938 563 9954 597
rect 9888 529 9954 563
rect 9888 495 9904 529
rect 9938 495 9954 529
rect 9888 461 9954 495
rect 9888 427 9904 461
rect 9938 427 9954 461
rect 9888 393 9954 427
rect 9888 359 9904 393
rect 9938 359 9954 393
rect 9888 325 9954 359
rect 9888 291 9904 325
rect 9938 291 9954 325
rect 9888 250 9954 291
rect 9984 1209 10050 1250
rect 9984 1175 10000 1209
rect 10034 1175 10050 1209
rect 9984 1141 10050 1175
rect 9984 1107 10000 1141
rect 10034 1107 10050 1141
rect 9984 1073 10050 1107
rect 9984 1039 10000 1073
rect 10034 1039 10050 1073
rect 9984 1005 10050 1039
rect 9984 971 10000 1005
rect 10034 971 10050 1005
rect 9984 937 10050 971
rect 9984 903 10000 937
rect 10034 903 10050 937
rect 9984 869 10050 903
rect 9984 835 10000 869
rect 10034 835 10050 869
rect 9984 801 10050 835
rect 9984 767 10000 801
rect 10034 767 10050 801
rect 9984 733 10050 767
rect 9984 699 10000 733
rect 10034 699 10050 733
rect 9984 665 10050 699
rect 9984 631 10000 665
rect 10034 631 10050 665
rect 9984 597 10050 631
rect 9984 563 10000 597
rect 10034 563 10050 597
rect 9984 529 10050 563
rect 9984 495 10000 529
rect 10034 495 10050 529
rect 9984 461 10050 495
rect 9984 427 10000 461
rect 10034 427 10050 461
rect 9984 393 10050 427
rect 9984 359 10000 393
rect 10034 359 10050 393
rect 9984 325 10050 359
rect 9984 291 10000 325
rect 10034 291 10050 325
rect 9984 250 10050 291
rect 10080 1209 10146 1250
rect 10080 1175 10096 1209
rect 10130 1175 10146 1209
rect 10080 1141 10146 1175
rect 10080 1107 10096 1141
rect 10130 1107 10146 1141
rect 10080 1073 10146 1107
rect 10080 1039 10096 1073
rect 10130 1039 10146 1073
rect 10080 1005 10146 1039
rect 10080 971 10096 1005
rect 10130 971 10146 1005
rect 10080 937 10146 971
rect 10080 903 10096 937
rect 10130 903 10146 937
rect 10080 869 10146 903
rect 10080 835 10096 869
rect 10130 835 10146 869
rect 10080 801 10146 835
rect 10080 767 10096 801
rect 10130 767 10146 801
rect 10080 733 10146 767
rect 10080 699 10096 733
rect 10130 699 10146 733
rect 10080 665 10146 699
rect 10080 631 10096 665
rect 10130 631 10146 665
rect 10080 597 10146 631
rect 10080 563 10096 597
rect 10130 563 10146 597
rect 10080 529 10146 563
rect 10080 495 10096 529
rect 10130 495 10146 529
rect 10080 461 10146 495
rect 10080 427 10096 461
rect 10130 427 10146 461
rect 10080 393 10146 427
rect 10080 359 10096 393
rect 10130 359 10146 393
rect 10080 325 10146 359
rect 10080 291 10096 325
rect 10130 291 10146 325
rect 10080 250 10146 291
rect 10176 1209 10242 1250
rect 10176 1175 10192 1209
rect 10226 1175 10242 1209
rect 10176 1141 10242 1175
rect 10176 1107 10192 1141
rect 10226 1107 10242 1141
rect 10176 1073 10242 1107
rect 10176 1039 10192 1073
rect 10226 1039 10242 1073
rect 10176 1005 10242 1039
rect 10176 971 10192 1005
rect 10226 971 10242 1005
rect 10176 937 10242 971
rect 10176 903 10192 937
rect 10226 903 10242 937
rect 10176 869 10242 903
rect 10176 835 10192 869
rect 10226 835 10242 869
rect 10176 801 10242 835
rect 10176 767 10192 801
rect 10226 767 10242 801
rect 10176 733 10242 767
rect 10176 699 10192 733
rect 10226 699 10242 733
rect 10176 665 10242 699
rect 10176 631 10192 665
rect 10226 631 10242 665
rect 10176 597 10242 631
rect 10176 563 10192 597
rect 10226 563 10242 597
rect 10176 529 10242 563
rect 10176 495 10192 529
rect 10226 495 10242 529
rect 10176 461 10242 495
rect 10176 427 10192 461
rect 10226 427 10242 461
rect 10176 393 10242 427
rect 10176 359 10192 393
rect 10226 359 10242 393
rect 10176 325 10242 359
rect 10176 291 10192 325
rect 10226 291 10242 325
rect 10176 250 10242 291
rect 10272 1209 10338 1250
rect 10272 1175 10288 1209
rect 10322 1175 10338 1209
rect 10272 1141 10338 1175
rect 10272 1107 10288 1141
rect 10322 1107 10338 1141
rect 10272 1073 10338 1107
rect 10272 1039 10288 1073
rect 10322 1039 10338 1073
rect 10272 1005 10338 1039
rect 10272 971 10288 1005
rect 10322 971 10338 1005
rect 10272 937 10338 971
rect 10272 903 10288 937
rect 10322 903 10338 937
rect 10272 869 10338 903
rect 10272 835 10288 869
rect 10322 835 10338 869
rect 10272 801 10338 835
rect 10272 767 10288 801
rect 10322 767 10338 801
rect 10272 733 10338 767
rect 10272 699 10288 733
rect 10322 699 10338 733
rect 10272 665 10338 699
rect 10272 631 10288 665
rect 10322 631 10338 665
rect 10272 597 10338 631
rect 10272 563 10288 597
rect 10322 563 10338 597
rect 10272 529 10338 563
rect 10272 495 10288 529
rect 10322 495 10338 529
rect 10272 461 10338 495
rect 10272 427 10288 461
rect 10322 427 10338 461
rect 10272 393 10338 427
rect 10272 359 10288 393
rect 10322 359 10338 393
rect 10272 325 10338 359
rect 10272 291 10288 325
rect 10322 291 10338 325
rect 10272 250 10338 291
rect 10368 1209 10430 1250
rect 10368 1175 10384 1209
rect 10418 1175 10430 1209
rect 10368 1141 10430 1175
rect 10368 1107 10384 1141
rect 10418 1107 10430 1141
rect 10368 1073 10430 1107
rect 10368 1039 10384 1073
rect 10418 1039 10430 1073
rect 10368 1005 10430 1039
rect 10368 971 10384 1005
rect 10418 971 10430 1005
rect 10368 937 10430 971
rect 10368 903 10384 937
rect 10418 903 10430 937
rect 10368 869 10430 903
rect 10368 835 10384 869
rect 10418 835 10430 869
rect 10368 801 10430 835
rect 10368 767 10384 801
rect 10418 767 10430 801
rect 10368 733 10430 767
rect 10368 699 10384 733
rect 10418 699 10430 733
rect 10368 665 10430 699
rect 10368 631 10384 665
rect 10418 631 10430 665
rect 10368 597 10430 631
rect 10368 563 10384 597
rect 10418 563 10430 597
rect 10368 529 10430 563
rect 10368 495 10384 529
rect 10418 495 10430 529
rect 10368 461 10430 495
rect 10368 427 10384 461
rect 10418 427 10430 461
rect 10368 393 10430 427
rect 10368 359 10384 393
rect 10418 359 10430 393
rect 10368 325 10430 359
rect 10368 291 10384 325
rect 10418 291 10430 325
rect 10368 250 10430 291
rect 10988 1209 11050 1250
rect 10988 1175 11000 1209
rect 11034 1175 11050 1209
rect 10988 1141 11050 1175
rect 10988 1107 11000 1141
rect 11034 1107 11050 1141
rect 10988 1073 11050 1107
rect 10988 1039 11000 1073
rect 11034 1039 11050 1073
rect 10988 1005 11050 1039
rect 10988 971 11000 1005
rect 11034 971 11050 1005
rect 10988 937 11050 971
rect 10988 903 11000 937
rect 11034 903 11050 937
rect 10988 869 11050 903
rect 10988 835 11000 869
rect 11034 835 11050 869
rect 10988 801 11050 835
rect 10988 767 11000 801
rect 11034 767 11050 801
rect 10988 733 11050 767
rect 10988 699 11000 733
rect 11034 699 11050 733
rect 10988 665 11050 699
rect 10988 631 11000 665
rect 11034 631 11050 665
rect 10988 597 11050 631
rect 10988 563 11000 597
rect 11034 563 11050 597
rect 10988 529 11050 563
rect 10988 495 11000 529
rect 11034 495 11050 529
rect 10988 461 11050 495
rect 10988 427 11000 461
rect 11034 427 11050 461
rect 10988 393 11050 427
rect 10988 359 11000 393
rect 11034 359 11050 393
rect 10988 325 11050 359
rect 10988 291 11000 325
rect 11034 291 11050 325
rect 10988 250 11050 291
rect 11080 1209 11146 1250
rect 11080 1175 11096 1209
rect 11130 1175 11146 1209
rect 11080 1141 11146 1175
rect 11080 1107 11096 1141
rect 11130 1107 11146 1141
rect 11080 1073 11146 1107
rect 11080 1039 11096 1073
rect 11130 1039 11146 1073
rect 11080 1005 11146 1039
rect 11080 971 11096 1005
rect 11130 971 11146 1005
rect 11080 937 11146 971
rect 11080 903 11096 937
rect 11130 903 11146 937
rect 11080 869 11146 903
rect 11080 835 11096 869
rect 11130 835 11146 869
rect 11080 801 11146 835
rect 11080 767 11096 801
rect 11130 767 11146 801
rect 11080 733 11146 767
rect 11080 699 11096 733
rect 11130 699 11146 733
rect 11080 665 11146 699
rect 11080 631 11096 665
rect 11130 631 11146 665
rect 11080 597 11146 631
rect 11080 563 11096 597
rect 11130 563 11146 597
rect 11080 529 11146 563
rect 11080 495 11096 529
rect 11130 495 11146 529
rect 11080 461 11146 495
rect 11080 427 11096 461
rect 11130 427 11146 461
rect 11080 393 11146 427
rect 11080 359 11096 393
rect 11130 359 11146 393
rect 11080 325 11146 359
rect 11080 291 11096 325
rect 11130 291 11146 325
rect 11080 250 11146 291
rect 11176 1209 11242 1250
rect 11176 1175 11192 1209
rect 11226 1175 11242 1209
rect 11176 1141 11242 1175
rect 11176 1107 11192 1141
rect 11226 1107 11242 1141
rect 11176 1073 11242 1107
rect 11176 1039 11192 1073
rect 11226 1039 11242 1073
rect 11176 1005 11242 1039
rect 11176 971 11192 1005
rect 11226 971 11242 1005
rect 11176 937 11242 971
rect 11176 903 11192 937
rect 11226 903 11242 937
rect 11176 869 11242 903
rect 11176 835 11192 869
rect 11226 835 11242 869
rect 11176 801 11242 835
rect 11176 767 11192 801
rect 11226 767 11242 801
rect 11176 733 11242 767
rect 11176 699 11192 733
rect 11226 699 11242 733
rect 11176 665 11242 699
rect 11176 631 11192 665
rect 11226 631 11242 665
rect 11176 597 11242 631
rect 11176 563 11192 597
rect 11226 563 11242 597
rect 11176 529 11242 563
rect 11176 495 11192 529
rect 11226 495 11242 529
rect 11176 461 11242 495
rect 11176 427 11192 461
rect 11226 427 11242 461
rect 11176 393 11242 427
rect 11176 359 11192 393
rect 11226 359 11242 393
rect 11176 325 11242 359
rect 11176 291 11192 325
rect 11226 291 11242 325
rect 11176 250 11242 291
rect 11272 1209 11338 1250
rect 11272 1175 11288 1209
rect 11322 1175 11338 1209
rect 11272 1141 11338 1175
rect 11272 1107 11288 1141
rect 11322 1107 11338 1141
rect 11272 1073 11338 1107
rect 11272 1039 11288 1073
rect 11322 1039 11338 1073
rect 11272 1005 11338 1039
rect 11272 971 11288 1005
rect 11322 971 11338 1005
rect 11272 937 11338 971
rect 11272 903 11288 937
rect 11322 903 11338 937
rect 11272 869 11338 903
rect 11272 835 11288 869
rect 11322 835 11338 869
rect 11272 801 11338 835
rect 11272 767 11288 801
rect 11322 767 11338 801
rect 11272 733 11338 767
rect 11272 699 11288 733
rect 11322 699 11338 733
rect 11272 665 11338 699
rect 11272 631 11288 665
rect 11322 631 11338 665
rect 11272 597 11338 631
rect 11272 563 11288 597
rect 11322 563 11338 597
rect 11272 529 11338 563
rect 11272 495 11288 529
rect 11322 495 11338 529
rect 11272 461 11338 495
rect 11272 427 11288 461
rect 11322 427 11338 461
rect 11272 393 11338 427
rect 11272 359 11288 393
rect 11322 359 11338 393
rect 11272 325 11338 359
rect 11272 291 11288 325
rect 11322 291 11338 325
rect 11272 250 11338 291
rect 11368 1209 11434 1250
rect 11368 1175 11384 1209
rect 11418 1175 11434 1209
rect 11368 1141 11434 1175
rect 11368 1107 11384 1141
rect 11418 1107 11434 1141
rect 11368 1073 11434 1107
rect 11368 1039 11384 1073
rect 11418 1039 11434 1073
rect 11368 1005 11434 1039
rect 11368 971 11384 1005
rect 11418 971 11434 1005
rect 11368 937 11434 971
rect 11368 903 11384 937
rect 11418 903 11434 937
rect 11368 869 11434 903
rect 11368 835 11384 869
rect 11418 835 11434 869
rect 11368 801 11434 835
rect 11368 767 11384 801
rect 11418 767 11434 801
rect 11368 733 11434 767
rect 11368 699 11384 733
rect 11418 699 11434 733
rect 11368 665 11434 699
rect 11368 631 11384 665
rect 11418 631 11434 665
rect 11368 597 11434 631
rect 11368 563 11384 597
rect 11418 563 11434 597
rect 11368 529 11434 563
rect 11368 495 11384 529
rect 11418 495 11434 529
rect 11368 461 11434 495
rect 11368 427 11384 461
rect 11418 427 11434 461
rect 11368 393 11434 427
rect 11368 359 11384 393
rect 11418 359 11434 393
rect 11368 325 11434 359
rect 11368 291 11384 325
rect 11418 291 11434 325
rect 11368 250 11434 291
rect 11464 1209 11530 1250
rect 11464 1175 11480 1209
rect 11514 1175 11530 1209
rect 11464 1141 11530 1175
rect 11464 1107 11480 1141
rect 11514 1107 11530 1141
rect 11464 1073 11530 1107
rect 11464 1039 11480 1073
rect 11514 1039 11530 1073
rect 11464 1005 11530 1039
rect 11464 971 11480 1005
rect 11514 971 11530 1005
rect 11464 937 11530 971
rect 11464 903 11480 937
rect 11514 903 11530 937
rect 11464 869 11530 903
rect 11464 835 11480 869
rect 11514 835 11530 869
rect 11464 801 11530 835
rect 11464 767 11480 801
rect 11514 767 11530 801
rect 11464 733 11530 767
rect 11464 699 11480 733
rect 11514 699 11530 733
rect 11464 665 11530 699
rect 11464 631 11480 665
rect 11514 631 11530 665
rect 11464 597 11530 631
rect 11464 563 11480 597
rect 11514 563 11530 597
rect 11464 529 11530 563
rect 11464 495 11480 529
rect 11514 495 11530 529
rect 11464 461 11530 495
rect 11464 427 11480 461
rect 11514 427 11530 461
rect 11464 393 11530 427
rect 11464 359 11480 393
rect 11514 359 11530 393
rect 11464 325 11530 359
rect 11464 291 11480 325
rect 11514 291 11530 325
rect 11464 250 11530 291
rect 11560 1209 11626 1250
rect 11560 1175 11576 1209
rect 11610 1175 11626 1209
rect 11560 1141 11626 1175
rect 11560 1107 11576 1141
rect 11610 1107 11626 1141
rect 11560 1073 11626 1107
rect 11560 1039 11576 1073
rect 11610 1039 11626 1073
rect 11560 1005 11626 1039
rect 11560 971 11576 1005
rect 11610 971 11626 1005
rect 11560 937 11626 971
rect 11560 903 11576 937
rect 11610 903 11626 937
rect 11560 869 11626 903
rect 11560 835 11576 869
rect 11610 835 11626 869
rect 11560 801 11626 835
rect 11560 767 11576 801
rect 11610 767 11626 801
rect 11560 733 11626 767
rect 11560 699 11576 733
rect 11610 699 11626 733
rect 11560 665 11626 699
rect 11560 631 11576 665
rect 11610 631 11626 665
rect 11560 597 11626 631
rect 11560 563 11576 597
rect 11610 563 11626 597
rect 11560 529 11626 563
rect 11560 495 11576 529
rect 11610 495 11626 529
rect 11560 461 11626 495
rect 11560 427 11576 461
rect 11610 427 11626 461
rect 11560 393 11626 427
rect 11560 359 11576 393
rect 11610 359 11626 393
rect 11560 325 11626 359
rect 11560 291 11576 325
rect 11610 291 11626 325
rect 11560 250 11626 291
rect 11656 1209 11722 1250
rect 11656 1175 11672 1209
rect 11706 1175 11722 1209
rect 11656 1141 11722 1175
rect 11656 1107 11672 1141
rect 11706 1107 11722 1141
rect 11656 1073 11722 1107
rect 11656 1039 11672 1073
rect 11706 1039 11722 1073
rect 11656 1005 11722 1039
rect 11656 971 11672 1005
rect 11706 971 11722 1005
rect 11656 937 11722 971
rect 11656 903 11672 937
rect 11706 903 11722 937
rect 11656 869 11722 903
rect 11656 835 11672 869
rect 11706 835 11722 869
rect 11656 801 11722 835
rect 11656 767 11672 801
rect 11706 767 11722 801
rect 11656 733 11722 767
rect 11656 699 11672 733
rect 11706 699 11722 733
rect 11656 665 11722 699
rect 11656 631 11672 665
rect 11706 631 11722 665
rect 11656 597 11722 631
rect 11656 563 11672 597
rect 11706 563 11722 597
rect 11656 529 11722 563
rect 11656 495 11672 529
rect 11706 495 11722 529
rect 11656 461 11722 495
rect 11656 427 11672 461
rect 11706 427 11722 461
rect 11656 393 11722 427
rect 11656 359 11672 393
rect 11706 359 11722 393
rect 11656 325 11722 359
rect 11656 291 11672 325
rect 11706 291 11722 325
rect 11656 250 11722 291
rect 11752 1209 11818 1250
rect 11752 1175 11768 1209
rect 11802 1175 11818 1209
rect 11752 1141 11818 1175
rect 11752 1107 11768 1141
rect 11802 1107 11818 1141
rect 11752 1073 11818 1107
rect 11752 1039 11768 1073
rect 11802 1039 11818 1073
rect 11752 1005 11818 1039
rect 11752 971 11768 1005
rect 11802 971 11818 1005
rect 11752 937 11818 971
rect 11752 903 11768 937
rect 11802 903 11818 937
rect 11752 869 11818 903
rect 11752 835 11768 869
rect 11802 835 11818 869
rect 11752 801 11818 835
rect 11752 767 11768 801
rect 11802 767 11818 801
rect 11752 733 11818 767
rect 11752 699 11768 733
rect 11802 699 11818 733
rect 11752 665 11818 699
rect 11752 631 11768 665
rect 11802 631 11818 665
rect 11752 597 11818 631
rect 11752 563 11768 597
rect 11802 563 11818 597
rect 11752 529 11818 563
rect 11752 495 11768 529
rect 11802 495 11818 529
rect 11752 461 11818 495
rect 11752 427 11768 461
rect 11802 427 11818 461
rect 11752 393 11818 427
rect 11752 359 11768 393
rect 11802 359 11818 393
rect 11752 325 11818 359
rect 11752 291 11768 325
rect 11802 291 11818 325
rect 11752 250 11818 291
rect 11848 1209 11914 1250
rect 11848 1175 11864 1209
rect 11898 1175 11914 1209
rect 11848 1141 11914 1175
rect 11848 1107 11864 1141
rect 11898 1107 11914 1141
rect 11848 1073 11914 1107
rect 11848 1039 11864 1073
rect 11898 1039 11914 1073
rect 11848 1005 11914 1039
rect 11848 971 11864 1005
rect 11898 971 11914 1005
rect 11848 937 11914 971
rect 11848 903 11864 937
rect 11898 903 11914 937
rect 11848 869 11914 903
rect 11848 835 11864 869
rect 11898 835 11914 869
rect 11848 801 11914 835
rect 11848 767 11864 801
rect 11898 767 11914 801
rect 11848 733 11914 767
rect 11848 699 11864 733
rect 11898 699 11914 733
rect 11848 665 11914 699
rect 11848 631 11864 665
rect 11898 631 11914 665
rect 11848 597 11914 631
rect 11848 563 11864 597
rect 11898 563 11914 597
rect 11848 529 11914 563
rect 11848 495 11864 529
rect 11898 495 11914 529
rect 11848 461 11914 495
rect 11848 427 11864 461
rect 11898 427 11914 461
rect 11848 393 11914 427
rect 11848 359 11864 393
rect 11898 359 11914 393
rect 11848 325 11914 359
rect 11848 291 11864 325
rect 11898 291 11914 325
rect 11848 250 11914 291
rect 11944 1209 12010 1250
rect 11944 1175 11960 1209
rect 11994 1175 12010 1209
rect 11944 1141 12010 1175
rect 11944 1107 11960 1141
rect 11994 1107 12010 1141
rect 11944 1073 12010 1107
rect 11944 1039 11960 1073
rect 11994 1039 12010 1073
rect 11944 1005 12010 1039
rect 11944 971 11960 1005
rect 11994 971 12010 1005
rect 11944 937 12010 971
rect 11944 903 11960 937
rect 11994 903 12010 937
rect 11944 869 12010 903
rect 11944 835 11960 869
rect 11994 835 12010 869
rect 11944 801 12010 835
rect 11944 767 11960 801
rect 11994 767 12010 801
rect 11944 733 12010 767
rect 11944 699 11960 733
rect 11994 699 12010 733
rect 11944 665 12010 699
rect 11944 631 11960 665
rect 11994 631 12010 665
rect 11944 597 12010 631
rect 11944 563 11960 597
rect 11994 563 12010 597
rect 11944 529 12010 563
rect 11944 495 11960 529
rect 11994 495 12010 529
rect 11944 461 12010 495
rect 11944 427 11960 461
rect 11994 427 12010 461
rect 11944 393 12010 427
rect 11944 359 11960 393
rect 11994 359 12010 393
rect 11944 325 12010 359
rect 11944 291 11960 325
rect 11994 291 12010 325
rect 11944 250 12010 291
rect 12040 1209 12102 1250
rect 15410 1261 15468 1300
rect 15410 1227 15422 1261
rect 15456 1227 15468 1261
rect 12040 1175 12056 1209
rect 12090 1175 12102 1209
rect 12040 1141 12102 1175
rect 12040 1107 12056 1141
rect 12090 1107 12102 1141
rect 12040 1073 12102 1107
rect 12040 1039 12056 1073
rect 12090 1039 12102 1073
rect 12040 1005 12102 1039
rect 12040 971 12056 1005
rect 12090 971 12102 1005
rect 12040 937 12102 971
rect 12040 903 12056 937
rect 12090 903 12102 937
rect 12040 869 12102 903
rect 12040 835 12056 869
rect 12090 835 12102 869
rect 12040 801 12102 835
rect 12040 767 12056 801
rect 12090 767 12102 801
rect 12040 733 12102 767
rect 12040 699 12056 733
rect 12090 699 12102 733
rect 12040 665 12102 699
rect 12040 631 12056 665
rect 12090 631 12102 665
rect 12040 597 12102 631
rect 12040 563 12056 597
rect 12090 563 12102 597
rect 12040 529 12102 563
rect 12040 495 12056 529
rect 12090 495 12102 529
rect 12040 461 12102 495
rect 12040 427 12056 461
rect 12090 427 12102 461
rect 12040 393 12102 427
rect 12040 359 12056 393
rect 12090 359 12102 393
rect 12040 325 12102 359
rect 12040 291 12056 325
rect 12090 291 12102 325
rect 12040 250 12102 291
rect 12376 1183 12438 1224
rect 12376 1149 12388 1183
rect 12422 1149 12438 1183
rect 12376 1115 12438 1149
rect 12376 1081 12388 1115
rect 12422 1081 12438 1115
rect 12376 1047 12438 1081
rect 12376 1013 12388 1047
rect 12422 1013 12438 1047
rect 12376 979 12438 1013
rect 12376 945 12388 979
rect 12422 945 12438 979
rect 12376 911 12438 945
rect 12376 877 12388 911
rect 12422 877 12438 911
rect 12376 843 12438 877
rect 12376 809 12388 843
rect 12422 809 12438 843
rect 12376 775 12438 809
rect 12376 741 12388 775
rect 12422 741 12438 775
rect 12376 707 12438 741
rect 12376 673 12388 707
rect 12422 673 12438 707
rect 12376 639 12438 673
rect 12376 605 12388 639
rect 12422 605 12438 639
rect 12376 571 12438 605
rect 12376 537 12388 571
rect 12422 537 12438 571
rect 12376 503 12438 537
rect 12376 469 12388 503
rect 12422 469 12438 503
rect 12376 435 12438 469
rect 12376 401 12388 435
rect 12422 401 12438 435
rect 12376 367 12438 401
rect 12376 333 12388 367
rect 12422 333 12438 367
rect 12376 299 12438 333
rect 12376 265 12388 299
rect 12422 265 12438 299
rect 12376 224 12438 265
rect 12468 1183 12534 1224
rect 12468 1149 12484 1183
rect 12518 1149 12534 1183
rect 12468 1115 12534 1149
rect 12468 1081 12484 1115
rect 12518 1081 12534 1115
rect 12468 1047 12534 1081
rect 12468 1013 12484 1047
rect 12518 1013 12534 1047
rect 12468 979 12534 1013
rect 12468 945 12484 979
rect 12518 945 12534 979
rect 12468 911 12534 945
rect 12468 877 12484 911
rect 12518 877 12534 911
rect 12468 843 12534 877
rect 12468 809 12484 843
rect 12518 809 12534 843
rect 12468 775 12534 809
rect 12468 741 12484 775
rect 12518 741 12534 775
rect 12468 707 12534 741
rect 12468 673 12484 707
rect 12518 673 12534 707
rect 12468 639 12534 673
rect 12468 605 12484 639
rect 12518 605 12534 639
rect 12468 571 12534 605
rect 12468 537 12484 571
rect 12518 537 12534 571
rect 12468 503 12534 537
rect 12468 469 12484 503
rect 12518 469 12534 503
rect 12468 435 12534 469
rect 12468 401 12484 435
rect 12518 401 12534 435
rect 12468 367 12534 401
rect 12468 333 12484 367
rect 12518 333 12534 367
rect 12468 299 12534 333
rect 12468 265 12484 299
rect 12518 265 12534 299
rect 12468 224 12534 265
rect 12564 1183 12630 1224
rect 12564 1149 12580 1183
rect 12614 1149 12630 1183
rect 12564 1115 12630 1149
rect 12564 1081 12580 1115
rect 12614 1081 12630 1115
rect 12564 1047 12630 1081
rect 12564 1013 12580 1047
rect 12614 1013 12630 1047
rect 12564 979 12630 1013
rect 12564 945 12580 979
rect 12614 945 12630 979
rect 12564 911 12630 945
rect 12564 877 12580 911
rect 12614 877 12630 911
rect 12564 843 12630 877
rect 12564 809 12580 843
rect 12614 809 12630 843
rect 12564 775 12630 809
rect 12564 741 12580 775
rect 12614 741 12630 775
rect 12564 707 12630 741
rect 12564 673 12580 707
rect 12614 673 12630 707
rect 12564 639 12630 673
rect 12564 605 12580 639
rect 12614 605 12630 639
rect 12564 571 12630 605
rect 12564 537 12580 571
rect 12614 537 12630 571
rect 12564 503 12630 537
rect 12564 469 12580 503
rect 12614 469 12630 503
rect 12564 435 12630 469
rect 12564 401 12580 435
rect 12614 401 12630 435
rect 12564 367 12630 401
rect 12564 333 12580 367
rect 12614 333 12630 367
rect 12564 299 12630 333
rect 12564 265 12580 299
rect 12614 265 12630 299
rect 12564 224 12630 265
rect 12660 1183 12726 1224
rect 12660 1149 12676 1183
rect 12710 1149 12726 1183
rect 12660 1115 12726 1149
rect 12660 1081 12676 1115
rect 12710 1081 12726 1115
rect 12660 1047 12726 1081
rect 12660 1013 12676 1047
rect 12710 1013 12726 1047
rect 12660 979 12726 1013
rect 12660 945 12676 979
rect 12710 945 12726 979
rect 12660 911 12726 945
rect 12660 877 12676 911
rect 12710 877 12726 911
rect 12660 843 12726 877
rect 12660 809 12676 843
rect 12710 809 12726 843
rect 12660 775 12726 809
rect 12660 741 12676 775
rect 12710 741 12726 775
rect 12660 707 12726 741
rect 12660 673 12676 707
rect 12710 673 12726 707
rect 12660 639 12726 673
rect 12660 605 12676 639
rect 12710 605 12726 639
rect 12660 571 12726 605
rect 12660 537 12676 571
rect 12710 537 12726 571
rect 12660 503 12726 537
rect 12660 469 12676 503
rect 12710 469 12726 503
rect 12660 435 12726 469
rect 12660 401 12676 435
rect 12710 401 12726 435
rect 12660 367 12726 401
rect 12660 333 12676 367
rect 12710 333 12726 367
rect 12660 299 12726 333
rect 12660 265 12676 299
rect 12710 265 12726 299
rect 12660 224 12726 265
rect 12756 1183 12822 1224
rect 12756 1149 12772 1183
rect 12806 1149 12822 1183
rect 12756 1115 12822 1149
rect 12756 1081 12772 1115
rect 12806 1081 12822 1115
rect 12756 1047 12822 1081
rect 12756 1013 12772 1047
rect 12806 1013 12822 1047
rect 12756 979 12822 1013
rect 12756 945 12772 979
rect 12806 945 12822 979
rect 12756 911 12822 945
rect 12756 877 12772 911
rect 12806 877 12822 911
rect 12756 843 12822 877
rect 12756 809 12772 843
rect 12806 809 12822 843
rect 12756 775 12822 809
rect 12756 741 12772 775
rect 12806 741 12822 775
rect 12756 707 12822 741
rect 12756 673 12772 707
rect 12806 673 12822 707
rect 12756 639 12822 673
rect 12756 605 12772 639
rect 12806 605 12822 639
rect 12756 571 12822 605
rect 12756 537 12772 571
rect 12806 537 12822 571
rect 12756 503 12822 537
rect 12756 469 12772 503
rect 12806 469 12822 503
rect 12756 435 12822 469
rect 12756 401 12772 435
rect 12806 401 12822 435
rect 12756 367 12822 401
rect 12756 333 12772 367
rect 12806 333 12822 367
rect 12756 299 12822 333
rect 12756 265 12772 299
rect 12806 265 12822 299
rect 12756 224 12822 265
rect 12852 1183 12918 1224
rect 12852 1149 12868 1183
rect 12902 1149 12918 1183
rect 12852 1115 12918 1149
rect 12852 1081 12868 1115
rect 12902 1081 12918 1115
rect 12852 1047 12918 1081
rect 12852 1013 12868 1047
rect 12902 1013 12918 1047
rect 12852 979 12918 1013
rect 12852 945 12868 979
rect 12902 945 12918 979
rect 12852 911 12918 945
rect 12852 877 12868 911
rect 12902 877 12918 911
rect 12852 843 12918 877
rect 12852 809 12868 843
rect 12902 809 12918 843
rect 12852 775 12918 809
rect 12852 741 12868 775
rect 12902 741 12918 775
rect 12852 707 12918 741
rect 12852 673 12868 707
rect 12902 673 12918 707
rect 12852 639 12918 673
rect 12852 605 12868 639
rect 12902 605 12918 639
rect 12852 571 12918 605
rect 12852 537 12868 571
rect 12902 537 12918 571
rect 12852 503 12918 537
rect 12852 469 12868 503
rect 12902 469 12918 503
rect 12852 435 12918 469
rect 12852 401 12868 435
rect 12902 401 12918 435
rect 12852 367 12918 401
rect 12852 333 12868 367
rect 12902 333 12918 367
rect 12852 299 12918 333
rect 12852 265 12868 299
rect 12902 265 12918 299
rect 12852 224 12918 265
rect 12948 1183 13014 1224
rect 12948 1149 12964 1183
rect 12998 1149 13014 1183
rect 12948 1115 13014 1149
rect 12948 1081 12964 1115
rect 12998 1081 13014 1115
rect 12948 1047 13014 1081
rect 12948 1013 12964 1047
rect 12998 1013 13014 1047
rect 12948 979 13014 1013
rect 12948 945 12964 979
rect 12998 945 13014 979
rect 12948 911 13014 945
rect 12948 877 12964 911
rect 12998 877 13014 911
rect 12948 843 13014 877
rect 12948 809 12964 843
rect 12998 809 13014 843
rect 12948 775 13014 809
rect 12948 741 12964 775
rect 12998 741 13014 775
rect 12948 707 13014 741
rect 12948 673 12964 707
rect 12998 673 13014 707
rect 12948 639 13014 673
rect 12948 605 12964 639
rect 12998 605 13014 639
rect 12948 571 13014 605
rect 12948 537 12964 571
rect 12998 537 13014 571
rect 12948 503 13014 537
rect 12948 469 12964 503
rect 12998 469 13014 503
rect 12948 435 13014 469
rect 12948 401 12964 435
rect 12998 401 13014 435
rect 12948 367 13014 401
rect 12948 333 12964 367
rect 12998 333 13014 367
rect 12948 299 13014 333
rect 12948 265 12964 299
rect 12998 265 13014 299
rect 12948 224 13014 265
rect 13044 1183 13110 1224
rect 13044 1149 13060 1183
rect 13094 1149 13110 1183
rect 13044 1115 13110 1149
rect 13044 1081 13060 1115
rect 13094 1081 13110 1115
rect 13044 1047 13110 1081
rect 13044 1013 13060 1047
rect 13094 1013 13110 1047
rect 13044 979 13110 1013
rect 13044 945 13060 979
rect 13094 945 13110 979
rect 13044 911 13110 945
rect 13044 877 13060 911
rect 13094 877 13110 911
rect 13044 843 13110 877
rect 13044 809 13060 843
rect 13094 809 13110 843
rect 13044 775 13110 809
rect 13044 741 13060 775
rect 13094 741 13110 775
rect 13044 707 13110 741
rect 13044 673 13060 707
rect 13094 673 13110 707
rect 13044 639 13110 673
rect 13044 605 13060 639
rect 13094 605 13110 639
rect 13044 571 13110 605
rect 13044 537 13060 571
rect 13094 537 13110 571
rect 13044 503 13110 537
rect 13044 469 13060 503
rect 13094 469 13110 503
rect 13044 435 13110 469
rect 13044 401 13060 435
rect 13094 401 13110 435
rect 13044 367 13110 401
rect 13044 333 13060 367
rect 13094 333 13110 367
rect 13044 299 13110 333
rect 13044 265 13060 299
rect 13094 265 13110 299
rect 13044 224 13110 265
rect 13140 1183 13206 1224
rect 13140 1149 13156 1183
rect 13190 1149 13206 1183
rect 13140 1115 13206 1149
rect 13140 1081 13156 1115
rect 13190 1081 13206 1115
rect 13140 1047 13206 1081
rect 13140 1013 13156 1047
rect 13190 1013 13206 1047
rect 13140 979 13206 1013
rect 13140 945 13156 979
rect 13190 945 13206 979
rect 13140 911 13206 945
rect 13140 877 13156 911
rect 13190 877 13206 911
rect 13140 843 13206 877
rect 13140 809 13156 843
rect 13190 809 13206 843
rect 13140 775 13206 809
rect 13140 741 13156 775
rect 13190 741 13206 775
rect 13140 707 13206 741
rect 13140 673 13156 707
rect 13190 673 13206 707
rect 13140 639 13206 673
rect 13140 605 13156 639
rect 13190 605 13206 639
rect 13140 571 13206 605
rect 13140 537 13156 571
rect 13190 537 13206 571
rect 13140 503 13206 537
rect 13140 469 13156 503
rect 13190 469 13206 503
rect 13140 435 13206 469
rect 13140 401 13156 435
rect 13190 401 13206 435
rect 13140 367 13206 401
rect 13140 333 13156 367
rect 13190 333 13206 367
rect 13140 299 13206 333
rect 13140 265 13156 299
rect 13190 265 13206 299
rect 13140 224 13206 265
rect 13236 1183 13302 1224
rect 13236 1149 13252 1183
rect 13286 1149 13302 1183
rect 13236 1115 13302 1149
rect 13236 1081 13252 1115
rect 13286 1081 13302 1115
rect 13236 1047 13302 1081
rect 13236 1013 13252 1047
rect 13286 1013 13302 1047
rect 13236 979 13302 1013
rect 13236 945 13252 979
rect 13286 945 13302 979
rect 13236 911 13302 945
rect 13236 877 13252 911
rect 13286 877 13302 911
rect 13236 843 13302 877
rect 13236 809 13252 843
rect 13286 809 13302 843
rect 13236 775 13302 809
rect 13236 741 13252 775
rect 13286 741 13302 775
rect 13236 707 13302 741
rect 13236 673 13252 707
rect 13286 673 13302 707
rect 13236 639 13302 673
rect 13236 605 13252 639
rect 13286 605 13302 639
rect 13236 571 13302 605
rect 13236 537 13252 571
rect 13286 537 13302 571
rect 13236 503 13302 537
rect 13236 469 13252 503
rect 13286 469 13302 503
rect 13236 435 13302 469
rect 13236 401 13252 435
rect 13286 401 13302 435
rect 13236 367 13302 401
rect 13236 333 13252 367
rect 13286 333 13302 367
rect 13236 299 13302 333
rect 13236 265 13252 299
rect 13286 265 13302 299
rect 13236 224 13302 265
rect 13332 1183 13398 1224
rect 13332 1149 13348 1183
rect 13382 1149 13398 1183
rect 13332 1115 13398 1149
rect 13332 1081 13348 1115
rect 13382 1081 13398 1115
rect 13332 1047 13398 1081
rect 13332 1013 13348 1047
rect 13382 1013 13398 1047
rect 13332 979 13398 1013
rect 13332 945 13348 979
rect 13382 945 13398 979
rect 13332 911 13398 945
rect 13332 877 13348 911
rect 13382 877 13398 911
rect 13332 843 13398 877
rect 13332 809 13348 843
rect 13382 809 13398 843
rect 13332 775 13398 809
rect 13332 741 13348 775
rect 13382 741 13398 775
rect 13332 707 13398 741
rect 13332 673 13348 707
rect 13382 673 13398 707
rect 13332 639 13398 673
rect 13332 605 13348 639
rect 13382 605 13398 639
rect 13332 571 13398 605
rect 13332 537 13348 571
rect 13382 537 13398 571
rect 13332 503 13398 537
rect 13332 469 13348 503
rect 13382 469 13398 503
rect 13332 435 13398 469
rect 13332 401 13348 435
rect 13382 401 13398 435
rect 13332 367 13398 401
rect 13332 333 13348 367
rect 13382 333 13398 367
rect 13332 299 13398 333
rect 13332 265 13348 299
rect 13382 265 13398 299
rect 13332 224 13398 265
rect 13428 1183 13494 1224
rect 13428 1149 13444 1183
rect 13478 1149 13494 1183
rect 13428 1115 13494 1149
rect 13428 1081 13444 1115
rect 13478 1081 13494 1115
rect 13428 1047 13494 1081
rect 13428 1013 13444 1047
rect 13478 1013 13494 1047
rect 13428 979 13494 1013
rect 13428 945 13444 979
rect 13478 945 13494 979
rect 13428 911 13494 945
rect 13428 877 13444 911
rect 13478 877 13494 911
rect 13428 843 13494 877
rect 13428 809 13444 843
rect 13478 809 13494 843
rect 13428 775 13494 809
rect 13428 741 13444 775
rect 13478 741 13494 775
rect 13428 707 13494 741
rect 13428 673 13444 707
rect 13478 673 13494 707
rect 13428 639 13494 673
rect 13428 605 13444 639
rect 13478 605 13494 639
rect 13428 571 13494 605
rect 13428 537 13444 571
rect 13478 537 13494 571
rect 13428 503 13494 537
rect 13428 469 13444 503
rect 13478 469 13494 503
rect 13428 435 13494 469
rect 13428 401 13444 435
rect 13478 401 13494 435
rect 13428 367 13494 401
rect 13428 333 13444 367
rect 13478 333 13494 367
rect 13428 299 13494 333
rect 13428 265 13444 299
rect 13478 265 13494 299
rect 13428 224 13494 265
rect 13524 1183 13586 1224
rect 13524 1149 13540 1183
rect 13574 1149 13586 1183
rect 13524 1115 13586 1149
rect 13524 1081 13540 1115
rect 13574 1081 13586 1115
rect 13524 1047 13586 1081
rect 13524 1013 13540 1047
rect 13574 1013 13586 1047
rect 13524 979 13586 1013
rect 13524 945 13540 979
rect 13574 945 13586 979
rect 13524 911 13586 945
rect 13524 877 13540 911
rect 13574 877 13586 911
rect 13524 843 13586 877
rect 13524 809 13540 843
rect 13574 809 13586 843
rect 13524 775 13586 809
rect 13524 741 13540 775
rect 13574 741 13586 775
rect 13524 707 13586 741
rect 13524 673 13540 707
rect 13574 673 13586 707
rect 13524 639 13586 673
rect 13524 605 13540 639
rect 13574 605 13586 639
rect 13524 571 13586 605
rect 13524 537 13540 571
rect 13574 537 13586 571
rect 13524 503 13586 537
rect 13524 469 13540 503
rect 13574 469 13586 503
rect 13524 435 13586 469
rect 13524 401 13540 435
rect 13574 401 13586 435
rect 13524 367 13586 401
rect 13524 333 13540 367
rect 13574 333 13586 367
rect 13524 299 13586 333
rect 13524 265 13540 299
rect 13574 265 13586 299
rect 13524 224 13586 265
rect 14144 1183 14206 1224
rect 14144 1149 14156 1183
rect 14190 1149 14206 1183
rect 14144 1115 14206 1149
rect 14144 1081 14156 1115
rect 14190 1081 14206 1115
rect 14144 1047 14206 1081
rect 14144 1013 14156 1047
rect 14190 1013 14206 1047
rect 14144 979 14206 1013
rect 14144 945 14156 979
rect 14190 945 14206 979
rect 14144 911 14206 945
rect 14144 877 14156 911
rect 14190 877 14206 911
rect 14144 843 14206 877
rect 14144 809 14156 843
rect 14190 809 14206 843
rect 14144 775 14206 809
rect 14144 741 14156 775
rect 14190 741 14206 775
rect 14144 707 14206 741
rect 14144 673 14156 707
rect 14190 673 14206 707
rect 14144 639 14206 673
rect 14144 605 14156 639
rect 14190 605 14206 639
rect 14144 571 14206 605
rect 14144 537 14156 571
rect 14190 537 14206 571
rect 14144 503 14206 537
rect 14144 469 14156 503
rect 14190 469 14206 503
rect 14144 435 14206 469
rect 14144 401 14156 435
rect 14190 401 14206 435
rect 14144 367 14206 401
rect 14144 333 14156 367
rect 14190 333 14206 367
rect 14144 299 14206 333
rect 14144 265 14156 299
rect 14190 265 14206 299
rect 14144 224 14206 265
rect 14236 1183 14302 1224
rect 14236 1149 14252 1183
rect 14286 1149 14302 1183
rect 14236 1115 14302 1149
rect 14236 1081 14252 1115
rect 14286 1081 14302 1115
rect 14236 1047 14302 1081
rect 14236 1013 14252 1047
rect 14286 1013 14302 1047
rect 14236 979 14302 1013
rect 14236 945 14252 979
rect 14286 945 14302 979
rect 14236 911 14302 945
rect 14236 877 14252 911
rect 14286 877 14302 911
rect 14236 843 14302 877
rect 14236 809 14252 843
rect 14286 809 14302 843
rect 14236 775 14302 809
rect 14236 741 14252 775
rect 14286 741 14302 775
rect 14236 707 14302 741
rect 14236 673 14252 707
rect 14286 673 14302 707
rect 14236 639 14302 673
rect 14236 605 14252 639
rect 14286 605 14302 639
rect 14236 571 14302 605
rect 14236 537 14252 571
rect 14286 537 14302 571
rect 14236 503 14302 537
rect 14236 469 14252 503
rect 14286 469 14302 503
rect 14236 435 14302 469
rect 14236 401 14252 435
rect 14286 401 14302 435
rect 14236 367 14302 401
rect 14236 333 14252 367
rect 14286 333 14302 367
rect 14236 299 14302 333
rect 14236 265 14252 299
rect 14286 265 14302 299
rect 14236 224 14302 265
rect 14332 1183 14398 1224
rect 14332 1149 14348 1183
rect 14382 1149 14398 1183
rect 14332 1115 14398 1149
rect 14332 1081 14348 1115
rect 14382 1081 14398 1115
rect 14332 1047 14398 1081
rect 14332 1013 14348 1047
rect 14382 1013 14398 1047
rect 14332 979 14398 1013
rect 14332 945 14348 979
rect 14382 945 14398 979
rect 14332 911 14398 945
rect 14332 877 14348 911
rect 14382 877 14398 911
rect 14332 843 14398 877
rect 14332 809 14348 843
rect 14382 809 14398 843
rect 14332 775 14398 809
rect 14332 741 14348 775
rect 14382 741 14398 775
rect 14332 707 14398 741
rect 14332 673 14348 707
rect 14382 673 14398 707
rect 14332 639 14398 673
rect 14332 605 14348 639
rect 14382 605 14398 639
rect 14332 571 14398 605
rect 14332 537 14348 571
rect 14382 537 14398 571
rect 14332 503 14398 537
rect 14332 469 14348 503
rect 14382 469 14398 503
rect 14332 435 14398 469
rect 14332 401 14348 435
rect 14382 401 14398 435
rect 14332 367 14398 401
rect 14332 333 14348 367
rect 14382 333 14398 367
rect 14332 299 14398 333
rect 14332 265 14348 299
rect 14382 265 14398 299
rect 14332 224 14398 265
rect 14428 1183 14494 1224
rect 14428 1149 14444 1183
rect 14478 1149 14494 1183
rect 14428 1115 14494 1149
rect 14428 1081 14444 1115
rect 14478 1081 14494 1115
rect 14428 1047 14494 1081
rect 14428 1013 14444 1047
rect 14478 1013 14494 1047
rect 14428 979 14494 1013
rect 14428 945 14444 979
rect 14478 945 14494 979
rect 14428 911 14494 945
rect 14428 877 14444 911
rect 14478 877 14494 911
rect 14428 843 14494 877
rect 14428 809 14444 843
rect 14478 809 14494 843
rect 14428 775 14494 809
rect 14428 741 14444 775
rect 14478 741 14494 775
rect 14428 707 14494 741
rect 14428 673 14444 707
rect 14478 673 14494 707
rect 14428 639 14494 673
rect 14428 605 14444 639
rect 14478 605 14494 639
rect 14428 571 14494 605
rect 14428 537 14444 571
rect 14478 537 14494 571
rect 14428 503 14494 537
rect 14428 469 14444 503
rect 14478 469 14494 503
rect 14428 435 14494 469
rect 14428 401 14444 435
rect 14478 401 14494 435
rect 14428 367 14494 401
rect 14428 333 14444 367
rect 14478 333 14494 367
rect 14428 299 14494 333
rect 14428 265 14444 299
rect 14478 265 14494 299
rect 14428 224 14494 265
rect 14524 1183 14590 1224
rect 14524 1149 14540 1183
rect 14574 1149 14590 1183
rect 14524 1115 14590 1149
rect 14524 1081 14540 1115
rect 14574 1081 14590 1115
rect 14524 1047 14590 1081
rect 14524 1013 14540 1047
rect 14574 1013 14590 1047
rect 14524 979 14590 1013
rect 14524 945 14540 979
rect 14574 945 14590 979
rect 14524 911 14590 945
rect 14524 877 14540 911
rect 14574 877 14590 911
rect 14524 843 14590 877
rect 14524 809 14540 843
rect 14574 809 14590 843
rect 14524 775 14590 809
rect 14524 741 14540 775
rect 14574 741 14590 775
rect 14524 707 14590 741
rect 14524 673 14540 707
rect 14574 673 14590 707
rect 14524 639 14590 673
rect 14524 605 14540 639
rect 14574 605 14590 639
rect 14524 571 14590 605
rect 14524 537 14540 571
rect 14574 537 14590 571
rect 14524 503 14590 537
rect 14524 469 14540 503
rect 14574 469 14590 503
rect 14524 435 14590 469
rect 14524 401 14540 435
rect 14574 401 14590 435
rect 14524 367 14590 401
rect 14524 333 14540 367
rect 14574 333 14590 367
rect 14524 299 14590 333
rect 14524 265 14540 299
rect 14574 265 14590 299
rect 14524 224 14590 265
rect 14620 1183 14686 1224
rect 14620 1149 14636 1183
rect 14670 1149 14686 1183
rect 14620 1115 14686 1149
rect 14620 1081 14636 1115
rect 14670 1081 14686 1115
rect 14620 1047 14686 1081
rect 14620 1013 14636 1047
rect 14670 1013 14686 1047
rect 14620 979 14686 1013
rect 14620 945 14636 979
rect 14670 945 14686 979
rect 14620 911 14686 945
rect 14620 877 14636 911
rect 14670 877 14686 911
rect 14620 843 14686 877
rect 14620 809 14636 843
rect 14670 809 14686 843
rect 14620 775 14686 809
rect 14620 741 14636 775
rect 14670 741 14686 775
rect 14620 707 14686 741
rect 14620 673 14636 707
rect 14670 673 14686 707
rect 14620 639 14686 673
rect 14620 605 14636 639
rect 14670 605 14686 639
rect 14620 571 14686 605
rect 14620 537 14636 571
rect 14670 537 14686 571
rect 14620 503 14686 537
rect 14620 469 14636 503
rect 14670 469 14686 503
rect 14620 435 14686 469
rect 14620 401 14636 435
rect 14670 401 14686 435
rect 14620 367 14686 401
rect 14620 333 14636 367
rect 14670 333 14686 367
rect 14620 299 14686 333
rect 14620 265 14636 299
rect 14670 265 14686 299
rect 14620 224 14686 265
rect 14716 1183 14782 1224
rect 14716 1149 14732 1183
rect 14766 1149 14782 1183
rect 14716 1115 14782 1149
rect 14716 1081 14732 1115
rect 14766 1081 14782 1115
rect 14716 1047 14782 1081
rect 14716 1013 14732 1047
rect 14766 1013 14782 1047
rect 14716 979 14782 1013
rect 14716 945 14732 979
rect 14766 945 14782 979
rect 14716 911 14782 945
rect 14716 877 14732 911
rect 14766 877 14782 911
rect 14716 843 14782 877
rect 14716 809 14732 843
rect 14766 809 14782 843
rect 14716 775 14782 809
rect 14716 741 14732 775
rect 14766 741 14782 775
rect 14716 707 14782 741
rect 14716 673 14732 707
rect 14766 673 14782 707
rect 14716 639 14782 673
rect 14716 605 14732 639
rect 14766 605 14782 639
rect 14716 571 14782 605
rect 14716 537 14732 571
rect 14766 537 14782 571
rect 14716 503 14782 537
rect 14716 469 14732 503
rect 14766 469 14782 503
rect 14716 435 14782 469
rect 14716 401 14732 435
rect 14766 401 14782 435
rect 14716 367 14782 401
rect 14716 333 14732 367
rect 14766 333 14782 367
rect 14716 299 14782 333
rect 14716 265 14732 299
rect 14766 265 14782 299
rect 14716 224 14782 265
rect 14812 1183 14878 1224
rect 14812 1149 14828 1183
rect 14862 1149 14878 1183
rect 14812 1115 14878 1149
rect 14812 1081 14828 1115
rect 14862 1081 14878 1115
rect 14812 1047 14878 1081
rect 14812 1013 14828 1047
rect 14862 1013 14878 1047
rect 14812 979 14878 1013
rect 14812 945 14828 979
rect 14862 945 14878 979
rect 14812 911 14878 945
rect 14812 877 14828 911
rect 14862 877 14878 911
rect 14812 843 14878 877
rect 14812 809 14828 843
rect 14862 809 14878 843
rect 14812 775 14878 809
rect 14812 741 14828 775
rect 14862 741 14878 775
rect 14812 707 14878 741
rect 14812 673 14828 707
rect 14862 673 14878 707
rect 14812 639 14878 673
rect 14812 605 14828 639
rect 14862 605 14878 639
rect 14812 571 14878 605
rect 14812 537 14828 571
rect 14862 537 14878 571
rect 14812 503 14878 537
rect 14812 469 14828 503
rect 14862 469 14878 503
rect 14812 435 14878 469
rect 14812 401 14828 435
rect 14862 401 14878 435
rect 14812 367 14878 401
rect 14812 333 14828 367
rect 14862 333 14878 367
rect 14812 299 14878 333
rect 14812 265 14828 299
rect 14862 265 14878 299
rect 14812 224 14878 265
rect 14908 1183 14974 1224
rect 14908 1149 14924 1183
rect 14958 1149 14974 1183
rect 14908 1115 14974 1149
rect 14908 1081 14924 1115
rect 14958 1081 14974 1115
rect 14908 1047 14974 1081
rect 14908 1013 14924 1047
rect 14958 1013 14974 1047
rect 14908 979 14974 1013
rect 14908 945 14924 979
rect 14958 945 14974 979
rect 14908 911 14974 945
rect 14908 877 14924 911
rect 14958 877 14974 911
rect 14908 843 14974 877
rect 14908 809 14924 843
rect 14958 809 14974 843
rect 14908 775 14974 809
rect 14908 741 14924 775
rect 14958 741 14974 775
rect 14908 707 14974 741
rect 14908 673 14924 707
rect 14958 673 14974 707
rect 14908 639 14974 673
rect 14908 605 14924 639
rect 14958 605 14974 639
rect 14908 571 14974 605
rect 14908 537 14924 571
rect 14958 537 14974 571
rect 14908 503 14974 537
rect 14908 469 14924 503
rect 14958 469 14974 503
rect 14908 435 14974 469
rect 14908 401 14924 435
rect 14958 401 14974 435
rect 14908 367 14974 401
rect 14908 333 14924 367
rect 14958 333 14974 367
rect 14908 299 14974 333
rect 14908 265 14924 299
rect 14958 265 14974 299
rect 14908 224 14974 265
rect 15004 1183 15070 1224
rect 15004 1149 15020 1183
rect 15054 1149 15070 1183
rect 15004 1115 15070 1149
rect 15004 1081 15020 1115
rect 15054 1081 15070 1115
rect 15004 1047 15070 1081
rect 15004 1013 15020 1047
rect 15054 1013 15070 1047
rect 15004 979 15070 1013
rect 15004 945 15020 979
rect 15054 945 15070 979
rect 15004 911 15070 945
rect 15004 877 15020 911
rect 15054 877 15070 911
rect 15004 843 15070 877
rect 15004 809 15020 843
rect 15054 809 15070 843
rect 15004 775 15070 809
rect 15004 741 15020 775
rect 15054 741 15070 775
rect 15004 707 15070 741
rect 15004 673 15020 707
rect 15054 673 15070 707
rect 15004 639 15070 673
rect 15004 605 15020 639
rect 15054 605 15070 639
rect 15004 571 15070 605
rect 15004 537 15020 571
rect 15054 537 15070 571
rect 15004 503 15070 537
rect 15004 469 15020 503
rect 15054 469 15070 503
rect 15004 435 15070 469
rect 15004 401 15020 435
rect 15054 401 15070 435
rect 15004 367 15070 401
rect 15004 333 15020 367
rect 15054 333 15070 367
rect 15004 299 15070 333
rect 15004 265 15020 299
rect 15054 265 15070 299
rect 15004 224 15070 265
rect 15100 1183 15166 1224
rect 15100 1149 15116 1183
rect 15150 1149 15166 1183
rect 15100 1115 15166 1149
rect 15100 1081 15116 1115
rect 15150 1081 15166 1115
rect 15100 1047 15166 1081
rect 15100 1013 15116 1047
rect 15150 1013 15166 1047
rect 15100 979 15166 1013
rect 15100 945 15116 979
rect 15150 945 15166 979
rect 15100 911 15166 945
rect 15100 877 15116 911
rect 15150 877 15166 911
rect 15100 843 15166 877
rect 15100 809 15116 843
rect 15150 809 15166 843
rect 15100 775 15166 809
rect 15100 741 15116 775
rect 15150 741 15166 775
rect 15100 707 15166 741
rect 15100 673 15116 707
rect 15150 673 15166 707
rect 15100 639 15166 673
rect 15100 605 15116 639
rect 15150 605 15166 639
rect 15100 571 15166 605
rect 15100 537 15116 571
rect 15150 537 15166 571
rect 15100 503 15166 537
rect 15100 469 15116 503
rect 15150 469 15166 503
rect 15100 435 15166 469
rect 15100 401 15116 435
rect 15150 401 15166 435
rect 15100 367 15166 401
rect 15100 333 15116 367
rect 15150 333 15166 367
rect 15100 299 15166 333
rect 15100 265 15116 299
rect 15150 265 15166 299
rect 15100 224 15166 265
rect 15196 1183 15258 1224
rect 15196 1149 15212 1183
rect 15246 1149 15258 1183
rect 15196 1115 15258 1149
rect 15196 1081 15212 1115
rect 15246 1081 15258 1115
rect 15196 1047 15258 1081
rect 15196 1013 15212 1047
rect 15246 1013 15258 1047
rect 15196 979 15258 1013
rect 15196 945 15212 979
rect 15246 945 15258 979
rect 15196 911 15258 945
rect 15196 877 15212 911
rect 15246 877 15258 911
rect 15196 843 15258 877
rect 15196 809 15212 843
rect 15246 809 15258 843
rect 15196 775 15258 809
rect 15196 741 15212 775
rect 15246 741 15258 775
rect 15196 707 15258 741
rect 15196 673 15212 707
rect 15246 673 15258 707
rect 15196 639 15258 673
rect 15196 605 15212 639
rect 15246 605 15258 639
rect 15196 571 15258 605
rect 15196 537 15212 571
rect 15246 537 15258 571
rect 15196 503 15258 537
rect 15196 469 15212 503
rect 15246 469 15258 503
rect 15196 435 15258 469
rect 15196 401 15212 435
rect 15246 401 15258 435
rect 15196 367 15258 401
rect 15196 333 15212 367
rect 15246 333 15258 367
rect 15196 299 15258 333
rect 15196 265 15212 299
rect 15246 265 15258 299
rect 15196 224 15258 265
rect 15410 1193 15468 1227
rect 15410 1159 15422 1193
rect 15456 1159 15468 1193
rect 15410 1125 15468 1159
rect 15410 1091 15422 1125
rect 15456 1091 15468 1125
rect 15410 1057 15468 1091
rect 15410 1023 15422 1057
rect 15456 1023 15468 1057
rect 15410 989 15468 1023
rect 15410 955 15422 989
rect 15456 955 15468 989
rect 15410 921 15468 955
rect 15410 887 15422 921
rect 15456 887 15468 921
rect 15410 853 15468 887
rect 15410 819 15422 853
rect 15456 819 15468 853
rect 15410 785 15468 819
rect 15410 751 15422 785
rect 15456 751 15468 785
rect 15410 717 15468 751
rect 15410 683 15422 717
rect 15456 683 15468 717
rect 15410 649 15468 683
rect 15410 615 15422 649
rect 15456 615 15468 649
rect 15410 581 15468 615
rect 15410 547 15422 581
rect 15456 547 15468 581
rect 15410 513 15468 547
rect 15410 479 15422 513
rect 15456 479 15468 513
rect 15410 445 15468 479
rect 15410 411 15422 445
rect 15456 411 15468 445
rect 15410 377 15468 411
rect 15410 343 15422 377
rect 15456 343 15468 377
rect 15410 309 15468 343
rect 15410 275 15422 309
rect 15456 275 15468 309
rect 15410 241 15468 275
rect 15410 207 15422 241
rect 15456 207 15468 241
rect 15410 173 15468 207
rect 15410 139 15422 173
rect 15456 139 15468 173
rect 15410 100 15468 139
rect 15498 1261 15556 1300
rect 15498 1227 15510 1261
rect 15544 1227 15556 1261
rect 15498 1193 15556 1227
rect 15498 1159 15510 1193
rect 15544 1159 15556 1193
rect 15498 1125 15556 1159
rect 15498 1091 15510 1125
rect 15544 1091 15556 1125
rect 15498 1057 15556 1091
rect 15498 1023 15510 1057
rect 15544 1023 15556 1057
rect 15498 989 15556 1023
rect 15498 955 15510 989
rect 15544 955 15556 989
rect 15498 921 15556 955
rect 15498 887 15510 921
rect 15544 887 15556 921
rect 15498 853 15556 887
rect 15498 819 15510 853
rect 15544 819 15556 853
rect 15498 785 15556 819
rect 15498 751 15510 785
rect 15544 751 15556 785
rect 15498 717 15556 751
rect 15498 683 15510 717
rect 15544 683 15556 717
rect 15498 649 15556 683
rect 15498 615 15510 649
rect 15544 615 15556 649
rect 15498 581 15556 615
rect 15498 547 15510 581
rect 15544 547 15556 581
rect 15498 513 15556 547
rect 15498 479 15510 513
rect 15544 479 15556 513
rect 15498 445 15556 479
rect 15498 411 15510 445
rect 15544 411 15556 445
rect 15498 377 15556 411
rect 15498 343 15510 377
rect 15544 343 15556 377
rect 15498 309 15556 343
rect 15498 275 15510 309
rect 15544 275 15556 309
rect 15498 241 15556 275
rect 15498 207 15510 241
rect 15544 207 15556 241
rect 15498 173 15556 207
rect 15498 139 15510 173
rect 15544 139 15556 173
rect 15498 100 15556 139
<< pdiff >>
rect 182 6565 244 6606
rect 182 6531 194 6565
rect 228 6531 244 6565
rect 182 6497 244 6531
rect 182 6463 194 6497
rect 228 6463 244 6497
rect 182 6429 244 6463
rect 182 6395 194 6429
rect 228 6395 244 6429
rect 182 6361 244 6395
rect 182 6327 194 6361
rect 228 6327 244 6361
rect 182 6293 244 6327
rect 182 6259 194 6293
rect 228 6259 244 6293
rect 182 6225 244 6259
rect 182 6191 194 6225
rect 228 6191 244 6225
rect 182 6157 244 6191
rect 182 6123 194 6157
rect 228 6123 244 6157
rect 182 6089 244 6123
rect 182 6055 194 6089
rect 228 6055 244 6089
rect 182 6021 244 6055
rect 182 5987 194 6021
rect 228 5987 244 6021
rect 182 5953 244 5987
rect -1664 5895 -1606 5936
rect -1664 5861 -1652 5895
rect -1618 5861 -1606 5895
rect -1664 5827 -1606 5861
rect -1664 5793 -1652 5827
rect -1618 5793 -1606 5827
rect -1664 5759 -1606 5793
rect -1664 5725 -1652 5759
rect -1618 5725 -1606 5759
rect -1664 5691 -1606 5725
rect -1664 5657 -1652 5691
rect -1618 5657 -1606 5691
rect -1664 5623 -1606 5657
rect -1664 5589 -1652 5623
rect -1618 5589 -1606 5623
rect -1664 5555 -1606 5589
rect -1664 5521 -1652 5555
rect -1618 5521 -1606 5555
rect -1664 5487 -1606 5521
rect -1664 5453 -1652 5487
rect -1618 5453 -1606 5487
rect -1664 5419 -1606 5453
rect -1664 5385 -1652 5419
rect -1618 5385 -1606 5419
rect -1664 5351 -1606 5385
rect -1664 5317 -1652 5351
rect -1618 5317 -1606 5351
rect -1664 5283 -1606 5317
rect -1664 5249 -1652 5283
rect -1618 5249 -1606 5283
rect -1664 5215 -1606 5249
rect -1664 5181 -1652 5215
rect -1618 5181 -1606 5215
rect -1664 5147 -1606 5181
rect -1664 5113 -1652 5147
rect -1618 5113 -1606 5147
rect -1664 5079 -1606 5113
rect -1664 5045 -1652 5079
rect -1618 5045 -1606 5079
rect -1664 5011 -1606 5045
rect -1664 4977 -1652 5011
rect -1618 4977 -1606 5011
rect -1664 4936 -1606 4977
rect -1566 5895 -1508 5936
rect -1566 5861 -1554 5895
rect -1520 5861 -1508 5895
rect -1566 5827 -1508 5861
rect -1566 5793 -1554 5827
rect -1520 5793 -1508 5827
rect -1566 5759 -1508 5793
rect -1566 5725 -1554 5759
rect -1520 5725 -1508 5759
rect -1566 5691 -1508 5725
rect -1566 5657 -1554 5691
rect -1520 5657 -1508 5691
rect -1566 5623 -1508 5657
rect -1566 5589 -1554 5623
rect -1520 5589 -1508 5623
rect -1566 5555 -1508 5589
rect -1566 5521 -1554 5555
rect -1520 5521 -1508 5555
rect -1566 5487 -1508 5521
rect -1566 5453 -1554 5487
rect -1520 5453 -1508 5487
rect -1566 5419 -1508 5453
rect -1566 5385 -1554 5419
rect -1520 5385 -1508 5419
rect -1566 5351 -1508 5385
rect -1566 5317 -1554 5351
rect -1520 5317 -1508 5351
rect -1566 5283 -1508 5317
rect -1566 5249 -1554 5283
rect -1520 5249 -1508 5283
rect -1566 5215 -1508 5249
rect -1566 5181 -1554 5215
rect -1520 5181 -1508 5215
rect -1566 5147 -1508 5181
rect -1566 5113 -1554 5147
rect -1520 5113 -1508 5147
rect -1566 5079 -1508 5113
rect -1566 5045 -1554 5079
rect -1520 5045 -1508 5079
rect -1566 5011 -1508 5045
rect -1566 4977 -1554 5011
rect -1520 4977 -1508 5011
rect -1566 4936 -1508 4977
rect -1468 5895 -1410 5936
rect -1468 5861 -1456 5895
rect -1422 5861 -1410 5895
rect -1468 5827 -1410 5861
rect -1468 5793 -1456 5827
rect -1422 5793 -1410 5827
rect -1468 5759 -1410 5793
rect -1468 5725 -1456 5759
rect -1422 5725 -1410 5759
rect -1468 5691 -1410 5725
rect -1468 5657 -1456 5691
rect -1422 5657 -1410 5691
rect -1468 5623 -1410 5657
rect -1468 5589 -1456 5623
rect -1422 5589 -1410 5623
rect -1468 5555 -1410 5589
rect -1468 5521 -1456 5555
rect -1422 5521 -1410 5555
rect -1468 5487 -1410 5521
rect -1468 5453 -1456 5487
rect -1422 5453 -1410 5487
rect -1468 5419 -1410 5453
rect -1468 5385 -1456 5419
rect -1422 5385 -1410 5419
rect -1468 5351 -1410 5385
rect -1468 5317 -1456 5351
rect -1422 5317 -1410 5351
rect -1468 5283 -1410 5317
rect -1468 5249 -1456 5283
rect -1422 5249 -1410 5283
rect -1468 5215 -1410 5249
rect -1468 5181 -1456 5215
rect -1422 5181 -1410 5215
rect -1468 5147 -1410 5181
rect -1468 5113 -1456 5147
rect -1422 5113 -1410 5147
rect -1468 5079 -1410 5113
rect -1468 5045 -1456 5079
rect -1422 5045 -1410 5079
rect -1468 5011 -1410 5045
rect -1468 4977 -1456 5011
rect -1422 4977 -1410 5011
rect -1468 4936 -1410 4977
rect -1370 5895 -1312 5936
rect -1370 5861 -1358 5895
rect -1324 5861 -1312 5895
rect -1370 5827 -1312 5861
rect -1370 5793 -1358 5827
rect -1324 5793 -1312 5827
rect -1370 5759 -1312 5793
rect -1370 5725 -1358 5759
rect -1324 5725 -1312 5759
rect -1370 5691 -1312 5725
rect -1370 5657 -1358 5691
rect -1324 5657 -1312 5691
rect -1370 5623 -1312 5657
rect -1370 5589 -1358 5623
rect -1324 5589 -1312 5623
rect -1370 5555 -1312 5589
rect -1370 5521 -1358 5555
rect -1324 5521 -1312 5555
rect -1370 5487 -1312 5521
rect -1370 5453 -1358 5487
rect -1324 5453 -1312 5487
rect -1370 5419 -1312 5453
rect -1370 5385 -1358 5419
rect -1324 5385 -1312 5419
rect -1370 5351 -1312 5385
rect -1370 5317 -1358 5351
rect -1324 5317 -1312 5351
rect -1370 5283 -1312 5317
rect -1370 5249 -1358 5283
rect -1324 5249 -1312 5283
rect -1370 5215 -1312 5249
rect -1370 5181 -1358 5215
rect -1324 5181 -1312 5215
rect -1370 5147 -1312 5181
rect -1370 5113 -1358 5147
rect -1324 5113 -1312 5147
rect -1370 5079 -1312 5113
rect -1370 5045 -1358 5079
rect -1324 5045 -1312 5079
rect -1370 5011 -1312 5045
rect -1370 4977 -1358 5011
rect -1324 4977 -1312 5011
rect -1370 4936 -1312 4977
rect -1272 5895 -1214 5936
rect -1272 5861 -1260 5895
rect -1226 5861 -1214 5895
rect -1272 5827 -1214 5861
rect -1272 5793 -1260 5827
rect -1226 5793 -1214 5827
rect -1272 5759 -1214 5793
rect -1272 5725 -1260 5759
rect -1226 5725 -1214 5759
rect -1272 5691 -1214 5725
rect -1272 5657 -1260 5691
rect -1226 5657 -1214 5691
rect -1272 5623 -1214 5657
rect -1272 5589 -1260 5623
rect -1226 5589 -1214 5623
rect -1272 5555 -1214 5589
rect -1272 5521 -1260 5555
rect -1226 5521 -1214 5555
rect -1272 5487 -1214 5521
rect -1272 5453 -1260 5487
rect -1226 5453 -1214 5487
rect -1272 5419 -1214 5453
rect -1272 5385 -1260 5419
rect -1226 5385 -1214 5419
rect -1272 5351 -1214 5385
rect -1272 5317 -1260 5351
rect -1226 5317 -1214 5351
rect -1272 5283 -1214 5317
rect -1272 5249 -1260 5283
rect -1226 5249 -1214 5283
rect -1272 5215 -1214 5249
rect -1272 5181 -1260 5215
rect -1226 5181 -1214 5215
rect -1272 5147 -1214 5181
rect -1272 5113 -1260 5147
rect -1226 5113 -1214 5147
rect -1272 5079 -1214 5113
rect -1272 5045 -1260 5079
rect -1226 5045 -1214 5079
rect -1272 5011 -1214 5045
rect -1272 4977 -1260 5011
rect -1226 4977 -1214 5011
rect -1272 4936 -1214 4977
rect -1174 5895 -1116 5936
rect -1174 5861 -1162 5895
rect -1128 5861 -1116 5895
rect -1174 5827 -1116 5861
rect -1174 5793 -1162 5827
rect -1128 5793 -1116 5827
rect -1174 5759 -1116 5793
rect -1174 5725 -1162 5759
rect -1128 5725 -1116 5759
rect -1174 5691 -1116 5725
rect -1174 5657 -1162 5691
rect -1128 5657 -1116 5691
rect -1174 5623 -1116 5657
rect -1174 5589 -1162 5623
rect -1128 5589 -1116 5623
rect -1174 5555 -1116 5589
rect -1174 5521 -1162 5555
rect -1128 5521 -1116 5555
rect -1174 5487 -1116 5521
rect -1174 5453 -1162 5487
rect -1128 5453 -1116 5487
rect -1174 5419 -1116 5453
rect -1174 5385 -1162 5419
rect -1128 5385 -1116 5419
rect -1174 5351 -1116 5385
rect -1174 5317 -1162 5351
rect -1128 5317 -1116 5351
rect -1174 5283 -1116 5317
rect -1174 5249 -1162 5283
rect -1128 5249 -1116 5283
rect -1174 5215 -1116 5249
rect -1174 5181 -1162 5215
rect -1128 5181 -1116 5215
rect -1174 5147 -1116 5181
rect -1174 5113 -1162 5147
rect -1128 5113 -1116 5147
rect -1174 5079 -1116 5113
rect -1174 5045 -1162 5079
rect -1128 5045 -1116 5079
rect -1174 5011 -1116 5045
rect -1174 4977 -1162 5011
rect -1128 4977 -1116 5011
rect -1174 4936 -1116 4977
rect -1076 5895 -1018 5936
rect -1076 5861 -1064 5895
rect -1030 5861 -1018 5895
rect -1076 5827 -1018 5861
rect -1076 5793 -1064 5827
rect -1030 5793 -1018 5827
rect -1076 5759 -1018 5793
rect -1076 5725 -1064 5759
rect -1030 5725 -1018 5759
rect -1076 5691 -1018 5725
rect -1076 5657 -1064 5691
rect -1030 5657 -1018 5691
rect -1076 5623 -1018 5657
rect -1076 5589 -1064 5623
rect -1030 5589 -1018 5623
rect -1076 5555 -1018 5589
rect -1076 5521 -1064 5555
rect -1030 5521 -1018 5555
rect -1076 5487 -1018 5521
rect -1076 5453 -1064 5487
rect -1030 5453 -1018 5487
rect -1076 5419 -1018 5453
rect -1076 5385 -1064 5419
rect -1030 5385 -1018 5419
rect -1076 5351 -1018 5385
rect -1076 5317 -1064 5351
rect -1030 5317 -1018 5351
rect -1076 5283 -1018 5317
rect -1076 5249 -1064 5283
rect -1030 5249 -1018 5283
rect -1076 5215 -1018 5249
rect -1076 5181 -1064 5215
rect -1030 5181 -1018 5215
rect -1076 5147 -1018 5181
rect -1076 5113 -1064 5147
rect -1030 5113 -1018 5147
rect -1076 5079 -1018 5113
rect -1076 5045 -1064 5079
rect -1030 5045 -1018 5079
rect -1076 5011 -1018 5045
rect -1076 4977 -1064 5011
rect -1030 4977 -1018 5011
rect -1076 4936 -1018 4977
rect -978 5895 -920 5936
rect -978 5861 -966 5895
rect -932 5861 -920 5895
rect -978 5827 -920 5861
rect -978 5793 -966 5827
rect -932 5793 -920 5827
rect -978 5759 -920 5793
rect -978 5725 -966 5759
rect -932 5725 -920 5759
rect -978 5691 -920 5725
rect -978 5657 -966 5691
rect -932 5657 -920 5691
rect -978 5623 -920 5657
rect -978 5589 -966 5623
rect -932 5589 -920 5623
rect -978 5555 -920 5589
rect -978 5521 -966 5555
rect -932 5521 -920 5555
rect -978 5487 -920 5521
rect -978 5453 -966 5487
rect -932 5453 -920 5487
rect -978 5419 -920 5453
rect -978 5385 -966 5419
rect -932 5385 -920 5419
rect -978 5351 -920 5385
rect -978 5317 -966 5351
rect -932 5317 -920 5351
rect -978 5283 -920 5317
rect -978 5249 -966 5283
rect -932 5249 -920 5283
rect -978 5215 -920 5249
rect -978 5181 -966 5215
rect -932 5181 -920 5215
rect -978 5147 -920 5181
rect -978 5113 -966 5147
rect -932 5113 -920 5147
rect -978 5079 -920 5113
rect -978 5045 -966 5079
rect -932 5045 -920 5079
rect -978 5011 -920 5045
rect -978 4977 -966 5011
rect -932 4977 -920 5011
rect -978 4936 -920 4977
rect -880 5895 -822 5936
rect -880 5861 -868 5895
rect -834 5861 -822 5895
rect -880 5827 -822 5861
rect -880 5793 -868 5827
rect -834 5793 -822 5827
rect -880 5759 -822 5793
rect -880 5725 -868 5759
rect -834 5725 -822 5759
rect -880 5691 -822 5725
rect -880 5657 -868 5691
rect -834 5657 -822 5691
rect -880 5623 -822 5657
rect -880 5589 -868 5623
rect -834 5589 -822 5623
rect 182 5919 194 5953
rect 228 5919 244 5953
rect 182 5885 244 5919
rect 182 5851 194 5885
rect 228 5851 244 5885
rect 182 5817 244 5851
rect 182 5783 194 5817
rect 228 5783 244 5817
rect 182 5749 244 5783
rect 182 5715 194 5749
rect 228 5715 244 5749
rect 182 5681 244 5715
rect 182 5647 194 5681
rect 228 5647 244 5681
rect 182 5606 244 5647
rect 274 6565 340 6606
rect 274 6531 290 6565
rect 324 6531 340 6565
rect 274 6497 340 6531
rect 274 6463 290 6497
rect 324 6463 340 6497
rect 274 6429 340 6463
rect 274 6395 290 6429
rect 324 6395 340 6429
rect 274 6361 340 6395
rect 274 6327 290 6361
rect 324 6327 340 6361
rect 274 6293 340 6327
rect 274 6259 290 6293
rect 324 6259 340 6293
rect 274 6225 340 6259
rect 274 6191 290 6225
rect 324 6191 340 6225
rect 274 6157 340 6191
rect 274 6123 290 6157
rect 324 6123 340 6157
rect 274 6089 340 6123
rect 274 6055 290 6089
rect 324 6055 340 6089
rect 274 6021 340 6055
rect 274 5987 290 6021
rect 324 5987 340 6021
rect 274 5953 340 5987
rect 274 5919 290 5953
rect 324 5919 340 5953
rect 274 5885 340 5919
rect 274 5851 290 5885
rect 324 5851 340 5885
rect 274 5817 340 5851
rect 274 5783 290 5817
rect 324 5783 340 5817
rect 274 5749 340 5783
rect 274 5715 290 5749
rect 324 5715 340 5749
rect 274 5681 340 5715
rect 274 5647 290 5681
rect 324 5647 340 5681
rect 274 5606 340 5647
rect 370 6565 436 6606
rect 370 6531 386 6565
rect 420 6531 436 6565
rect 370 6497 436 6531
rect 370 6463 386 6497
rect 420 6463 436 6497
rect 370 6429 436 6463
rect 370 6395 386 6429
rect 420 6395 436 6429
rect 370 6361 436 6395
rect 370 6327 386 6361
rect 420 6327 436 6361
rect 370 6293 436 6327
rect 370 6259 386 6293
rect 420 6259 436 6293
rect 370 6225 436 6259
rect 370 6191 386 6225
rect 420 6191 436 6225
rect 370 6157 436 6191
rect 370 6123 386 6157
rect 420 6123 436 6157
rect 370 6089 436 6123
rect 370 6055 386 6089
rect 420 6055 436 6089
rect 370 6021 436 6055
rect 370 5987 386 6021
rect 420 5987 436 6021
rect 370 5953 436 5987
rect 370 5919 386 5953
rect 420 5919 436 5953
rect 370 5885 436 5919
rect 370 5851 386 5885
rect 420 5851 436 5885
rect 370 5817 436 5851
rect 370 5783 386 5817
rect 420 5783 436 5817
rect 370 5749 436 5783
rect 370 5715 386 5749
rect 420 5715 436 5749
rect 370 5681 436 5715
rect 370 5647 386 5681
rect 420 5647 436 5681
rect 370 5606 436 5647
rect 466 6565 532 6606
rect 466 6531 482 6565
rect 516 6531 532 6565
rect 466 6497 532 6531
rect 466 6463 482 6497
rect 516 6463 532 6497
rect 466 6429 532 6463
rect 466 6395 482 6429
rect 516 6395 532 6429
rect 466 6361 532 6395
rect 466 6327 482 6361
rect 516 6327 532 6361
rect 466 6293 532 6327
rect 466 6259 482 6293
rect 516 6259 532 6293
rect 466 6225 532 6259
rect 466 6191 482 6225
rect 516 6191 532 6225
rect 466 6157 532 6191
rect 466 6123 482 6157
rect 516 6123 532 6157
rect 466 6089 532 6123
rect 466 6055 482 6089
rect 516 6055 532 6089
rect 466 6021 532 6055
rect 466 5987 482 6021
rect 516 5987 532 6021
rect 466 5953 532 5987
rect 466 5919 482 5953
rect 516 5919 532 5953
rect 466 5885 532 5919
rect 466 5851 482 5885
rect 516 5851 532 5885
rect 466 5817 532 5851
rect 466 5783 482 5817
rect 516 5783 532 5817
rect 466 5749 532 5783
rect 466 5715 482 5749
rect 516 5715 532 5749
rect 466 5681 532 5715
rect 466 5647 482 5681
rect 516 5647 532 5681
rect 466 5606 532 5647
rect 562 6565 628 6606
rect 562 6531 578 6565
rect 612 6531 628 6565
rect 562 6497 628 6531
rect 562 6463 578 6497
rect 612 6463 628 6497
rect 562 6429 628 6463
rect 562 6395 578 6429
rect 612 6395 628 6429
rect 562 6361 628 6395
rect 562 6327 578 6361
rect 612 6327 628 6361
rect 562 6293 628 6327
rect 562 6259 578 6293
rect 612 6259 628 6293
rect 562 6225 628 6259
rect 562 6191 578 6225
rect 612 6191 628 6225
rect 562 6157 628 6191
rect 562 6123 578 6157
rect 612 6123 628 6157
rect 562 6089 628 6123
rect 562 6055 578 6089
rect 612 6055 628 6089
rect 562 6021 628 6055
rect 562 5987 578 6021
rect 612 5987 628 6021
rect 562 5953 628 5987
rect 562 5919 578 5953
rect 612 5919 628 5953
rect 562 5885 628 5919
rect 562 5851 578 5885
rect 612 5851 628 5885
rect 562 5817 628 5851
rect 562 5783 578 5817
rect 612 5783 628 5817
rect 562 5749 628 5783
rect 562 5715 578 5749
rect 612 5715 628 5749
rect 562 5681 628 5715
rect 562 5647 578 5681
rect 612 5647 628 5681
rect 562 5606 628 5647
rect 658 6565 724 6606
rect 658 6531 674 6565
rect 708 6531 724 6565
rect 658 6497 724 6531
rect 658 6463 674 6497
rect 708 6463 724 6497
rect 658 6429 724 6463
rect 658 6395 674 6429
rect 708 6395 724 6429
rect 658 6361 724 6395
rect 658 6327 674 6361
rect 708 6327 724 6361
rect 658 6293 724 6327
rect 658 6259 674 6293
rect 708 6259 724 6293
rect 658 6225 724 6259
rect 658 6191 674 6225
rect 708 6191 724 6225
rect 658 6157 724 6191
rect 658 6123 674 6157
rect 708 6123 724 6157
rect 658 6089 724 6123
rect 658 6055 674 6089
rect 708 6055 724 6089
rect 658 6021 724 6055
rect 658 5987 674 6021
rect 708 5987 724 6021
rect 658 5953 724 5987
rect 658 5919 674 5953
rect 708 5919 724 5953
rect 658 5885 724 5919
rect 658 5851 674 5885
rect 708 5851 724 5885
rect 658 5817 724 5851
rect 658 5783 674 5817
rect 708 5783 724 5817
rect 658 5749 724 5783
rect 658 5715 674 5749
rect 708 5715 724 5749
rect 658 5681 724 5715
rect 658 5647 674 5681
rect 708 5647 724 5681
rect 658 5606 724 5647
rect 754 6565 820 6606
rect 754 6531 770 6565
rect 804 6531 820 6565
rect 754 6497 820 6531
rect 754 6463 770 6497
rect 804 6463 820 6497
rect 754 6429 820 6463
rect 754 6395 770 6429
rect 804 6395 820 6429
rect 754 6361 820 6395
rect 754 6327 770 6361
rect 804 6327 820 6361
rect 754 6293 820 6327
rect 754 6259 770 6293
rect 804 6259 820 6293
rect 754 6225 820 6259
rect 754 6191 770 6225
rect 804 6191 820 6225
rect 754 6157 820 6191
rect 754 6123 770 6157
rect 804 6123 820 6157
rect 754 6089 820 6123
rect 754 6055 770 6089
rect 804 6055 820 6089
rect 754 6021 820 6055
rect 754 5987 770 6021
rect 804 5987 820 6021
rect 754 5953 820 5987
rect 754 5919 770 5953
rect 804 5919 820 5953
rect 754 5885 820 5919
rect 754 5851 770 5885
rect 804 5851 820 5885
rect 754 5817 820 5851
rect 754 5783 770 5817
rect 804 5783 820 5817
rect 754 5749 820 5783
rect 754 5715 770 5749
rect 804 5715 820 5749
rect 754 5681 820 5715
rect 754 5647 770 5681
rect 804 5647 820 5681
rect 754 5606 820 5647
rect 850 6565 916 6606
rect 850 6531 866 6565
rect 900 6531 916 6565
rect 850 6497 916 6531
rect 850 6463 866 6497
rect 900 6463 916 6497
rect 850 6429 916 6463
rect 850 6395 866 6429
rect 900 6395 916 6429
rect 850 6361 916 6395
rect 850 6327 866 6361
rect 900 6327 916 6361
rect 850 6293 916 6327
rect 850 6259 866 6293
rect 900 6259 916 6293
rect 850 6225 916 6259
rect 850 6191 866 6225
rect 900 6191 916 6225
rect 850 6157 916 6191
rect 850 6123 866 6157
rect 900 6123 916 6157
rect 850 6089 916 6123
rect 850 6055 866 6089
rect 900 6055 916 6089
rect 850 6021 916 6055
rect 850 5987 866 6021
rect 900 5987 916 6021
rect 850 5953 916 5987
rect 850 5919 866 5953
rect 900 5919 916 5953
rect 850 5885 916 5919
rect 850 5851 866 5885
rect 900 5851 916 5885
rect 850 5817 916 5851
rect 850 5783 866 5817
rect 900 5783 916 5817
rect 850 5749 916 5783
rect 850 5715 866 5749
rect 900 5715 916 5749
rect 850 5681 916 5715
rect 850 5647 866 5681
rect 900 5647 916 5681
rect 850 5606 916 5647
rect 946 6565 1012 6606
rect 946 6531 962 6565
rect 996 6531 1012 6565
rect 946 6497 1012 6531
rect 946 6463 962 6497
rect 996 6463 1012 6497
rect 946 6429 1012 6463
rect 946 6395 962 6429
rect 996 6395 1012 6429
rect 946 6361 1012 6395
rect 946 6327 962 6361
rect 996 6327 1012 6361
rect 946 6293 1012 6327
rect 946 6259 962 6293
rect 996 6259 1012 6293
rect 946 6225 1012 6259
rect 946 6191 962 6225
rect 996 6191 1012 6225
rect 946 6157 1012 6191
rect 946 6123 962 6157
rect 996 6123 1012 6157
rect 946 6089 1012 6123
rect 946 6055 962 6089
rect 996 6055 1012 6089
rect 946 6021 1012 6055
rect 946 5987 962 6021
rect 996 5987 1012 6021
rect 946 5953 1012 5987
rect 946 5919 962 5953
rect 996 5919 1012 5953
rect 946 5885 1012 5919
rect 946 5851 962 5885
rect 996 5851 1012 5885
rect 946 5817 1012 5851
rect 946 5783 962 5817
rect 996 5783 1012 5817
rect 946 5749 1012 5783
rect 946 5715 962 5749
rect 996 5715 1012 5749
rect 946 5681 1012 5715
rect 946 5647 962 5681
rect 996 5647 1012 5681
rect 946 5606 1012 5647
rect 1042 6565 1108 6606
rect 1042 6531 1058 6565
rect 1092 6531 1108 6565
rect 1042 6497 1108 6531
rect 1042 6463 1058 6497
rect 1092 6463 1108 6497
rect 1042 6429 1108 6463
rect 1042 6395 1058 6429
rect 1092 6395 1108 6429
rect 1042 6361 1108 6395
rect 1042 6327 1058 6361
rect 1092 6327 1108 6361
rect 1042 6293 1108 6327
rect 1042 6259 1058 6293
rect 1092 6259 1108 6293
rect 1042 6225 1108 6259
rect 1042 6191 1058 6225
rect 1092 6191 1108 6225
rect 1042 6157 1108 6191
rect 1042 6123 1058 6157
rect 1092 6123 1108 6157
rect 1042 6089 1108 6123
rect 1042 6055 1058 6089
rect 1092 6055 1108 6089
rect 1042 6021 1108 6055
rect 1042 5987 1058 6021
rect 1092 5987 1108 6021
rect 1042 5953 1108 5987
rect 1042 5919 1058 5953
rect 1092 5919 1108 5953
rect 1042 5885 1108 5919
rect 1042 5851 1058 5885
rect 1092 5851 1108 5885
rect 1042 5817 1108 5851
rect 1042 5783 1058 5817
rect 1092 5783 1108 5817
rect 1042 5749 1108 5783
rect 1042 5715 1058 5749
rect 1092 5715 1108 5749
rect 1042 5681 1108 5715
rect 1042 5647 1058 5681
rect 1092 5647 1108 5681
rect 1042 5606 1108 5647
rect 1138 6565 1204 6606
rect 1138 6531 1154 6565
rect 1188 6531 1204 6565
rect 1138 6497 1204 6531
rect 1138 6463 1154 6497
rect 1188 6463 1204 6497
rect 1138 6429 1204 6463
rect 1138 6395 1154 6429
rect 1188 6395 1204 6429
rect 1138 6361 1204 6395
rect 1138 6327 1154 6361
rect 1188 6327 1204 6361
rect 1138 6293 1204 6327
rect 1138 6259 1154 6293
rect 1188 6259 1204 6293
rect 1138 6225 1204 6259
rect 1138 6191 1154 6225
rect 1188 6191 1204 6225
rect 1138 6157 1204 6191
rect 1138 6123 1154 6157
rect 1188 6123 1204 6157
rect 1138 6089 1204 6123
rect 1138 6055 1154 6089
rect 1188 6055 1204 6089
rect 1138 6021 1204 6055
rect 1138 5987 1154 6021
rect 1188 5987 1204 6021
rect 1138 5953 1204 5987
rect 1138 5919 1154 5953
rect 1188 5919 1204 5953
rect 1138 5885 1204 5919
rect 1138 5851 1154 5885
rect 1188 5851 1204 5885
rect 1138 5817 1204 5851
rect 1138 5783 1154 5817
rect 1188 5783 1204 5817
rect 1138 5749 1204 5783
rect 1138 5715 1154 5749
rect 1188 5715 1204 5749
rect 1138 5681 1204 5715
rect 1138 5647 1154 5681
rect 1188 5647 1204 5681
rect 1138 5606 1204 5647
rect 1234 6565 1300 6606
rect 1234 6531 1250 6565
rect 1284 6531 1300 6565
rect 1234 6497 1300 6531
rect 1234 6463 1250 6497
rect 1284 6463 1300 6497
rect 1234 6429 1300 6463
rect 1234 6395 1250 6429
rect 1284 6395 1300 6429
rect 1234 6361 1300 6395
rect 1234 6327 1250 6361
rect 1284 6327 1300 6361
rect 1234 6293 1300 6327
rect 1234 6259 1250 6293
rect 1284 6259 1300 6293
rect 1234 6225 1300 6259
rect 1234 6191 1250 6225
rect 1284 6191 1300 6225
rect 1234 6157 1300 6191
rect 1234 6123 1250 6157
rect 1284 6123 1300 6157
rect 1234 6089 1300 6123
rect 1234 6055 1250 6089
rect 1284 6055 1300 6089
rect 1234 6021 1300 6055
rect 1234 5987 1250 6021
rect 1284 5987 1300 6021
rect 1234 5953 1300 5987
rect 1234 5919 1250 5953
rect 1284 5919 1300 5953
rect 1234 5885 1300 5919
rect 1234 5851 1250 5885
rect 1284 5851 1300 5885
rect 1234 5817 1300 5851
rect 1234 5783 1250 5817
rect 1284 5783 1300 5817
rect 1234 5749 1300 5783
rect 1234 5715 1250 5749
rect 1284 5715 1300 5749
rect 1234 5681 1300 5715
rect 1234 5647 1250 5681
rect 1284 5647 1300 5681
rect 1234 5606 1300 5647
rect 1330 6565 1392 6606
rect 1330 6531 1346 6565
rect 1380 6531 1392 6565
rect 1330 6497 1392 6531
rect 1330 6463 1346 6497
rect 1380 6463 1392 6497
rect 1330 6429 1392 6463
rect 1330 6395 1346 6429
rect 1380 6395 1392 6429
rect 1330 6361 1392 6395
rect 1330 6327 1346 6361
rect 1380 6327 1392 6361
rect 1330 6293 1392 6327
rect 1330 6259 1346 6293
rect 1380 6259 1392 6293
rect 1330 6225 1392 6259
rect 1330 6191 1346 6225
rect 1380 6191 1392 6225
rect 1330 6157 1392 6191
rect 1330 6123 1346 6157
rect 1380 6123 1392 6157
rect 1330 6089 1392 6123
rect 1330 6055 1346 6089
rect 1380 6055 1392 6089
rect 1330 6021 1392 6055
rect 1330 5987 1346 6021
rect 1380 5987 1392 6021
rect 1330 5953 1392 5987
rect 1330 5919 1346 5953
rect 1380 5919 1392 5953
rect 1330 5885 1392 5919
rect 1330 5851 1346 5885
rect 1380 5851 1392 5885
rect 1330 5817 1392 5851
rect 1330 5783 1346 5817
rect 1380 5783 1392 5817
rect 1330 5749 1392 5783
rect 1330 5715 1346 5749
rect 1380 5715 1392 5749
rect 1330 5681 1392 5715
rect 1330 5647 1346 5681
rect 1380 5647 1392 5681
rect 1330 5606 1392 5647
rect 1948 6561 2010 6602
rect 1948 6527 1960 6561
rect 1994 6527 2010 6561
rect 1948 6493 2010 6527
rect 1948 6459 1960 6493
rect 1994 6459 2010 6493
rect 1948 6425 2010 6459
rect 1948 6391 1960 6425
rect 1994 6391 2010 6425
rect 1948 6357 2010 6391
rect 1948 6323 1960 6357
rect 1994 6323 2010 6357
rect 1948 6289 2010 6323
rect 1948 6255 1960 6289
rect 1994 6255 2010 6289
rect 1948 6221 2010 6255
rect 1948 6187 1960 6221
rect 1994 6187 2010 6221
rect 1948 6153 2010 6187
rect 1948 6119 1960 6153
rect 1994 6119 2010 6153
rect 1948 6085 2010 6119
rect 1948 6051 1960 6085
rect 1994 6051 2010 6085
rect 1948 6017 2010 6051
rect 1948 5983 1960 6017
rect 1994 5983 2010 6017
rect 1948 5949 2010 5983
rect 1948 5915 1960 5949
rect 1994 5915 2010 5949
rect 1948 5881 2010 5915
rect 1948 5847 1960 5881
rect 1994 5847 2010 5881
rect 1948 5813 2010 5847
rect 1948 5779 1960 5813
rect 1994 5779 2010 5813
rect 1948 5745 2010 5779
rect 1948 5711 1960 5745
rect 1994 5711 2010 5745
rect 1948 5677 2010 5711
rect 1948 5643 1960 5677
rect 1994 5643 2010 5677
rect -880 5555 -822 5589
rect 1948 5602 2010 5643
rect 2040 6561 2106 6602
rect 2040 6527 2056 6561
rect 2090 6527 2106 6561
rect 2040 6493 2106 6527
rect 2040 6459 2056 6493
rect 2090 6459 2106 6493
rect 2040 6425 2106 6459
rect 2040 6391 2056 6425
rect 2090 6391 2106 6425
rect 2040 6357 2106 6391
rect 2040 6323 2056 6357
rect 2090 6323 2106 6357
rect 2040 6289 2106 6323
rect 2040 6255 2056 6289
rect 2090 6255 2106 6289
rect 2040 6221 2106 6255
rect 2040 6187 2056 6221
rect 2090 6187 2106 6221
rect 2040 6153 2106 6187
rect 2040 6119 2056 6153
rect 2090 6119 2106 6153
rect 2040 6085 2106 6119
rect 2040 6051 2056 6085
rect 2090 6051 2106 6085
rect 2040 6017 2106 6051
rect 2040 5983 2056 6017
rect 2090 5983 2106 6017
rect 2040 5949 2106 5983
rect 2040 5915 2056 5949
rect 2090 5915 2106 5949
rect 2040 5881 2106 5915
rect 2040 5847 2056 5881
rect 2090 5847 2106 5881
rect 2040 5813 2106 5847
rect 2040 5779 2056 5813
rect 2090 5779 2106 5813
rect 2040 5745 2106 5779
rect 2040 5711 2056 5745
rect 2090 5711 2106 5745
rect 2040 5677 2106 5711
rect 2040 5643 2056 5677
rect 2090 5643 2106 5677
rect 2040 5602 2106 5643
rect 2136 6561 2202 6602
rect 2136 6527 2152 6561
rect 2186 6527 2202 6561
rect 2136 6493 2202 6527
rect 2136 6459 2152 6493
rect 2186 6459 2202 6493
rect 2136 6425 2202 6459
rect 2136 6391 2152 6425
rect 2186 6391 2202 6425
rect 2136 6357 2202 6391
rect 2136 6323 2152 6357
rect 2186 6323 2202 6357
rect 2136 6289 2202 6323
rect 2136 6255 2152 6289
rect 2186 6255 2202 6289
rect 2136 6221 2202 6255
rect 2136 6187 2152 6221
rect 2186 6187 2202 6221
rect 2136 6153 2202 6187
rect 2136 6119 2152 6153
rect 2186 6119 2202 6153
rect 2136 6085 2202 6119
rect 2136 6051 2152 6085
rect 2186 6051 2202 6085
rect 2136 6017 2202 6051
rect 2136 5983 2152 6017
rect 2186 5983 2202 6017
rect 2136 5949 2202 5983
rect 2136 5915 2152 5949
rect 2186 5915 2202 5949
rect 2136 5881 2202 5915
rect 2136 5847 2152 5881
rect 2186 5847 2202 5881
rect 2136 5813 2202 5847
rect 2136 5779 2152 5813
rect 2186 5779 2202 5813
rect 2136 5745 2202 5779
rect 2136 5711 2152 5745
rect 2186 5711 2202 5745
rect 2136 5677 2202 5711
rect 2136 5643 2152 5677
rect 2186 5643 2202 5677
rect 2136 5602 2202 5643
rect 2232 6561 2298 6602
rect 2232 6527 2248 6561
rect 2282 6527 2298 6561
rect 2232 6493 2298 6527
rect 2232 6459 2248 6493
rect 2282 6459 2298 6493
rect 2232 6425 2298 6459
rect 2232 6391 2248 6425
rect 2282 6391 2298 6425
rect 2232 6357 2298 6391
rect 2232 6323 2248 6357
rect 2282 6323 2298 6357
rect 2232 6289 2298 6323
rect 2232 6255 2248 6289
rect 2282 6255 2298 6289
rect 2232 6221 2298 6255
rect 2232 6187 2248 6221
rect 2282 6187 2298 6221
rect 2232 6153 2298 6187
rect 2232 6119 2248 6153
rect 2282 6119 2298 6153
rect 2232 6085 2298 6119
rect 2232 6051 2248 6085
rect 2282 6051 2298 6085
rect 2232 6017 2298 6051
rect 2232 5983 2248 6017
rect 2282 5983 2298 6017
rect 2232 5949 2298 5983
rect 2232 5915 2248 5949
rect 2282 5915 2298 5949
rect 2232 5881 2298 5915
rect 2232 5847 2248 5881
rect 2282 5847 2298 5881
rect 2232 5813 2298 5847
rect 2232 5779 2248 5813
rect 2282 5779 2298 5813
rect 2232 5745 2298 5779
rect 2232 5711 2248 5745
rect 2282 5711 2298 5745
rect 2232 5677 2298 5711
rect 2232 5643 2248 5677
rect 2282 5643 2298 5677
rect 2232 5602 2298 5643
rect 2328 6561 2394 6602
rect 2328 6527 2344 6561
rect 2378 6527 2394 6561
rect 2328 6493 2394 6527
rect 2328 6459 2344 6493
rect 2378 6459 2394 6493
rect 2328 6425 2394 6459
rect 2328 6391 2344 6425
rect 2378 6391 2394 6425
rect 2328 6357 2394 6391
rect 2328 6323 2344 6357
rect 2378 6323 2394 6357
rect 2328 6289 2394 6323
rect 2328 6255 2344 6289
rect 2378 6255 2394 6289
rect 2328 6221 2394 6255
rect 2328 6187 2344 6221
rect 2378 6187 2394 6221
rect 2328 6153 2394 6187
rect 2328 6119 2344 6153
rect 2378 6119 2394 6153
rect 2328 6085 2394 6119
rect 2328 6051 2344 6085
rect 2378 6051 2394 6085
rect 2328 6017 2394 6051
rect 2328 5983 2344 6017
rect 2378 5983 2394 6017
rect 2328 5949 2394 5983
rect 2328 5915 2344 5949
rect 2378 5915 2394 5949
rect 2328 5881 2394 5915
rect 2328 5847 2344 5881
rect 2378 5847 2394 5881
rect 2328 5813 2394 5847
rect 2328 5779 2344 5813
rect 2378 5779 2394 5813
rect 2328 5745 2394 5779
rect 2328 5711 2344 5745
rect 2378 5711 2394 5745
rect 2328 5677 2394 5711
rect 2328 5643 2344 5677
rect 2378 5643 2394 5677
rect 2328 5602 2394 5643
rect 2424 6561 2490 6602
rect 2424 6527 2440 6561
rect 2474 6527 2490 6561
rect 2424 6493 2490 6527
rect 2424 6459 2440 6493
rect 2474 6459 2490 6493
rect 2424 6425 2490 6459
rect 2424 6391 2440 6425
rect 2474 6391 2490 6425
rect 2424 6357 2490 6391
rect 2424 6323 2440 6357
rect 2474 6323 2490 6357
rect 2424 6289 2490 6323
rect 2424 6255 2440 6289
rect 2474 6255 2490 6289
rect 2424 6221 2490 6255
rect 2424 6187 2440 6221
rect 2474 6187 2490 6221
rect 2424 6153 2490 6187
rect 2424 6119 2440 6153
rect 2474 6119 2490 6153
rect 2424 6085 2490 6119
rect 2424 6051 2440 6085
rect 2474 6051 2490 6085
rect 2424 6017 2490 6051
rect 2424 5983 2440 6017
rect 2474 5983 2490 6017
rect 2424 5949 2490 5983
rect 2424 5915 2440 5949
rect 2474 5915 2490 5949
rect 2424 5881 2490 5915
rect 2424 5847 2440 5881
rect 2474 5847 2490 5881
rect 2424 5813 2490 5847
rect 2424 5779 2440 5813
rect 2474 5779 2490 5813
rect 2424 5745 2490 5779
rect 2424 5711 2440 5745
rect 2474 5711 2490 5745
rect 2424 5677 2490 5711
rect 2424 5643 2440 5677
rect 2474 5643 2490 5677
rect 2424 5602 2490 5643
rect 2520 6561 2586 6602
rect 2520 6527 2536 6561
rect 2570 6527 2586 6561
rect 2520 6493 2586 6527
rect 2520 6459 2536 6493
rect 2570 6459 2586 6493
rect 2520 6425 2586 6459
rect 2520 6391 2536 6425
rect 2570 6391 2586 6425
rect 2520 6357 2586 6391
rect 2520 6323 2536 6357
rect 2570 6323 2586 6357
rect 2520 6289 2586 6323
rect 2520 6255 2536 6289
rect 2570 6255 2586 6289
rect 2520 6221 2586 6255
rect 2520 6187 2536 6221
rect 2570 6187 2586 6221
rect 2520 6153 2586 6187
rect 2520 6119 2536 6153
rect 2570 6119 2586 6153
rect 2520 6085 2586 6119
rect 2520 6051 2536 6085
rect 2570 6051 2586 6085
rect 2520 6017 2586 6051
rect 2520 5983 2536 6017
rect 2570 5983 2586 6017
rect 2520 5949 2586 5983
rect 2520 5915 2536 5949
rect 2570 5915 2586 5949
rect 2520 5881 2586 5915
rect 2520 5847 2536 5881
rect 2570 5847 2586 5881
rect 2520 5813 2586 5847
rect 2520 5779 2536 5813
rect 2570 5779 2586 5813
rect 2520 5745 2586 5779
rect 2520 5711 2536 5745
rect 2570 5711 2586 5745
rect 2520 5677 2586 5711
rect 2520 5643 2536 5677
rect 2570 5643 2586 5677
rect 2520 5602 2586 5643
rect 2616 6561 2682 6602
rect 2616 6527 2632 6561
rect 2666 6527 2682 6561
rect 2616 6493 2682 6527
rect 2616 6459 2632 6493
rect 2666 6459 2682 6493
rect 2616 6425 2682 6459
rect 2616 6391 2632 6425
rect 2666 6391 2682 6425
rect 2616 6357 2682 6391
rect 2616 6323 2632 6357
rect 2666 6323 2682 6357
rect 2616 6289 2682 6323
rect 2616 6255 2632 6289
rect 2666 6255 2682 6289
rect 2616 6221 2682 6255
rect 2616 6187 2632 6221
rect 2666 6187 2682 6221
rect 2616 6153 2682 6187
rect 2616 6119 2632 6153
rect 2666 6119 2682 6153
rect 2616 6085 2682 6119
rect 2616 6051 2632 6085
rect 2666 6051 2682 6085
rect 2616 6017 2682 6051
rect 2616 5983 2632 6017
rect 2666 5983 2682 6017
rect 2616 5949 2682 5983
rect 2616 5915 2632 5949
rect 2666 5915 2682 5949
rect 2616 5881 2682 5915
rect 2616 5847 2632 5881
rect 2666 5847 2682 5881
rect 2616 5813 2682 5847
rect 2616 5779 2632 5813
rect 2666 5779 2682 5813
rect 2616 5745 2682 5779
rect 2616 5711 2632 5745
rect 2666 5711 2682 5745
rect 2616 5677 2682 5711
rect 2616 5643 2632 5677
rect 2666 5643 2682 5677
rect 2616 5602 2682 5643
rect 2712 6561 2774 6602
rect 2712 6527 2728 6561
rect 2762 6527 2774 6561
rect 2712 6493 2774 6527
rect 2712 6459 2728 6493
rect 2762 6459 2774 6493
rect 2712 6425 2774 6459
rect 2712 6391 2728 6425
rect 2762 6391 2774 6425
rect 2712 6357 2774 6391
rect 2712 6323 2728 6357
rect 2762 6323 2774 6357
rect 2712 6289 2774 6323
rect 2712 6255 2728 6289
rect 2762 6255 2774 6289
rect 2712 6221 2774 6255
rect 2712 6187 2728 6221
rect 2762 6187 2774 6221
rect 2712 6153 2774 6187
rect 2712 6119 2728 6153
rect 2762 6119 2774 6153
rect 2712 6085 2774 6119
rect 2712 6051 2728 6085
rect 2762 6051 2774 6085
rect 2712 6017 2774 6051
rect 2712 5983 2728 6017
rect 2762 5983 2774 6017
rect 2712 5949 2774 5983
rect 2712 5915 2728 5949
rect 2762 5915 2774 5949
rect 2712 5881 2774 5915
rect 2712 5847 2728 5881
rect 2762 5847 2774 5881
rect 2712 5813 2774 5847
rect 2712 5779 2728 5813
rect 2762 5779 2774 5813
rect 2712 5745 2774 5779
rect 2712 5711 2728 5745
rect 2762 5711 2774 5745
rect 2712 5677 2774 5711
rect 2712 5643 2728 5677
rect 2762 5643 2774 5677
rect 2712 5602 2774 5643
rect 3138 6549 3200 6590
rect 3138 6515 3150 6549
rect 3184 6515 3200 6549
rect 3138 6481 3200 6515
rect 3138 6447 3150 6481
rect 3184 6447 3200 6481
rect 3138 6413 3200 6447
rect 3138 6379 3150 6413
rect 3184 6379 3200 6413
rect 3138 6345 3200 6379
rect 3138 6311 3150 6345
rect 3184 6311 3200 6345
rect 3138 6277 3200 6311
rect 3138 6243 3150 6277
rect 3184 6243 3200 6277
rect 3138 6209 3200 6243
rect 3138 6175 3150 6209
rect 3184 6175 3200 6209
rect 3138 6141 3200 6175
rect 3138 6107 3150 6141
rect 3184 6107 3200 6141
rect 3138 6073 3200 6107
rect 3138 6039 3150 6073
rect 3184 6039 3200 6073
rect 3138 6005 3200 6039
rect 3138 5971 3150 6005
rect 3184 5971 3200 6005
rect 3138 5937 3200 5971
rect 3138 5903 3150 5937
rect 3184 5903 3200 5937
rect 3138 5869 3200 5903
rect 3138 5835 3150 5869
rect 3184 5835 3200 5869
rect 3138 5801 3200 5835
rect 3138 5767 3150 5801
rect 3184 5767 3200 5801
rect 3138 5733 3200 5767
rect 3138 5699 3150 5733
rect 3184 5699 3200 5733
rect 3138 5665 3200 5699
rect 3138 5631 3150 5665
rect 3184 5631 3200 5665
rect 3138 5590 3200 5631
rect 3230 6549 3296 6590
rect 3230 6515 3246 6549
rect 3280 6515 3296 6549
rect 3230 6481 3296 6515
rect 3230 6447 3246 6481
rect 3280 6447 3296 6481
rect 3230 6413 3296 6447
rect 3230 6379 3246 6413
rect 3280 6379 3296 6413
rect 3230 6345 3296 6379
rect 3230 6311 3246 6345
rect 3280 6311 3296 6345
rect 3230 6277 3296 6311
rect 3230 6243 3246 6277
rect 3280 6243 3296 6277
rect 3230 6209 3296 6243
rect 3230 6175 3246 6209
rect 3280 6175 3296 6209
rect 3230 6141 3296 6175
rect 3230 6107 3246 6141
rect 3280 6107 3296 6141
rect 3230 6073 3296 6107
rect 3230 6039 3246 6073
rect 3280 6039 3296 6073
rect 3230 6005 3296 6039
rect 3230 5971 3246 6005
rect 3280 5971 3296 6005
rect 3230 5937 3296 5971
rect 3230 5903 3246 5937
rect 3280 5903 3296 5937
rect 3230 5869 3296 5903
rect 3230 5835 3246 5869
rect 3280 5835 3296 5869
rect 3230 5801 3296 5835
rect 3230 5767 3246 5801
rect 3280 5767 3296 5801
rect 3230 5733 3296 5767
rect 3230 5699 3246 5733
rect 3280 5699 3296 5733
rect 3230 5665 3296 5699
rect 3230 5631 3246 5665
rect 3280 5631 3296 5665
rect 3230 5590 3296 5631
rect 3326 6549 3392 6590
rect 3326 6515 3342 6549
rect 3376 6515 3392 6549
rect 3326 6481 3392 6515
rect 3326 6447 3342 6481
rect 3376 6447 3392 6481
rect 3326 6413 3392 6447
rect 3326 6379 3342 6413
rect 3376 6379 3392 6413
rect 3326 6345 3392 6379
rect 3326 6311 3342 6345
rect 3376 6311 3392 6345
rect 3326 6277 3392 6311
rect 3326 6243 3342 6277
rect 3376 6243 3392 6277
rect 3326 6209 3392 6243
rect 3326 6175 3342 6209
rect 3376 6175 3392 6209
rect 3326 6141 3392 6175
rect 3326 6107 3342 6141
rect 3376 6107 3392 6141
rect 3326 6073 3392 6107
rect 3326 6039 3342 6073
rect 3376 6039 3392 6073
rect 3326 6005 3392 6039
rect 3326 5971 3342 6005
rect 3376 5971 3392 6005
rect 3326 5937 3392 5971
rect 3326 5903 3342 5937
rect 3376 5903 3392 5937
rect 3326 5869 3392 5903
rect 3326 5835 3342 5869
rect 3376 5835 3392 5869
rect 3326 5801 3392 5835
rect 3326 5767 3342 5801
rect 3376 5767 3392 5801
rect 3326 5733 3392 5767
rect 3326 5699 3342 5733
rect 3376 5699 3392 5733
rect 3326 5665 3392 5699
rect 3326 5631 3342 5665
rect 3376 5631 3392 5665
rect 3326 5590 3392 5631
rect 3422 6549 3488 6590
rect 3422 6515 3438 6549
rect 3472 6515 3488 6549
rect 3422 6481 3488 6515
rect 3422 6447 3438 6481
rect 3472 6447 3488 6481
rect 3422 6413 3488 6447
rect 3422 6379 3438 6413
rect 3472 6379 3488 6413
rect 3422 6345 3488 6379
rect 3422 6311 3438 6345
rect 3472 6311 3488 6345
rect 3422 6277 3488 6311
rect 3422 6243 3438 6277
rect 3472 6243 3488 6277
rect 3422 6209 3488 6243
rect 3422 6175 3438 6209
rect 3472 6175 3488 6209
rect 3422 6141 3488 6175
rect 3422 6107 3438 6141
rect 3472 6107 3488 6141
rect 3422 6073 3488 6107
rect 3422 6039 3438 6073
rect 3472 6039 3488 6073
rect 3422 6005 3488 6039
rect 3422 5971 3438 6005
rect 3472 5971 3488 6005
rect 3422 5937 3488 5971
rect 3422 5903 3438 5937
rect 3472 5903 3488 5937
rect 3422 5869 3488 5903
rect 3422 5835 3438 5869
rect 3472 5835 3488 5869
rect 3422 5801 3488 5835
rect 3422 5767 3438 5801
rect 3472 5767 3488 5801
rect 3422 5733 3488 5767
rect 3422 5699 3438 5733
rect 3472 5699 3488 5733
rect 3422 5665 3488 5699
rect 3422 5631 3438 5665
rect 3472 5631 3488 5665
rect 3422 5590 3488 5631
rect 3518 6549 3584 6590
rect 3518 6515 3534 6549
rect 3568 6515 3584 6549
rect 3518 6481 3584 6515
rect 3518 6447 3534 6481
rect 3568 6447 3584 6481
rect 3518 6413 3584 6447
rect 3518 6379 3534 6413
rect 3568 6379 3584 6413
rect 3518 6345 3584 6379
rect 3518 6311 3534 6345
rect 3568 6311 3584 6345
rect 3518 6277 3584 6311
rect 3518 6243 3534 6277
rect 3568 6243 3584 6277
rect 3518 6209 3584 6243
rect 3518 6175 3534 6209
rect 3568 6175 3584 6209
rect 3518 6141 3584 6175
rect 3518 6107 3534 6141
rect 3568 6107 3584 6141
rect 3518 6073 3584 6107
rect 3518 6039 3534 6073
rect 3568 6039 3584 6073
rect 3518 6005 3584 6039
rect 3518 5971 3534 6005
rect 3568 5971 3584 6005
rect 3518 5937 3584 5971
rect 3518 5903 3534 5937
rect 3568 5903 3584 5937
rect 3518 5869 3584 5903
rect 3518 5835 3534 5869
rect 3568 5835 3584 5869
rect 3518 5801 3584 5835
rect 3518 5767 3534 5801
rect 3568 5767 3584 5801
rect 3518 5733 3584 5767
rect 3518 5699 3534 5733
rect 3568 5699 3584 5733
rect 3518 5665 3584 5699
rect 3518 5631 3534 5665
rect 3568 5631 3584 5665
rect 3518 5590 3584 5631
rect 3614 6549 3680 6590
rect 3614 6515 3630 6549
rect 3664 6515 3680 6549
rect 3614 6481 3680 6515
rect 3614 6447 3630 6481
rect 3664 6447 3680 6481
rect 3614 6413 3680 6447
rect 3614 6379 3630 6413
rect 3664 6379 3680 6413
rect 3614 6345 3680 6379
rect 3614 6311 3630 6345
rect 3664 6311 3680 6345
rect 3614 6277 3680 6311
rect 3614 6243 3630 6277
rect 3664 6243 3680 6277
rect 3614 6209 3680 6243
rect 3614 6175 3630 6209
rect 3664 6175 3680 6209
rect 3614 6141 3680 6175
rect 3614 6107 3630 6141
rect 3664 6107 3680 6141
rect 3614 6073 3680 6107
rect 3614 6039 3630 6073
rect 3664 6039 3680 6073
rect 3614 6005 3680 6039
rect 3614 5971 3630 6005
rect 3664 5971 3680 6005
rect 3614 5937 3680 5971
rect 3614 5903 3630 5937
rect 3664 5903 3680 5937
rect 3614 5869 3680 5903
rect 3614 5835 3630 5869
rect 3664 5835 3680 5869
rect 3614 5801 3680 5835
rect 3614 5767 3630 5801
rect 3664 5767 3680 5801
rect 3614 5733 3680 5767
rect 3614 5699 3630 5733
rect 3664 5699 3680 5733
rect 3614 5665 3680 5699
rect 3614 5631 3630 5665
rect 3664 5631 3680 5665
rect 3614 5590 3680 5631
rect 3710 6549 3776 6590
rect 3710 6515 3726 6549
rect 3760 6515 3776 6549
rect 3710 6481 3776 6515
rect 3710 6447 3726 6481
rect 3760 6447 3776 6481
rect 3710 6413 3776 6447
rect 3710 6379 3726 6413
rect 3760 6379 3776 6413
rect 3710 6345 3776 6379
rect 3710 6311 3726 6345
rect 3760 6311 3776 6345
rect 3710 6277 3776 6311
rect 3710 6243 3726 6277
rect 3760 6243 3776 6277
rect 3710 6209 3776 6243
rect 3710 6175 3726 6209
rect 3760 6175 3776 6209
rect 3710 6141 3776 6175
rect 3710 6107 3726 6141
rect 3760 6107 3776 6141
rect 3710 6073 3776 6107
rect 3710 6039 3726 6073
rect 3760 6039 3776 6073
rect 3710 6005 3776 6039
rect 3710 5971 3726 6005
rect 3760 5971 3776 6005
rect 3710 5937 3776 5971
rect 3710 5903 3726 5937
rect 3760 5903 3776 5937
rect 3710 5869 3776 5903
rect 3710 5835 3726 5869
rect 3760 5835 3776 5869
rect 3710 5801 3776 5835
rect 3710 5767 3726 5801
rect 3760 5767 3776 5801
rect 3710 5733 3776 5767
rect 3710 5699 3726 5733
rect 3760 5699 3776 5733
rect 3710 5665 3776 5699
rect 3710 5631 3726 5665
rect 3760 5631 3776 5665
rect 3710 5590 3776 5631
rect 3806 6549 3872 6590
rect 3806 6515 3822 6549
rect 3856 6515 3872 6549
rect 3806 6481 3872 6515
rect 3806 6447 3822 6481
rect 3856 6447 3872 6481
rect 3806 6413 3872 6447
rect 3806 6379 3822 6413
rect 3856 6379 3872 6413
rect 3806 6345 3872 6379
rect 3806 6311 3822 6345
rect 3856 6311 3872 6345
rect 3806 6277 3872 6311
rect 3806 6243 3822 6277
rect 3856 6243 3872 6277
rect 3806 6209 3872 6243
rect 3806 6175 3822 6209
rect 3856 6175 3872 6209
rect 3806 6141 3872 6175
rect 3806 6107 3822 6141
rect 3856 6107 3872 6141
rect 3806 6073 3872 6107
rect 3806 6039 3822 6073
rect 3856 6039 3872 6073
rect 3806 6005 3872 6039
rect 3806 5971 3822 6005
rect 3856 5971 3872 6005
rect 3806 5937 3872 5971
rect 3806 5903 3822 5937
rect 3856 5903 3872 5937
rect 3806 5869 3872 5903
rect 3806 5835 3822 5869
rect 3856 5835 3872 5869
rect 3806 5801 3872 5835
rect 3806 5767 3822 5801
rect 3856 5767 3872 5801
rect 3806 5733 3872 5767
rect 3806 5699 3822 5733
rect 3856 5699 3872 5733
rect 3806 5665 3872 5699
rect 3806 5631 3822 5665
rect 3856 5631 3872 5665
rect 3806 5590 3872 5631
rect 3902 6549 3968 6590
rect 3902 6515 3918 6549
rect 3952 6515 3968 6549
rect 3902 6481 3968 6515
rect 3902 6447 3918 6481
rect 3952 6447 3968 6481
rect 3902 6413 3968 6447
rect 3902 6379 3918 6413
rect 3952 6379 3968 6413
rect 3902 6345 3968 6379
rect 3902 6311 3918 6345
rect 3952 6311 3968 6345
rect 3902 6277 3968 6311
rect 3902 6243 3918 6277
rect 3952 6243 3968 6277
rect 3902 6209 3968 6243
rect 3902 6175 3918 6209
rect 3952 6175 3968 6209
rect 3902 6141 3968 6175
rect 3902 6107 3918 6141
rect 3952 6107 3968 6141
rect 3902 6073 3968 6107
rect 3902 6039 3918 6073
rect 3952 6039 3968 6073
rect 3902 6005 3968 6039
rect 3902 5971 3918 6005
rect 3952 5971 3968 6005
rect 3902 5937 3968 5971
rect 3902 5903 3918 5937
rect 3952 5903 3968 5937
rect 3902 5869 3968 5903
rect 3902 5835 3918 5869
rect 3952 5835 3968 5869
rect 3902 5801 3968 5835
rect 3902 5767 3918 5801
rect 3952 5767 3968 5801
rect 3902 5733 3968 5767
rect 3902 5699 3918 5733
rect 3952 5699 3968 5733
rect 3902 5665 3968 5699
rect 3902 5631 3918 5665
rect 3952 5631 3968 5665
rect 3902 5590 3968 5631
rect 3998 6549 4064 6590
rect 3998 6515 4014 6549
rect 4048 6515 4064 6549
rect 3998 6481 4064 6515
rect 3998 6447 4014 6481
rect 4048 6447 4064 6481
rect 3998 6413 4064 6447
rect 3998 6379 4014 6413
rect 4048 6379 4064 6413
rect 3998 6345 4064 6379
rect 3998 6311 4014 6345
rect 4048 6311 4064 6345
rect 3998 6277 4064 6311
rect 3998 6243 4014 6277
rect 4048 6243 4064 6277
rect 3998 6209 4064 6243
rect 3998 6175 4014 6209
rect 4048 6175 4064 6209
rect 3998 6141 4064 6175
rect 3998 6107 4014 6141
rect 4048 6107 4064 6141
rect 3998 6073 4064 6107
rect 3998 6039 4014 6073
rect 4048 6039 4064 6073
rect 3998 6005 4064 6039
rect 3998 5971 4014 6005
rect 4048 5971 4064 6005
rect 3998 5937 4064 5971
rect 3998 5903 4014 5937
rect 4048 5903 4064 5937
rect 3998 5869 4064 5903
rect 3998 5835 4014 5869
rect 4048 5835 4064 5869
rect 3998 5801 4064 5835
rect 3998 5767 4014 5801
rect 4048 5767 4064 5801
rect 3998 5733 4064 5767
rect 3998 5699 4014 5733
rect 4048 5699 4064 5733
rect 3998 5665 4064 5699
rect 3998 5631 4014 5665
rect 4048 5631 4064 5665
rect 3998 5590 4064 5631
rect 4094 6549 4160 6590
rect 4094 6515 4110 6549
rect 4144 6515 4160 6549
rect 4094 6481 4160 6515
rect 4094 6447 4110 6481
rect 4144 6447 4160 6481
rect 4094 6413 4160 6447
rect 4094 6379 4110 6413
rect 4144 6379 4160 6413
rect 4094 6345 4160 6379
rect 4094 6311 4110 6345
rect 4144 6311 4160 6345
rect 4094 6277 4160 6311
rect 4094 6243 4110 6277
rect 4144 6243 4160 6277
rect 4094 6209 4160 6243
rect 4094 6175 4110 6209
rect 4144 6175 4160 6209
rect 4094 6141 4160 6175
rect 4094 6107 4110 6141
rect 4144 6107 4160 6141
rect 4094 6073 4160 6107
rect 4094 6039 4110 6073
rect 4144 6039 4160 6073
rect 4094 6005 4160 6039
rect 4094 5971 4110 6005
rect 4144 5971 4160 6005
rect 4094 5937 4160 5971
rect 4094 5903 4110 5937
rect 4144 5903 4160 5937
rect 4094 5869 4160 5903
rect 4094 5835 4110 5869
rect 4144 5835 4160 5869
rect 4094 5801 4160 5835
rect 4094 5767 4110 5801
rect 4144 5767 4160 5801
rect 4094 5733 4160 5767
rect 4094 5699 4110 5733
rect 4144 5699 4160 5733
rect 4094 5665 4160 5699
rect 4094 5631 4110 5665
rect 4144 5631 4160 5665
rect 4094 5590 4160 5631
rect 4190 6549 4256 6590
rect 4190 6515 4206 6549
rect 4240 6515 4256 6549
rect 4190 6481 4256 6515
rect 4190 6447 4206 6481
rect 4240 6447 4256 6481
rect 4190 6413 4256 6447
rect 4190 6379 4206 6413
rect 4240 6379 4256 6413
rect 4190 6345 4256 6379
rect 4190 6311 4206 6345
rect 4240 6311 4256 6345
rect 4190 6277 4256 6311
rect 4190 6243 4206 6277
rect 4240 6243 4256 6277
rect 4190 6209 4256 6243
rect 4190 6175 4206 6209
rect 4240 6175 4256 6209
rect 4190 6141 4256 6175
rect 4190 6107 4206 6141
rect 4240 6107 4256 6141
rect 4190 6073 4256 6107
rect 4190 6039 4206 6073
rect 4240 6039 4256 6073
rect 4190 6005 4256 6039
rect 4190 5971 4206 6005
rect 4240 5971 4256 6005
rect 4190 5937 4256 5971
rect 4190 5903 4206 5937
rect 4240 5903 4256 5937
rect 4190 5869 4256 5903
rect 4190 5835 4206 5869
rect 4240 5835 4256 5869
rect 4190 5801 4256 5835
rect 4190 5767 4206 5801
rect 4240 5767 4256 5801
rect 4190 5733 4256 5767
rect 4190 5699 4206 5733
rect 4240 5699 4256 5733
rect 4190 5665 4256 5699
rect 4190 5631 4206 5665
rect 4240 5631 4256 5665
rect 4190 5590 4256 5631
rect 4286 6549 4348 6590
rect 4286 6515 4302 6549
rect 4336 6515 4348 6549
rect 4286 6481 4348 6515
rect 4286 6447 4302 6481
rect 4336 6447 4348 6481
rect 4286 6413 4348 6447
rect 4286 6379 4302 6413
rect 4336 6379 4348 6413
rect 4286 6345 4348 6379
rect 4286 6311 4302 6345
rect 4336 6311 4348 6345
rect 4286 6277 4348 6311
rect 4286 6243 4302 6277
rect 4336 6243 4348 6277
rect 4286 6209 4348 6243
rect 4286 6175 4302 6209
rect 4336 6175 4348 6209
rect 4286 6141 4348 6175
rect 4286 6107 4302 6141
rect 4336 6107 4348 6141
rect 4286 6073 4348 6107
rect 4286 6039 4302 6073
rect 4336 6039 4348 6073
rect 4286 6005 4348 6039
rect 4286 5971 4302 6005
rect 4336 5971 4348 6005
rect 4286 5937 4348 5971
rect 4286 5903 4302 5937
rect 4336 5903 4348 5937
rect 4286 5869 4348 5903
rect 4286 5835 4302 5869
rect 4336 5835 4348 5869
rect 4286 5801 4348 5835
rect 4286 5767 4302 5801
rect 4336 5767 4348 5801
rect 4286 5733 4348 5767
rect 4286 5699 4302 5733
rect 4336 5699 4348 5733
rect 4286 5665 4348 5699
rect 4286 5631 4302 5665
rect 4336 5631 4348 5665
rect 4286 5590 4348 5631
rect 4904 6545 4966 6586
rect 4904 6511 4916 6545
rect 4950 6511 4966 6545
rect 4904 6477 4966 6511
rect 4904 6443 4916 6477
rect 4950 6443 4966 6477
rect 4904 6409 4966 6443
rect 4904 6375 4916 6409
rect 4950 6375 4966 6409
rect 4904 6341 4966 6375
rect 4904 6307 4916 6341
rect 4950 6307 4966 6341
rect 4904 6273 4966 6307
rect 4904 6239 4916 6273
rect 4950 6239 4966 6273
rect 4904 6205 4966 6239
rect 4904 6171 4916 6205
rect 4950 6171 4966 6205
rect 4904 6137 4966 6171
rect 4904 6103 4916 6137
rect 4950 6103 4966 6137
rect 4904 6069 4966 6103
rect 4904 6035 4916 6069
rect 4950 6035 4966 6069
rect 4904 6001 4966 6035
rect 4904 5967 4916 6001
rect 4950 5967 4966 6001
rect 4904 5933 4966 5967
rect 4904 5899 4916 5933
rect 4950 5899 4966 5933
rect 4904 5865 4966 5899
rect 4904 5831 4916 5865
rect 4950 5831 4966 5865
rect 4904 5797 4966 5831
rect 4904 5763 4916 5797
rect 4950 5763 4966 5797
rect 4904 5729 4966 5763
rect 4904 5695 4916 5729
rect 4950 5695 4966 5729
rect 4904 5661 4966 5695
rect 4904 5627 4916 5661
rect 4950 5627 4966 5661
rect 4904 5586 4966 5627
rect 4996 6545 5062 6586
rect 4996 6511 5012 6545
rect 5046 6511 5062 6545
rect 4996 6477 5062 6511
rect 4996 6443 5012 6477
rect 5046 6443 5062 6477
rect 4996 6409 5062 6443
rect 4996 6375 5012 6409
rect 5046 6375 5062 6409
rect 4996 6341 5062 6375
rect 4996 6307 5012 6341
rect 5046 6307 5062 6341
rect 4996 6273 5062 6307
rect 4996 6239 5012 6273
rect 5046 6239 5062 6273
rect 4996 6205 5062 6239
rect 4996 6171 5012 6205
rect 5046 6171 5062 6205
rect 4996 6137 5062 6171
rect 4996 6103 5012 6137
rect 5046 6103 5062 6137
rect 4996 6069 5062 6103
rect 4996 6035 5012 6069
rect 5046 6035 5062 6069
rect 4996 6001 5062 6035
rect 4996 5967 5012 6001
rect 5046 5967 5062 6001
rect 4996 5933 5062 5967
rect 4996 5899 5012 5933
rect 5046 5899 5062 5933
rect 4996 5865 5062 5899
rect 4996 5831 5012 5865
rect 5046 5831 5062 5865
rect 4996 5797 5062 5831
rect 4996 5763 5012 5797
rect 5046 5763 5062 5797
rect 4996 5729 5062 5763
rect 4996 5695 5012 5729
rect 5046 5695 5062 5729
rect 4996 5661 5062 5695
rect 4996 5627 5012 5661
rect 5046 5627 5062 5661
rect 4996 5586 5062 5627
rect 5092 6545 5158 6586
rect 5092 6511 5108 6545
rect 5142 6511 5158 6545
rect 5092 6477 5158 6511
rect 5092 6443 5108 6477
rect 5142 6443 5158 6477
rect 5092 6409 5158 6443
rect 5092 6375 5108 6409
rect 5142 6375 5158 6409
rect 5092 6341 5158 6375
rect 5092 6307 5108 6341
rect 5142 6307 5158 6341
rect 5092 6273 5158 6307
rect 5092 6239 5108 6273
rect 5142 6239 5158 6273
rect 5092 6205 5158 6239
rect 5092 6171 5108 6205
rect 5142 6171 5158 6205
rect 5092 6137 5158 6171
rect 5092 6103 5108 6137
rect 5142 6103 5158 6137
rect 5092 6069 5158 6103
rect 5092 6035 5108 6069
rect 5142 6035 5158 6069
rect 5092 6001 5158 6035
rect 5092 5967 5108 6001
rect 5142 5967 5158 6001
rect 5092 5933 5158 5967
rect 5092 5899 5108 5933
rect 5142 5899 5158 5933
rect 5092 5865 5158 5899
rect 5092 5831 5108 5865
rect 5142 5831 5158 5865
rect 5092 5797 5158 5831
rect 5092 5763 5108 5797
rect 5142 5763 5158 5797
rect 5092 5729 5158 5763
rect 5092 5695 5108 5729
rect 5142 5695 5158 5729
rect 5092 5661 5158 5695
rect 5092 5627 5108 5661
rect 5142 5627 5158 5661
rect 5092 5586 5158 5627
rect 5188 6545 5254 6586
rect 5188 6511 5204 6545
rect 5238 6511 5254 6545
rect 5188 6477 5254 6511
rect 5188 6443 5204 6477
rect 5238 6443 5254 6477
rect 5188 6409 5254 6443
rect 5188 6375 5204 6409
rect 5238 6375 5254 6409
rect 5188 6341 5254 6375
rect 5188 6307 5204 6341
rect 5238 6307 5254 6341
rect 5188 6273 5254 6307
rect 5188 6239 5204 6273
rect 5238 6239 5254 6273
rect 5188 6205 5254 6239
rect 5188 6171 5204 6205
rect 5238 6171 5254 6205
rect 5188 6137 5254 6171
rect 5188 6103 5204 6137
rect 5238 6103 5254 6137
rect 5188 6069 5254 6103
rect 5188 6035 5204 6069
rect 5238 6035 5254 6069
rect 5188 6001 5254 6035
rect 5188 5967 5204 6001
rect 5238 5967 5254 6001
rect 5188 5933 5254 5967
rect 5188 5899 5204 5933
rect 5238 5899 5254 5933
rect 5188 5865 5254 5899
rect 5188 5831 5204 5865
rect 5238 5831 5254 5865
rect 5188 5797 5254 5831
rect 5188 5763 5204 5797
rect 5238 5763 5254 5797
rect 5188 5729 5254 5763
rect 5188 5695 5204 5729
rect 5238 5695 5254 5729
rect 5188 5661 5254 5695
rect 5188 5627 5204 5661
rect 5238 5627 5254 5661
rect 5188 5586 5254 5627
rect 5284 6545 5350 6586
rect 5284 6511 5300 6545
rect 5334 6511 5350 6545
rect 5284 6477 5350 6511
rect 5284 6443 5300 6477
rect 5334 6443 5350 6477
rect 5284 6409 5350 6443
rect 5284 6375 5300 6409
rect 5334 6375 5350 6409
rect 5284 6341 5350 6375
rect 5284 6307 5300 6341
rect 5334 6307 5350 6341
rect 5284 6273 5350 6307
rect 5284 6239 5300 6273
rect 5334 6239 5350 6273
rect 5284 6205 5350 6239
rect 5284 6171 5300 6205
rect 5334 6171 5350 6205
rect 5284 6137 5350 6171
rect 5284 6103 5300 6137
rect 5334 6103 5350 6137
rect 5284 6069 5350 6103
rect 5284 6035 5300 6069
rect 5334 6035 5350 6069
rect 5284 6001 5350 6035
rect 5284 5967 5300 6001
rect 5334 5967 5350 6001
rect 5284 5933 5350 5967
rect 5284 5899 5300 5933
rect 5334 5899 5350 5933
rect 5284 5865 5350 5899
rect 5284 5831 5300 5865
rect 5334 5831 5350 5865
rect 5284 5797 5350 5831
rect 5284 5763 5300 5797
rect 5334 5763 5350 5797
rect 5284 5729 5350 5763
rect 5284 5695 5300 5729
rect 5334 5695 5350 5729
rect 5284 5661 5350 5695
rect 5284 5627 5300 5661
rect 5334 5627 5350 5661
rect 5284 5586 5350 5627
rect 5380 6545 5446 6586
rect 5380 6511 5396 6545
rect 5430 6511 5446 6545
rect 5380 6477 5446 6511
rect 5380 6443 5396 6477
rect 5430 6443 5446 6477
rect 5380 6409 5446 6443
rect 5380 6375 5396 6409
rect 5430 6375 5446 6409
rect 5380 6341 5446 6375
rect 5380 6307 5396 6341
rect 5430 6307 5446 6341
rect 5380 6273 5446 6307
rect 5380 6239 5396 6273
rect 5430 6239 5446 6273
rect 5380 6205 5446 6239
rect 5380 6171 5396 6205
rect 5430 6171 5446 6205
rect 5380 6137 5446 6171
rect 5380 6103 5396 6137
rect 5430 6103 5446 6137
rect 5380 6069 5446 6103
rect 5380 6035 5396 6069
rect 5430 6035 5446 6069
rect 5380 6001 5446 6035
rect 5380 5967 5396 6001
rect 5430 5967 5446 6001
rect 5380 5933 5446 5967
rect 5380 5899 5396 5933
rect 5430 5899 5446 5933
rect 5380 5865 5446 5899
rect 5380 5831 5396 5865
rect 5430 5831 5446 5865
rect 5380 5797 5446 5831
rect 5380 5763 5396 5797
rect 5430 5763 5446 5797
rect 5380 5729 5446 5763
rect 5380 5695 5396 5729
rect 5430 5695 5446 5729
rect 5380 5661 5446 5695
rect 5380 5627 5396 5661
rect 5430 5627 5446 5661
rect 5380 5586 5446 5627
rect 5476 6545 5542 6586
rect 5476 6511 5492 6545
rect 5526 6511 5542 6545
rect 5476 6477 5542 6511
rect 5476 6443 5492 6477
rect 5526 6443 5542 6477
rect 5476 6409 5542 6443
rect 5476 6375 5492 6409
rect 5526 6375 5542 6409
rect 5476 6341 5542 6375
rect 5476 6307 5492 6341
rect 5526 6307 5542 6341
rect 5476 6273 5542 6307
rect 5476 6239 5492 6273
rect 5526 6239 5542 6273
rect 5476 6205 5542 6239
rect 5476 6171 5492 6205
rect 5526 6171 5542 6205
rect 5476 6137 5542 6171
rect 5476 6103 5492 6137
rect 5526 6103 5542 6137
rect 5476 6069 5542 6103
rect 5476 6035 5492 6069
rect 5526 6035 5542 6069
rect 5476 6001 5542 6035
rect 5476 5967 5492 6001
rect 5526 5967 5542 6001
rect 5476 5933 5542 5967
rect 5476 5899 5492 5933
rect 5526 5899 5542 5933
rect 5476 5865 5542 5899
rect 5476 5831 5492 5865
rect 5526 5831 5542 5865
rect 5476 5797 5542 5831
rect 5476 5763 5492 5797
rect 5526 5763 5542 5797
rect 5476 5729 5542 5763
rect 5476 5695 5492 5729
rect 5526 5695 5542 5729
rect 5476 5661 5542 5695
rect 5476 5627 5492 5661
rect 5526 5627 5542 5661
rect 5476 5586 5542 5627
rect 5572 6545 5638 6586
rect 5572 6511 5588 6545
rect 5622 6511 5638 6545
rect 5572 6477 5638 6511
rect 5572 6443 5588 6477
rect 5622 6443 5638 6477
rect 5572 6409 5638 6443
rect 5572 6375 5588 6409
rect 5622 6375 5638 6409
rect 5572 6341 5638 6375
rect 5572 6307 5588 6341
rect 5622 6307 5638 6341
rect 5572 6273 5638 6307
rect 5572 6239 5588 6273
rect 5622 6239 5638 6273
rect 5572 6205 5638 6239
rect 5572 6171 5588 6205
rect 5622 6171 5638 6205
rect 5572 6137 5638 6171
rect 5572 6103 5588 6137
rect 5622 6103 5638 6137
rect 5572 6069 5638 6103
rect 5572 6035 5588 6069
rect 5622 6035 5638 6069
rect 5572 6001 5638 6035
rect 5572 5967 5588 6001
rect 5622 5967 5638 6001
rect 5572 5933 5638 5967
rect 5572 5899 5588 5933
rect 5622 5899 5638 5933
rect 5572 5865 5638 5899
rect 5572 5831 5588 5865
rect 5622 5831 5638 5865
rect 5572 5797 5638 5831
rect 5572 5763 5588 5797
rect 5622 5763 5638 5797
rect 5572 5729 5638 5763
rect 5572 5695 5588 5729
rect 5622 5695 5638 5729
rect 5572 5661 5638 5695
rect 5572 5627 5588 5661
rect 5622 5627 5638 5661
rect 5572 5586 5638 5627
rect 5668 6545 5730 6586
rect 5668 6511 5684 6545
rect 5718 6511 5730 6545
rect 5668 6477 5730 6511
rect 5668 6443 5684 6477
rect 5718 6443 5730 6477
rect 5668 6409 5730 6443
rect 5668 6375 5684 6409
rect 5718 6375 5730 6409
rect 5668 6341 5730 6375
rect 5668 6307 5684 6341
rect 5718 6307 5730 6341
rect 5668 6273 5730 6307
rect 5668 6239 5684 6273
rect 5718 6239 5730 6273
rect 5668 6205 5730 6239
rect 5668 6171 5684 6205
rect 5718 6171 5730 6205
rect 5668 6137 5730 6171
rect 5668 6103 5684 6137
rect 5718 6103 5730 6137
rect 5668 6069 5730 6103
rect 5668 6035 5684 6069
rect 5718 6035 5730 6069
rect 5668 6001 5730 6035
rect 5668 5967 5684 6001
rect 5718 5967 5730 6001
rect 5668 5933 5730 5967
rect 5668 5899 5684 5933
rect 5718 5899 5730 5933
rect 5668 5865 5730 5899
rect 5668 5831 5684 5865
rect 5718 5831 5730 5865
rect 5668 5797 5730 5831
rect 5668 5763 5684 5797
rect 5718 5763 5730 5797
rect 5668 5729 5730 5763
rect 5668 5695 5684 5729
rect 5718 5695 5730 5729
rect 5668 5661 5730 5695
rect 5668 5627 5684 5661
rect 5718 5627 5730 5661
rect 5668 5586 5730 5627
rect 6168 6549 6230 6590
rect 6168 6515 6180 6549
rect 6214 6515 6230 6549
rect 6168 6481 6230 6515
rect 6168 6447 6180 6481
rect 6214 6447 6230 6481
rect 6168 6413 6230 6447
rect 6168 6379 6180 6413
rect 6214 6379 6230 6413
rect 6168 6345 6230 6379
rect 6168 6311 6180 6345
rect 6214 6311 6230 6345
rect 6168 6277 6230 6311
rect 6168 6243 6180 6277
rect 6214 6243 6230 6277
rect 6168 6209 6230 6243
rect 6168 6175 6180 6209
rect 6214 6175 6230 6209
rect 6168 6141 6230 6175
rect 6168 6107 6180 6141
rect 6214 6107 6230 6141
rect 6168 6073 6230 6107
rect 6168 6039 6180 6073
rect 6214 6039 6230 6073
rect 6168 6005 6230 6039
rect 6168 5971 6180 6005
rect 6214 5971 6230 6005
rect 6168 5937 6230 5971
rect 6168 5903 6180 5937
rect 6214 5903 6230 5937
rect 6168 5869 6230 5903
rect 6168 5835 6180 5869
rect 6214 5835 6230 5869
rect 6168 5801 6230 5835
rect 6168 5767 6180 5801
rect 6214 5767 6230 5801
rect 6168 5733 6230 5767
rect 6168 5699 6180 5733
rect 6214 5699 6230 5733
rect 6168 5665 6230 5699
rect 6168 5631 6180 5665
rect 6214 5631 6230 5665
rect 6168 5590 6230 5631
rect 6260 6549 6326 6590
rect 6260 6515 6276 6549
rect 6310 6515 6326 6549
rect 6260 6481 6326 6515
rect 6260 6447 6276 6481
rect 6310 6447 6326 6481
rect 6260 6413 6326 6447
rect 6260 6379 6276 6413
rect 6310 6379 6326 6413
rect 6260 6345 6326 6379
rect 6260 6311 6276 6345
rect 6310 6311 6326 6345
rect 6260 6277 6326 6311
rect 6260 6243 6276 6277
rect 6310 6243 6326 6277
rect 6260 6209 6326 6243
rect 6260 6175 6276 6209
rect 6310 6175 6326 6209
rect 6260 6141 6326 6175
rect 6260 6107 6276 6141
rect 6310 6107 6326 6141
rect 6260 6073 6326 6107
rect 6260 6039 6276 6073
rect 6310 6039 6326 6073
rect 6260 6005 6326 6039
rect 6260 5971 6276 6005
rect 6310 5971 6326 6005
rect 6260 5937 6326 5971
rect 6260 5903 6276 5937
rect 6310 5903 6326 5937
rect 6260 5869 6326 5903
rect 6260 5835 6276 5869
rect 6310 5835 6326 5869
rect 6260 5801 6326 5835
rect 6260 5767 6276 5801
rect 6310 5767 6326 5801
rect 6260 5733 6326 5767
rect 6260 5699 6276 5733
rect 6310 5699 6326 5733
rect 6260 5665 6326 5699
rect 6260 5631 6276 5665
rect 6310 5631 6326 5665
rect 6260 5590 6326 5631
rect 6356 6549 6422 6590
rect 6356 6515 6372 6549
rect 6406 6515 6422 6549
rect 6356 6481 6422 6515
rect 6356 6447 6372 6481
rect 6406 6447 6422 6481
rect 6356 6413 6422 6447
rect 6356 6379 6372 6413
rect 6406 6379 6422 6413
rect 6356 6345 6422 6379
rect 6356 6311 6372 6345
rect 6406 6311 6422 6345
rect 6356 6277 6422 6311
rect 6356 6243 6372 6277
rect 6406 6243 6422 6277
rect 6356 6209 6422 6243
rect 6356 6175 6372 6209
rect 6406 6175 6422 6209
rect 6356 6141 6422 6175
rect 6356 6107 6372 6141
rect 6406 6107 6422 6141
rect 6356 6073 6422 6107
rect 6356 6039 6372 6073
rect 6406 6039 6422 6073
rect 6356 6005 6422 6039
rect 6356 5971 6372 6005
rect 6406 5971 6422 6005
rect 6356 5937 6422 5971
rect 6356 5903 6372 5937
rect 6406 5903 6422 5937
rect 6356 5869 6422 5903
rect 6356 5835 6372 5869
rect 6406 5835 6422 5869
rect 6356 5801 6422 5835
rect 6356 5767 6372 5801
rect 6406 5767 6422 5801
rect 6356 5733 6422 5767
rect 6356 5699 6372 5733
rect 6406 5699 6422 5733
rect 6356 5665 6422 5699
rect 6356 5631 6372 5665
rect 6406 5631 6422 5665
rect 6356 5590 6422 5631
rect 6452 6549 6518 6590
rect 6452 6515 6468 6549
rect 6502 6515 6518 6549
rect 6452 6481 6518 6515
rect 6452 6447 6468 6481
rect 6502 6447 6518 6481
rect 6452 6413 6518 6447
rect 6452 6379 6468 6413
rect 6502 6379 6518 6413
rect 6452 6345 6518 6379
rect 6452 6311 6468 6345
rect 6502 6311 6518 6345
rect 6452 6277 6518 6311
rect 6452 6243 6468 6277
rect 6502 6243 6518 6277
rect 6452 6209 6518 6243
rect 6452 6175 6468 6209
rect 6502 6175 6518 6209
rect 6452 6141 6518 6175
rect 6452 6107 6468 6141
rect 6502 6107 6518 6141
rect 6452 6073 6518 6107
rect 6452 6039 6468 6073
rect 6502 6039 6518 6073
rect 6452 6005 6518 6039
rect 6452 5971 6468 6005
rect 6502 5971 6518 6005
rect 6452 5937 6518 5971
rect 6452 5903 6468 5937
rect 6502 5903 6518 5937
rect 6452 5869 6518 5903
rect 6452 5835 6468 5869
rect 6502 5835 6518 5869
rect 6452 5801 6518 5835
rect 6452 5767 6468 5801
rect 6502 5767 6518 5801
rect 6452 5733 6518 5767
rect 6452 5699 6468 5733
rect 6502 5699 6518 5733
rect 6452 5665 6518 5699
rect 6452 5631 6468 5665
rect 6502 5631 6518 5665
rect 6452 5590 6518 5631
rect 6548 6549 6614 6590
rect 6548 6515 6564 6549
rect 6598 6515 6614 6549
rect 6548 6481 6614 6515
rect 6548 6447 6564 6481
rect 6598 6447 6614 6481
rect 6548 6413 6614 6447
rect 6548 6379 6564 6413
rect 6598 6379 6614 6413
rect 6548 6345 6614 6379
rect 6548 6311 6564 6345
rect 6598 6311 6614 6345
rect 6548 6277 6614 6311
rect 6548 6243 6564 6277
rect 6598 6243 6614 6277
rect 6548 6209 6614 6243
rect 6548 6175 6564 6209
rect 6598 6175 6614 6209
rect 6548 6141 6614 6175
rect 6548 6107 6564 6141
rect 6598 6107 6614 6141
rect 6548 6073 6614 6107
rect 6548 6039 6564 6073
rect 6598 6039 6614 6073
rect 6548 6005 6614 6039
rect 6548 5971 6564 6005
rect 6598 5971 6614 6005
rect 6548 5937 6614 5971
rect 6548 5903 6564 5937
rect 6598 5903 6614 5937
rect 6548 5869 6614 5903
rect 6548 5835 6564 5869
rect 6598 5835 6614 5869
rect 6548 5801 6614 5835
rect 6548 5767 6564 5801
rect 6598 5767 6614 5801
rect 6548 5733 6614 5767
rect 6548 5699 6564 5733
rect 6598 5699 6614 5733
rect 6548 5665 6614 5699
rect 6548 5631 6564 5665
rect 6598 5631 6614 5665
rect 6548 5590 6614 5631
rect 6644 6549 6710 6590
rect 6644 6515 6660 6549
rect 6694 6515 6710 6549
rect 6644 6481 6710 6515
rect 6644 6447 6660 6481
rect 6694 6447 6710 6481
rect 6644 6413 6710 6447
rect 6644 6379 6660 6413
rect 6694 6379 6710 6413
rect 6644 6345 6710 6379
rect 6644 6311 6660 6345
rect 6694 6311 6710 6345
rect 6644 6277 6710 6311
rect 6644 6243 6660 6277
rect 6694 6243 6710 6277
rect 6644 6209 6710 6243
rect 6644 6175 6660 6209
rect 6694 6175 6710 6209
rect 6644 6141 6710 6175
rect 6644 6107 6660 6141
rect 6694 6107 6710 6141
rect 6644 6073 6710 6107
rect 6644 6039 6660 6073
rect 6694 6039 6710 6073
rect 6644 6005 6710 6039
rect 6644 5971 6660 6005
rect 6694 5971 6710 6005
rect 6644 5937 6710 5971
rect 6644 5903 6660 5937
rect 6694 5903 6710 5937
rect 6644 5869 6710 5903
rect 6644 5835 6660 5869
rect 6694 5835 6710 5869
rect 6644 5801 6710 5835
rect 6644 5767 6660 5801
rect 6694 5767 6710 5801
rect 6644 5733 6710 5767
rect 6644 5699 6660 5733
rect 6694 5699 6710 5733
rect 6644 5665 6710 5699
rect 6644 5631 6660 5665
rect 6694 5631 6710 5665
rect 6644 5590 6710 5631
rect 6740 6549 6806 6590
rect 6740 6515 6756 6549
rect 6790 6515 6806 6549
rect 6740 6481 6806 6515
rect 6740 6447 6756 6481
rect 6790 6447 6806 6481
rect 6740 6413 6806 6447
rect 6740 6379 6756 6413
rect 6790 6379 6806 6413
rect 6740 6345 6806 6379
rect 6740 6311 6756 6345
rect 6790 6311 6806 6345
rect 6740 6277 6806 6311
rect 6740 6243 6756 6277
rect 6790 6243 6806 6277
rect 6740 6209 6806 6243
rect 6740 6175 6756 6209
rect 6790 6175 6806 6209
rect 6740 6141 6806 6175
rect 6740 6107 6756 6141
rect 6790 6107 6806 6141
rect 6740 6073 6806 6107
rect 6740 6039 6756 6073
rect 6790 6039 6806 6073
rect 6740 6005 6806 6039
rect 6740 5971 6756 6005
rect 6790 5971 6806 6005
rect 6740 5937 6806 5971
rect 6740 5903 6756 5937
rect 6790 5903 6806 5937
rect 6740 5869 6806 5903
rect 6740 5835 6756 5869
rect 6790 5835 6806 5869
rect 6740 5801 6806 5835
rect 6740 5767 6756 5801
rect 6790 5767 6806 5801
rect 6740 5733 6806 5767
rect 6740 5699 6756 5733
rect 6790 5699 6806 5733
rect 6740 5665 6806 5699
rect 6740 5631 6756 5665
rect 6790 5631 6806 5665
rect 6740 5590 6806 5631
rect 6836 6549 6902 6590
rect 6836 6515 6852 6549
rect 6886 6515 6902 6549
rect 6836 6481 6902 6515
rect 6836 6447 6852 6481
rect 6886 6447 6902 6481
rect 6836 6413 6902 6447
rect 6836 6379 6852 6413
rect 6886 6379 6902 6413
rect 6836 6345 6902 6379
rect 6836 6311 6852 6345
rect 6886 6311 6902 6345
rect 6836 6277 6902 6311
rect 6836 6243 6852 6277
rect 6886 6243 6902 6277
rect 6836 6209 6902 6243
rect 6836 6175 6852 6209
rect 6886 6175 6902 6209
rect 6836 6141 6902 6175
rect 6836 6107 6852 6141
rect 6886 6107 6902 6141
rect 6836 6073 6902 6107
rect 6836 6039 6852 6073
rect 6886 6039 6902 6073
rect 6836 6005 6902 6039
rect 6836 5971 6852 6005
rect 6886 5971 6902 6005
rect 6836 5937 6902 5971
rect 6836 5903 6852 5937
rect 6886 5903 6902 5937
rect 6836 5869 6902 5903
rect 6836 5835 6852 5869
rect 6886 5835 6902 5869
rect 6836 5801 6902 5835
rect 6836 5767 6852 5801
rect 6886 5767 6902 5801
rect 6836 5733 6902 5767
rect 6836 5699 6852 5733
rect 6886 5699 6902 5733
rect 6836 5665 6902 5699
rect 6836 5631 6852 5665
rect 6886 5631 6902 5665
rect 6836 5590 6902 5631
rect 6932 6549 6998 6590
rect 6932 6515 6948 6549
rect 6982 6515 6998 6549
rect 6932 6481 6998 6515
rect 6932 6447 6948 6481
rect 6982 6447 6998 6481
rect 6932 6413 6998 6447
rect 6932 6379 6948 6413
rect 6982 6379 6998 6413
rect 6932 6345 6998 6379
rect 6932 6311 6948 6345
rect 6982 6311 6998 6345
rect 6932 6277 6998 6311
rect 6932 6243 6948 6277
rect 6982 6243 6998 6277
rect 6932 6209 6998 6243
rect 6932 6175 6948 6209
rect 6982 6175 6998 6209
rect 6932 6141 6998 6175
rect 6932 6107 6948 6141
rect 6982 6107 6998 6141
rect 6932 6073 6998 6107
rect 6932 6039 6948 6073
rect 6982 6039 6998 6073
rect 6932 6005 6998 6039
rect 6932 5971 6948 6005
rect 6982 5971 6998 6005
rect 6932 5937 6998 5971
rect 6932 5903 6948 5937
rect 6982 5903 6998 5937
rect 6932 5869 6998 5903
rect 6932 5835 6948 5869
rect 6982 5835 6998 5869
rect 6932 5801 6998 5835
rect 6932 5767 6948 5801
rect 6982 5767 6998 5801
rect 6932 5733 6998 5767
rect 6932 5699 6948 5733
rect 6982 5699 6998 5733
rect 6932 5665 6998 5699
rect 6932 5631 6948 5665
rect 6982 5631 6998 5665
rect 6932 5590 6998 5631
rect 7028 6549 7094 6590
rect 7028 6515 7044 6549
rect 7078 6515 7094 6549
rect 7028 6481 7094 6515
rect 7028 6447 7044 6481
rect 7078 6447 7094 6481
rect 7028 6413 7094 6447
rect 7028 6379 7044 6413
rect 7078 6379 7094 6413
rect 7028 6345 7094 6379
rect 7028 6311 7044 6345
rect 7078 6311 7094 6345
rect 7028 6277 7094 6311
rect 7028 6243 7044 6277
rect 7078 6243 7094 6277
rect 7028 6209 7094 6243
rect 7028 6175 7044 6209
rect 7078 6175 7094 6209
rect 7028 6141 7094 6175
rect 7028 6107 7044 6141
rect 7078 6107 7094 6141
rect 7028 6073 7094 6107
rect 7028 6039 7044 6073
rect 7078 6039 7094 6073
rect 7028 6005 7094 6039
rect 7028 5971 7044 6005
rect 7078 5971 7094 6005
rect 7028 5937 7094 5971
rect 7028 5903 7044 5937
rect 7078 5903 7094 5937
rect 7028 5869 7094 5903
rect 7028 5835 7044 5869
rect 7078 5835 7094 5869
rect 7028 5801 7094 5835
rect 7028 5767 7044 5801
rect 7078 5767 7094 5801
rect 7028 5733 7094 5767
rect 7028 5699 7044 5733
rect 7078 5699 7094 5733
rect 7028 5665 7094 5699
rect 7028 5631 7044 5665
rect 7078 5631 7094 5665
rect 7028 5590 7094 5631
rect 7124 6549 7190 6590
rect 7124 6515 7140 6549
rect 7174 6515 7190 6549
rect 7124 6481 7190 6515
rect 7124 6447 7140 6481
rect 7174 6447 7190 6481
rect 7124 6413 7190 6447
rect 7124 6379 7140 6413
rect 7174 6379 7190 6413
rect 7124 6345 7190 6379
rect 7124 6311 7140 6345
rect 7174 6311 7190 6345
rect 7124 6277 7190 6311
rect 7124 6243 7140 6277
rect 7174 6243 7190 6277
rect 7124 6209 7190 6243
rect 7124 6175 7140 6209
rect 7174 6175 7190 6209
rect 7124 6141 7190 6175
rect 7124 6107 7140 6141
rect 7174 6107 7190 6141
rect 7124 6073 7190 6107
rect 7124 6039 7140 6073
rect 7174 6039 7190 6073
rect 7124 6005 7190 6039
rect 7124 5971 7140 6005
rect 7174 5971 7190 6005
rect 7124 5937 7190 5971
rect 7124 5903 7140 5937
rect 7174 5903 7190 5937
rect 7124 5869 7190 5903
rect 7124 5835 7140 5869
rect 7174 5835 7190 5869
rect 7124 5801 7190 5835
rect 7124 5767 7140 5801
rect 7174 5767 7190 5801
rect 7124 5733 7190 5767
rect 7124 5699 7140 5733
rect 7174 5699 7190 5733
rect 7124 5665 7190 5699
rect 7124 5631 7140 5665
rect 7174 5631 7190 5665
rect 7124 5590 7190 5631
rect 7220 6549 7286 6590
rect 7220 6515 7236 6549
rect 7270 6515 7286 6549
rect 7220 6481 7286 6515
rect 7220 6447 7236 6481
rect 7270 6447 7286 6481
rect 7220 6413 7286 6447
rect 7220 6379 7236 6413
rect 7270 6379 7286 6413
rect 7220 6345 7286 6379
rect 7220 6311 7236 6345
rect 7270 6311 7286 6345
rect 7220 6277 7286 6311
rect 7220 6243 7236 6277
rect 7270 6243 7286 6277
rect 7220 6209 7286 6243
rect 7220 6175 7236 6209
rect 7270 6175 7286 6209
rect 7220 6141 7286 6175
rect 7220 6107 7236 6141
rect 7270 6107 7286 6141
rect 7220 6073 7286 6107
rect 7220 6039 7236 6073
rect 7270 6039 7286 6073
rect 7220 6005 7286 6039
rect 7220 5971 7236 6005
rect 7270 5971 7286 6005
rect 7220 5937 7286 5971
rect 7220 5903 7236 5937
rect 7270 5903 7286 5937
rect 7220 5869 7286 5903
rect 7220 5835 7236 5869
rect 7270 5835 7286 5869
rect 7220 5801 7286 5835
rect 7220 5767 7236 5801
rect 7270 5767 7286 5801
rect 7220 5733 7286 5767
rect 7220 5699 7236 5733
rect 7270 5699 7286 5733
rect 7220 5665 7286 5699
rect 7220 5631 7236 5665
rect 7270 5631 7286 5665
rect 7220 5590 7286 5631
rect 7316 6549 7378 6590
rect 7316 6515 7332 6549
rect 7366 6515 7378 6549
rect 7316 6481 7378 6515
rect 7316 6447 7332 6481
rect 7366 6447 7378 6481
rect 7316 6413 7378 6447
rect 7316 6379 7332 6413
rect 7366 6379 7378 6413
rect 7316 6345 7378 6379
rect 7316 6311 7332 6345
rect 7366 6311 7378 6345
rect 7316 6277 7378 6311
rect 7316 6243 7332 6277
rect 7366 6243 7378 6277
rect 7316 6209 7378 6243
rect 7316 6175 7332 6209
rect 7366 6175 7378 6209
rect 7316 6141 7378 6175
rect 7316 6107 7332 6141
rect 7366 6107 7378 6141
rect 7316 6073 7378 6107
rect 7316 6039 7332 6073
rect 7366 6039 7378 6073
rect 7316 6005 7378 6039
rect 7316 5971 7332 6005
rect 7366 5971 7378 6005
rect 7316 5937 7378 5971
rect 7316 5903 7332 5937
rect 7366 5903 7378 5937
rect 7316 5869 7378 5903
rect 7316 5835 7332 5869
rect 7366 5835 7378 5869
rect 7316 5801 7378 5835
rect 7316 5767 7332 5801
rect 7366 5767 7378 5801
rect 7316 5733 7378 5767
rect 7316 5699 7332 5733
rect 7366 5699 7378 5733
rect 7316 5665 7378 5699
rect 7316 5631 7332 5665
rect 7366 5631 7378 5665
rect 7316 5590 7378 5631
rect 7934 6545 7996 6586
rect 7934 6511 7946 6545
rect 7980 6511 7996 6545
rect 7934 6477 7996 6511
rect 7934 6443 7946 6477
rect 7980 6443 7996 6477
rect 7934 6409 7996 6443
rect 7934 6375 7946 6409
rect 7980 6375 7996 6409
rect 7934 6341 7996 6375
rect 7934 6307 7946 6341
rect 7980 6307 7996 6341
rect 7934 6273 7996 6307
rect 7934 6239 7946 6273
rect 7980 6239 7996 6273
rect 7934 6205 7996 6239
rect 7934 6171 7946 6205
rect 7980 6171 7996 6205
rect 7934 6137 7996 6171
rect 7934 6103 7946 6137
rect 7980 6103 7996 6137
rect 7934 6069 7996 6103
rect 7934 6035 7946 6069
rect 7980 6035 7996 6069
rect 7934 6001 7996 6035
rect 7934 5967 7946 6001
rect 7980 5967 7996 6001
rect 7934 5933 7996 5967
rect 7934 5899 7946 5933
rect 7980 5899 7996 5933
rect 7934 5865 7996 5899
rect 7934 5831 7946 5865
rect 7980 5831 7996 5865
rect 7934 5797 7996 5831
rect 7934 5763 7946 5797
rect 7980 5763 7996 5797
rect 7934 5729 7996 5763
rect 7934 5695 7946 5729
rect 7980 5695 7996 5729
rect 7934 5661 7996 5695
rect 7934 5627 7946 5661
rect 7980 5627 7996 5661
rect 7934 5586 7996 5627
rect 8026 6545 8092 6586
rect 8026 6511 8042 6545
rect 8076 6511 8092 6545
rect 8026 6477 8092 6511
rect 8026 6443 8042 6477
rect 8076 6443 8092 6477
rect 8026 6409 8092 6443
rect 8026 6375 8042 6409
rect 8076 6375 8092 6409
rect 8026 6341 8092 6375
rect 8026 6307 8042 6341
rect 8076 6307 8092 6341
rect 8026 6273 8092 6307
rect 8026 6239 8042 6273
rect 8076 6239 8092 6273
rect 8026 6205 8092 6239
rect 8026 6171 8042 6205
rect 8076 6171 8092 6205
rect 8026 6137 8092 6171
rect 8026 6103 8042 6137
rect 8076 6103 8092 6137
rect 8026 6069 8092 6103
rect 8026 6035 8042 6069
rect 8076 6035 8092 6069
rect 8026 6001 8092 6035
rect 8026 5967 8042 6001
rect 8076 5967 8092 6001
rect 8026 5933 8092 5967
rect 8026 5899 8042 5933
rect 8076 5899 8092 5933
rect 8026 5865 8092 5899
rect 8026 5831 8042 5865
rect 8076 5831 8092 5865
rect 8026 5797 8092 5831
rect 8026 5763 8042 5797
rect 8076 5763 8092 5797
rect 8026 5729 8092 5763
rect 8026 5695 8042 5729
rect 8076 5695 8092 5729
rect 8026 5661 8092 5695
rect 8026 5627 8042 5661
rect 8076 5627 8092 5661
rect 8026 5586 8092 5627
rect 8122 6545 8188 6586
rect 8122 6511 8138 6545
rect 8172 6511 8188 6545
rect 8122 6477 8188 6511
rect 8122 6443 8138 6477
rect 8172 6443 8188 6477
rect 8122 6409 8188 6443
rect 8122 6375 8138 6409
rect 8172 6375 8188 6409
rect 8122 6341 8188 6375
rect 8122 6307 8138 6341
rect 8172 6307 8188 6341
rect 8122 6273 8188 6307
rect 8122 6239 8138 6273
rect 8172 6239 8188 6273
rect 8122 6205 8188 6239
rect 8122 6171 8138 6205
rect 8172 6171 8188 6205
rect 8122 6137 8188 6171
rect 8122 6103 8138 6137
rect 8172 6103 8188 6137
rect 8122 6069 8188 6103
rect 8122 6035 8138 6069
rect 8172 6035 8188 6069
rect 8122 6001 8188 6035
rect 8122 5967 8138 6001
rect 8172 5967 8188 6001
rect 8122 5933 8188 5967
rect 8122 5899 8138 5933
rect 8172 5899 8188 5933
rect 8122 5865 8188 5899
rect 8122 5831 8138 5865
rect 8172 5831 8188 5865
rect 8122 5797 8188 5831
rect 8122 5763 8138 5797
rect 8172 5763 8188 5797
rect 8122 5729 8188 5763
rect 8122 5695 8138 5729
rect 8172 5695 8188 5729
rect 8122 5661 8188 5695
rect 8122 5627 8138 5661
rect 8172 5627 8188 5661
rect 8122 5586 8188 5627
rect 8218 6545 8284 6586
rect 8218 6511 8234 6545
rect 8268 6511 8284 6545
rect 8218 6477 8284 6511
rect 8218 6443 8234 6477
rect 8268 6443 8284 6477
rect 8218 6409 8284 6443
rect 8218 6375 8234 6409
rect 8268 6375 8284 6409
rect 8218 6341 8284 6375
rect 8218 6307 8234 6341
rect 8268 6307 8284 6341
rect 8218 6273 8284 6307
rect 8218 6239 8234 6273
rect 8268 6239 8284 6273
rect 8218 6205 8284 6239
rect 8218 6171 8234 6205
rect 8268 6171 8284 6205
rect 8218 6137 8284 6171
rect 8218 6103 8234 6137
rect 8268 6103 8284 6137
rect 8218 6069 8284 6103
rect 8218 6035 8234 6069
rect 8268 6035 8284 6069
rect 8218 6001 8284 6035
rect 8218 5967 8234 6001
rect 8268 5967 8284 6001
rect 8218 5933 8284 5967
rect 8218 5899 8234 5933
rect 8268 5899 8284 5933
rect 8218 5865 8284 5899
rect 8218 5831 8234 5865
rect 8268 5831 8284 5865
rect 8218 5797 8284 5831
rect 8218 5763 8234 5797
rect 8268 5763 8284 5797
rect 8218 5729 8284 5763
rect 8218 5695 8234 5729
rect 8268 5695 8284 5729
rect 8218 5661 8284 5695
rect 8218 5627 8234 5661
rect 8268 5627 8284 5661
rect 8218 5586 8284 5627
rect 8314 6545 8380 6586
rect 8314 6511 8330 6545
rect 8364 6511 8380 6545
rect 8314 6477 8380 6511
rect 8314 6443 8330 6477
rect 8364 6443 8380 6477
rect 8314 6409 8380 6443
rect 8314 6375 8330 6409
rect 8364 6375 8380 6409
rect 8314 6341 8380 6375
rect 8314 6307 8330 6341
rect 8364 6307 8380 6341
rect 8314 6273 8380 6307
rect 8314 6239 8330 6273
rect 8364 6239 8380 6273
rect 8314 6205 8380 6239
rect 8314 6171 8330 6205
rect 8364 6171 8380 6205
rect 8314 6137 8380 6171
rect 8314 6103 8330 6137
rect 8364 6103 8380 6137
rect 8314 6069 8380 6103
rect 8314 6035 8330 6069
rect 8364 6035 8380 6069
rect 8314 6001 8380 6035
rect 8314 5967 8330 6001
rect 8364 5967 8380 6001
rect 8314 5933 8380 5967
rect 8314 5899 8330 5933
rect 8364 5899 8380 5933
rect 8314 5865 8380 5899
rect 8314 5831 8330 5865
rect 8364 5831 8380 5865
rect 8314 5797 8380 5831
rect 8314 5763 8330 5797
rect 8364 5763 8380 5797
rect 8314 5729 8380 5763
rect 8314 5695 8330 5729
rect 8364 5695 8380 5729
rect 8314 5661 8380 5695
rect 8314 5627 8330 5661
rect 8364 5627 8380 5661
rect 8314 5586 8380 5627
rect 8410 6545 8476 6586
rect 8410 6511 8426 6545
rect 8460 6511 8476 6545
rect 8410 6477 8476 6511
rect 8410 6443 8426 6477
rect 8460 6443 8476 6477
rect 8410 6409 8476 6443
rect 8410 6375 8426 6409
rect 8460 6375 8476 6409
rect 8410 6341 8476 6375
rect 8410 6307 8426 6341
rect 8460 6307 8476 6341
rect 8410 6273 8476 6307
rect 8410 6239 8426 6273
rect 8460 6239 8476 6273
rect 8410 6205 8476 6239
rect 8410 6171 8426 6205
rect 8460 6171 8476 6205
rect 8410 6137 8476 6171
rect 8410 6103 8426 6137
rect 8460 6103 8476 6137
rect 8410 6069 8476 6103
rect 8410 6035 8426 6069
rect 8460 6035 8476 6069
rect 8410 6001 8476 6035
rect 8410 5967 8426 6001
rect 8460 5967 8476 6001
rect 8410 5933 8476 5967
rect 8410 5899 8426 5933
rect 8460 5899 8476 5933
rect 8410 5865 8476 5899
rect 8410 5831 8426 5865
rect 8460 5831 8476 5865
rect 8410 5797 8476 5831
rect 8410 5763 8426 5797
rect 8460 5763 8476 5797
rect 8410 5729 8476 5763
rect 8410 5695 8426 5729
rect 8460 5695 8476 5729
rect 8410 5661 8476 5695
rect 8410 5627 8426 5661
rect 8460 5627 8476 5661
rect 8410 5586 8476 5627
rect 8506 6545 8572 6586
rect 8506 6511 8522 6545
rect 8556 6511 8572 6545
rect 8506 6477 8572 6511
rect 8506 6443 8522 6477
rect 8556 6443 8572 6477
rect 8506 6409 8572 6443
rect 8506 6375 8522 6409
rect 8556 6375 8572 6409
rect 8506 6341 8572 6375
rect 8506 6307 8522 6341
rect 8556 6307 8572 6341
rect 8506 6273 8572 6307
rect 8506 6239 8522 6273
rect 8556 6239 8572 6273
rect 8506 6205 8572 6239
rect 8506 6171 8522 6205
rect 8556 6171 8572 6205
rect 8506 6137 8572 6171
rect 8506 6103 8522 6137
rect 8556 6103 8572 6137
rect 8506 6069 8572 6103
rect 8506 6035 8522 6069
rect 8556 6035 8572 6069
rect 8506 6001 8572 6035
rect 8506 5967 8522 6001
rect 8556 5967 8572 6001
rect 8506 5933 8572 5967
rect 8506 5899 8522 5933
rect 8556 5899 8572 5933
rect 8506 5865 8572 5899
rect 8506 5831 8522 5865
rect 8556 5831 8572 5865
rect 8506 5797 8572 5831
rect 8506 5763 8522 5797
rect 8556 5763 8572 5797
rect 8506 5729 8572 5763
rect 8506 5695 8522 5729
rect 8556 5695 8572 5729
rect 8506 5661 8572 5695
rect 8506 5627 8522 5661
rect 8556 5627 8572 5661
rect 8506 5586 8572 5627
rect 8602 6545 8668 6586
rect 8602 6511 8618 6545
rect 8652 6511 8668 6545
rect 8602 6477 8668 6511
rect 8602 6443 8618 6477
rect 8652 6443 8668 6477
rect 8602 6409 8668 6443
rect 8602 6375 8618 6409
rect 8652 6375 8668 6409
rect 8602 6341 8668 6375
rect 8602 6307 8618 6341
rect 8652 6307 8668 6341
rect 8602 6273 8668 6307
rect 8602 6239 8618 6273
rect 8652 6239 8668 6273
rect 8602 6205 8668 6239
rect 8602 6171 8618 6205
rect 8652 6171 8668 6205
rect 8602 6137 8668 6171
rect 8602 6103 8618 6137
rect 8652 6103 8668 6137
rect 8602 6069 8668 6103
rect 8602 6035 8618 6069
rect 8652 6035 8668 6069
rect 8602 6001 8668 6035
rect 8602 5967 8618 6001
rect 8652 5967 8668 6001
rect 8602 5933 8668 5967
rect 8602 5899 8618 5933
rect 8652 5899 8668 5933
rect 8602 5865 8668 5899
rect 8602 5831 8618 5865
rect 8652 5831 8668 5865
rect 8602 5797 8668 5831
rect 8602 5763 8618 5797
rect 8652 5763 8668 5797
rect 8602 5729 8668 5763
rect 8602 5695 8618 5729
rect 8652 5695 8668 5729
rect 8602 5661 8668 5695
rect 8602 5627 8618 5661
rect 8652 5627 8668 5661
rect 8602 5586 8668 5627
rect 8698 6545 8760 6586
rect 8698 6511 8714 6545
rect 8748 6511 8760 6545
rect 8698 6477 8760 6511
rect 8698 6443 8714 6477
rect 8748 6443 8760 6477
rect 8698 6409 8760 6443
rect 8698 6375 8714 6409
rect 8748 6375 8760 6409
rect 8698 6341 8760 6375
rect 8698 6307 8714 6341
rect 8748 6307 8760 6341
rect 8698 6273 8760 6307
rect 8698 6239 8714 6273
rect 8748 6239 8760 6273
rect 8698 6205 8760 6239
rect 8698 6171 8714 6205
rect 8748 6171 8760 6205
rect 8698 6137 8760 6171
rect 8698 6103 8714 6137
rect 8748 6103 8760 6137
rect 8698 6069 8760 6103
rect 8698 6035 8714 6069
rect 8748 6035 8760 6069
rect 8698 6001 8760 6035
rect 8698 5967 8714 6001
rect 8748 5967 8760 6001
rect 8698 5933 8760 5967
rect 8698 5899 8714 5933
rect 8748 5899 8760 5933
rect 8698 5865 8760 5899
rect 8698 5831 8714 5865
rect 8748 5831 8760 5865
rect 8698 5797 8760 5831
rect 8698 5763 8714 5797
rect 8748 5763 8760 5797
rect 8698 5729 8760 5763
rect 8698 5695 8714 5729
rect 8748 5695 8760 5729
rect 8698 5661 8760 5695
rect 8698 5627 8714 5661
rect 8748 5627 8760 5661
rect 8698 5586 8760 5627
rect 9256 6547 9318 6588
rect 9256 6513 9268 6547
rect 9302 6513 9318 6547
rect 9256 6479 9318 6513
rect 9256 6445 9268 6479
rect 9302 6445 9318 6479
rect 9256 6411 9318 6445
rect 9256 6377 9268 6411
rect 9302 6377 9318 6411
rect 9256 6343 9318 6377
rect 9256 6309 9268 6343
rect 9302 6309 9318 6343
rect 9256 6275 9318 6309
rect 9256 6241 9268 6275
rect 9302 6241 9318 6275
rect 9256 6207 9318 6241
rect 9256 6173 9268 6207
rect 9302 6173 9318 6207
rect 9256 6139 9318 6173
rect 9256 6105 9268 6139
rect 9302 6105 9318 6139
rect 9256 6071 9318 6105
rect 9256 6037 9268 6071
rect 9302 6037 9318 6071
rect 9256 6003 9318 6037
rect 9256 5969 9268 6003
rect 9302 5969 9318 6003
rect 9256 5935 9318 5969
rect 9256 5901 9268 5935
rect 9302 5901 9318 5935
rect 9256 5867 9318 5901
rect 9256 5833 9268 5867
rect 9302 5833 9318 5867
rect 9256 5799 9318 5833
rect 9256 5765 9268 5799
rect 9302 5765 9318 5799
rect 9256 5731 9318 5765
rect 9256 5697 9268 5731
rect 9302 5697 9318 5731
rect 9256 5663 9318 5697
rect 9256 5629 9268 5663
rect 9302 5629 9318 5663
rect 9256 5588 9318 5629
rect 9348 6547 9414 6588
rect 9348 6513 9364 6547
rect 9398 6513 9414 6547
rect 9348 6479 9414 6513
rect 9348 6445 9364 6479
rect 9398 6445 9414 6479
rect 9348 6411 9414 6445
rect 9348 6377 9364 6411
rect 9398 6377 9414 6411
rect 9348 6343 9414 6377
rect 9348 6309 9364 6343
rect 9398 6309 9414 6343
rect 9348 6275 9414 6309
rect 9348 6241 9364 6275
rect 9398 6241 9414 6275
rect 9348 6207 9414 6241
rect 9348 6173 9364 6207
rect 9398 6173 9414 6207
rect 9348 6139 9414 6173
rect 9348 6105 9364 6139
rect 9398 6105 9414 6139
rect 9348 6071 9414 6105
rect 9348 6037 9364 6071
rect 9398 6037 9414 6071
rect 9348 6003 9414 6037
rect 9348 5969 9364 6003
rect 9398 5969 9414 6003
rect 9348 5935 9414 5969
rect 9348 5901 9364 5935
rect 9398 5901 9414 5935
rect 9348 5867 9414 5901
rect 9348 5833 9364 5867
rect 9398 5833 9414 5867
rect 9348 5799 9414 5833
rect 9348 5765 9364 5799
rect 9398 5765 9414 5799
rect 9348 5731 9414 5765
rect 9348 5697 9364 5731
rect 9398 5697 9414 5731
rect 9348 5663 9414 5697
rect 9348 5629 9364 5663
rect 9398 5629 9414 5663
rect 9348 5588 9414 5629
rect 9444 6547 9510 6588
rect 9444 6513 9460 6547
rect 9494 6513 9510 6547
rect 9444 6479 9510 6513
rect 9444 6445 9460 6479
rect 9494 6445 9510 6479
rect 9444 6411 9510 6445
rect 9444 6377 9460 6411
rect 9494 6377 9510 6411
rect 9444 6343 9510 6377
rect 9444 6309 9460 6343
rect 9494 6309 9510 6343
rect 9444 6275 9510 6309
rect 9444 6241 9460 6275
rect 9494 6241 9510 6275
rect 9444 6207 9510 6241
rect 9444 6173 9460 6207
rect 9494 6173 9510 6207
rect 9444 6139 9510 6173
rect 9444 6105 9460 6139
rect 9494 6105 9510 6139
rect 9444 6071 9510 6105
rect 9444 6037 9460 6071
rect 9494 6037 9510 6071
rect 9444 6003 9510 6037
rect 9444 5969 9460 6003
rect 9494 5969 9510 6003
rect 9444 5935 9510 5969
rect 9444 5901 9460 5935
rect 9494 5901 9510 5935
rect 9444 5867 9510 5901
rect 9444 5833 9460 5867
rect 9494 5833 9510 5867
rect 9444 5799 9510 5833
rect 9444 5765 9460 5799
rect 9494 5765 9510 5799
rect 9444 5731 9510 5765
rect 9444 5697 9460 5731
rect 9494 5697 9510 5731
rect 9444 5663 9510 5697
rect 9444 5629 9460 5663
rect 9494 5629 9510 5663
rect 9444 5588 9510 5629
rect 9540 6547 9606 6588
rect 9540 6513 9556 6547
rect 9590 6513 9606 6547
rect 9540 6479 9606 6513
rect 9540 6445 9556 6479
rect 9590 6445 9606 6479
rect 9540 6411 9606 6445
rect 9540 6377 9556 6411
rect 9590 6377 9606 6411
rect 9540 6343 9606 6377
rect 9540 6309 9556 6343
rect 9590 6309 9606 6343
rect 9540 6275 9606 6309
rect 9540 6241 9556 6275
rect 9590 6241 9606 6275
rect 9540 6207 9606 6241
rect 9540 6173 9556 6207
rect 9590 6173 9606 6207
rect 9540 6139 9606 6173
rect 9540 6105 9556 6139
rect 9590 6105 9606 6139
rect 9540 6071 9606 6105
rect 9540 6037 9556 6071
rect 9590 6037 9606 6071
rect 9540 6003 9606 6037
rect 9540 5969 9556 6003
rect 9590 5969 9606 6003
rect 9540 5935 9606 5969
rect 9540 5901 9556 5935
rect 9590 5901 9606 5935
rect 9540 5867 9606 5901
rect 9540 5833 9556 5867
rect 9590 5833 9606 5867
rect 9540 5799 9606 5833
rect 9540 5765 9556 5799
rect 9590 5765 9606 5799
rect 9540 5731 9606 5765
rect 9540 5697 9556 5731
rect 9590 5697 9606 5731
rect 9540 5663 9606 5697
rect 9540 5629 9556 5663
rect 9590 5629 9606 5663
rect 9540 5588 9606 5629
rect 9636 6547 9702 6588
rect 9636 6513 9652 6547
rect 9686 6513 9702 6547
rect 9636 6479 9702 6513
rect 9636 6445 9652 6479
rect 9686 6445 9702 6479
rect 9636 6411 9702 6445
rect 9636 6377 9652 6411
rect 9686 6377 9702 6411
rect 9636 6343 9702 6377
rect 9636 6309 9652 6343
rect 9686 6309 9702 6343
rect 9636 6275 9702 6309
rect 9636 6241 9652 6275
rect 9686 6241 9702 6275
rect 9636 6207 9702 6241
rect 9636 6173 9652 6207
rect 9686 6173 9702 6207
rect 9636 6139 9702 6173
rect 9636 6105 9652 6139
rect 9686 6105 9702 6139
rect 9636 6071 9702 6105
rect 9636 6037 9652 6071
rect 9686 6037 9702 6071
rect 9636 6003 9702 6037
rect 9636 5969 9652 6003
rect 9686 5969 9702 6003
rect 9636 5935 9702 5969
rect 9636 5901 9652 5935
rect 9686 5901 9702 5935
rect 9636 5867 9702 5901
rect 9636 5833 9652 5867
rect 9686 5833 9702 5867
rect 9636 5799 9702 5833
rect 9636 5765 9652 5799
rect 9686 5765 9702 5799
rect 9636 5731 9702 5765
rect 9636 5697 9652 5731
rect 9686 5697 9702 5731
rect 9636 5663 9702 5697
rect 9636 5629 9652 5663
rect 9686 5629 9702 5663
rect 9636 5588 9702 5629
rect 9732 6547 9798 6588
rect 9732 6513 9748 6547
rect 9782 6513 9798 6547
rect 9732 6479 9798 6513
rect 9732 6445 9748 6479
rect 9782 6445 9798 6479
rect 9732 6411 9798 6445
rect 9732 6377 9748 6411
rect 9782 6377 9798 6411
rect 9732 6343 9798 6377
rect 9732 6309 9748 6343
rect 9782 6309 9798 6343
rect 9732 6275 9798 6309
rect 9732 6241 9748 6275
rect 9782 6241 9798 6275
rect 9732 6207 9798 6241
rect 9732 6173 9748 6207
rect 9782 6173 9798 6207
rect 9732 6139 9798 6173
rect 9732 6105 9748 6139
rect 9782 6105 9798 6139
rect 9732 6071 9798 6105
rect 9732 6037 9748 6071
rect 9782 6037 9798 6071
rect 9732 6003 9798 6037
rect 9732 5969 9748 6003
rect 9782 5969 9798 6003
rect 9732 5935 9798 5969
rect 9732 5901 9748 5935
rect 9782 5901 9798 5935
rect 9732 5867 9798 5901
rect 9732 5833 9748 5867
rect 9782 5833 9798 5867
rect 9732 5799 9798 5833
rect 9732 5765 9748 5799
rect 9782 5765 9798 5799
rect 9732 5731 9798 5765
rect 9732 5697 9748 5731
rect 9782 5697 9798 5731
rect 9732 5663 9798 5697
rect 9732 5629 9748 5663
rect 9782 5629 9798 5663
rect 9732 5588 9798 5629
rect 9828 6547 9894 6588
rect 9828 6513 9844 6547
rect 9878 6513 9894 6547
rect 9828 6479 9894 6513
rect 9828 6445 9844 6479
rect 9878 6445 9894 6479
rect 9828 6411 9894 6445
rect 9828 6377 9844 6411
rect 9878 6377 9894 6411
rect 9828 6343 9894 6377
rect 9828 6309 9844 6343
rect 9878 6309 9894 6343
rect 9828 6275 9894 6309
rect 9828 6241 9844 6275
rect 9878 6241 9894 6275
rect 9828 6207 9894 6241
rect 9828 6173 9844 6207
rect 9878 6173 9894 6207
rect 9828 6139 9894 6173
rect 9828 6105 9844 6139
rect 9878 6105 9894 6139
rect 9828 6071 9894 6105
rect 9828 6037 9844 6071
rect 9878 6037 9894 6071
rect 9828 6003 9894 6037
rect 9828 5969 9844 6003
rect 9878 5969 9894 6003
rect 9828 5935 9894 5969
rect 9828 5901 9844 5935
rect 9878 5901 9894 5935
rect 9828 5867 9894 5901
rect 9828 5833 9844 5867
rect 9878 5833 9894 5867
rect 9828 5799 9894 5833
rect 9828 5765 9844 5799
rect 9878 5765 9894 5799
rect 9828 5731 9894 5765
rect 9828 5697 9844 5731
rect 9878 5697 9894 5731
rect 9828 5663 9894 5697
rect 9828 5629 9844 5663
rect 9878 5629 9894 5663
rect 9828 5588 9894 5629
rect 9924 6547 9990 6588
rect 9924 6513 9940 6547
rect 9974 6513 9990 6547
rect 9924 6479 9990 6513
rect 9924 6445 9940 6479
rect 9974 6445 9990 6479
rect 9924 6411 9990 6445
rect 9924 6377 9940 6411
rect 9974 6377 9990 6411
rect 9924 6343 9990 6377
rect 9924 6309 9940 6343
rect 9974 6309 9990 6343
rect 9924 6275 9990 6309
rect 9924 6241 9940 6275
rect 9974 6241 9990 6275
rect 9924 6207 9990 6241
rect 9924 6173 9940 6207
rect 9974 6173 9990 6207
rect 9924 6139 9990 6173
rect 9924 6105 9940 6139
rect 9974 6105 9990 6139
rect 9924 6071 9990 6105
rect 9924 6037 9940 6071
rect 9974 6037 9990 6071
rect 9924 6003 9990 6037
rect 9924 5969 9940 6003
rect 9974 5969 9990 6003
rect 9924 5935 9990 5969
rect 9924 5901 9940 5935
rect 9974 5901 9990 5935
rect 9924 5867 9990 5901
rect 9924 5833 9940 5867
rect 9974 5833 9990 5867
rect 9924 5799 9990 5833
rect 9924 5765 9940 5799
rect 9974 5765 9990 5799
rect 9924 5731 9990 5765
rect 9924 5697 9940 5731
rect 9974 5697 9990 5731
rect 9924 5663 9990 5697
rect 9924 5629 9940 5663
rect 9974 5629 9990 5663
rect 9924 5588 9990 5629
rect 10020 6547 10086 6588
rect 10020 6513 10036 6547
rect 10070 6513 10086 6547
rect 10020 6479 10086 6513
rect 10020 6445 10036 6479
rect 10070 6445 10086 6479
rect 10020 6411 10086 6445
rect 10020 6377 10036 6411
rect 10070 6377 10086 6411
rect 10020 6343 10086 6377
rect 10020 6309 10036 6343
rect 10070 6309 10086 6343
rect 10020 6275 10086 6309
rect 10020 6241 10036 6275
rect 10070 6241 10086 6275
rect 10020 6207 10086 6241
rect 10020 6173 10036 6207
rect 10070 6173 10086 6207
rect 10020 6139 10086 6173
rect 10020 6105 10036 6139
rect 10070 6105 10086 6139
rect 10020 6071 10086 6105
rect 10020 6037 10036 6071
rect 10070 6037 10086 6071
rect 10020 6003 10086 6037
rect 10020 5969 10036 6003
rect 10070 5969 10086 6003
rect 10020 5935 10086 5969
rect 10020 5901 10036 5935
rect 10070 5901 10086 5935
rect 10020 5867 10086 5901
rect 10020 5833 10036 5867
rect 10070 5833 10086 5867
rect 10020 5799 10086 5833
rect 10020 5765 10036 5799
rect 10070 5765 10086 5799
rect 10020 5731 10086 5765
rect 10020 5697 10036 5731
rect 10070 5697 10086 5731
rect 10020 5663 10086 5697
rect 10020 5629 10036 5663
rect 10070 5629 10086 5663
rect 10020 5588 10086 5629
rect 10116 6547 10182 6588
rect 10116 6513 10132 6547
rect 10166 6513 10182 6547
rect 10116 6479 10182 6513
rect 10116 6445 10132 6479
rect 10166 6445 10182 6479
rect 10116 6411 10182 6445
rect 10116 6377 10132 6411
rect 10166 6377 10182 6411
rect 10116 6343 10182 6377
rect 10116 6309 10132 6343
rect 10166 6309 10182 6343
rect 10116 6275 10182 6309
rect 10116 6241 10132 6275
rect 10166 6241 10182 6275
rect 10116 6207 10182 6241
rect 10116 6173 10132 6207
rect 10166 6173 10182 6207
rect 10116 6139 10182 6173
rect 10116 6105 10132 6139
rect 10166 6105 10182 6139
rect 10116 6071 10182 6105
rect 10116 6037 10132 6071
rect 10166 6037 10182 6071
rect 10116 6003 10182 6037
rect 10116 5969 10132 6003
rect 10166 5969 10182 6003
rect 10116 5935 10182 5969
rect 10116 5901 10132 5935
rect 10166 5901 10182 5935
rect 10116 5867 10182 5901
rect 10116 5833 10132 5867
rect 10166 5833 10182 5867
rect 10116 5799 10182 5833
rect 10116 5765 10132 5799
rect 10166 5765 10182 5799
rect 10116 5731 10182 5765
rect 10116 5697 10132 5731
rect 10166 5697 10182 5731
rect 10116 5663 10182 5697
rect 10116 5629 10132 5663
rect 10166 5629 10182 5663
rect 10116 5588 10182 5629
rect 10212 6547 10278 6588
rect 10212 6513 10228 6547
rect 10262 6513 10278 6547
rect 10212 6479 10278 6513
rect 10212 6445 10228 6479
rect 10262 6445 10278 6479
rect 10212 6411 10278 6445
rect 10212 6377 10228 6411
rect 10262 6377 10278 6411
rect 10212 6343 10278 6377
rect 10212 6309 10228 6343
rect 10262 6309 10278 6343
rect 10212 6275 10278 6309
rect 10212 6241 10228 6275
rect 10262 6241 10278 6275
rect 10212 6207 10278 6241
rect 10212 6173 10228 6207
rect 10262 6173 10278 6207
rect 10212 6139 10278 6173
rect 10212 6105 10228 6139
rect 10262 6105 10278 6139
rect 10212 6071 10278 6105
rect 10212 6037 10228 6071
rect 10262 6037 10278 6071
rect 10212 6003 10278 6037
rect 10212 5969 10228 6003
rect 10262 5969 10278 6003
rect 10212 5935 10278 5969
rect 10212 5901 10228 5935
rect 10262 5901 10278 5935
rect 10212 5867 10278 5901
rect 10212 5833 10228 5867
rect 10262 5833 10278 5867
rect 10212 5799 10278 5833
rect 10212 5765 10228 5799
rect 10262 5765 10278 5799
rect 10212 5731 10278 5765
rect 10212 5697 10228 5731
rect 10262 5697 10278 5731
rect 10212 5663 10278 5697
rect 10212 5629 10228 5663
rect 10262 5629 10278 5663
rect 10212 5588 10278 5629
rect 10308 6547 10374 6588
rect 10308 6513 10324 6547
rect 10358 6513 10374 6547
rect 10308 6479 10374 6513
rect 10308 6445 10324 6479
rect 10358 6445 10374 6479
rect 10308 6411 10374 6445
rect 10308 6377 10324 6411
rect 10358 6377 10374 6411
rect 10308 6343 10374 6377
rect 10308 6309 10324 6343
rect 10358 6309 10374 6343
rect 10308 6275 10374 6309
rect 10308 6241 10324 6275
rect 10358 6241 10374 6275
rect 10308 6207 10374 6241
rect 10308 6173 10324 6207
rect 10358 6173 10374 6207
rect 10308 6139 10374 6173
rect 10308 6105 10324 6139
rect 10358 6105 10374 6139
rect 10308 6071 10374 6105
rect 10308 6037 10324 6071
rect 10358 6037 10374 6071
rect 10308 6003 10374 6037
rect 10308 5969 10324 6003
rect 10358 5969 10374 6003
rect 10308 5935 10374 5969
rect 10308 5901 10324 5935
rect 10358 5901 10374 5935
rect 10308 5867 10374 5901
rect 10308 5833 10324 5867
rect 10358 5833 10374 5867
rect 10308 5799 10374 5833
rect 10308 5765 10324 5799
rect 10358 5765 10374 5799
rect 10308 5731 10374 5765
rect 10308 5697 10324 5731
rect 10358 5697 10374 5731
rect 10308 5663 10374 5697
rect 10308 5629 10324 5663
rect 10358 5629 10374 5663
rect 10308 5588 10374 5629
rect 10404 6547 10466 6588
rect 10404 6513 10420 6547
rect 10454 6513 10466 6547
rect 10404 6479 10466 6513
rect 10404 6445 10420 6479
rect 10454 6445 10466 6479
rect 10404 6411 10466 6445
rect 10404 6377 10420 6411
rect 10454 6377 10466 6411
rect 10404 6343 10466 6377
rect 10404 6309 10420 6343
rect 10454 6309 10466 6343
rect 10404 6275 10466 6309
rect 10404 6241 10420 6275
rect 10454 6241 10466 6275
rect 10404 6207 10466 6241
rect 10404 6173 10420 6207
rect 10454 6173 10466 6207
rect 10404 6139 10466 6173
rect 10404 6105 10420 6139
rect 10454 6105 10466 6139
rect 10404 6071 10466 6105
rect 10404 6037 10420 6071
rect 10454 6037 10466 6071
rect 10404 6003 10466 6037
rect 10404 5969 10420 6003
rect 10454 5969 10466 6003
rect 10404 5935 10466 5969
rect 10404 5901 10420 5935
rect 10454 5901 10466 5935
rect 10404 5867 10466 5901
rect 10404 5833 10420 5867
rect 10454 5833 10466 5867
rect 10404 5799 10466 5833
rect 10404 5765 10420 5799
rect 10454 5765 10466 5799
rect 10404 5731 10466 5765
rect 10404 5697 10420 5731
rect 10454 5697 10466 5731
rect 10404 5663 10466 5697
rect 10404 5629 10420 5663
rect 10454 5629 10466 5663
rect 10404 5588 10466 5629
rect 11022 6543 11084 6584
rect 11022 6509 11034 6543
rect 11068 6509 11084 6543
rect 11022 6475 11084 6509
rect 11022 6441 11034 6475
rect 11068 6441 11084 6475
rect 11022 6407 11084 6441
rect 11022 6373 11034 6407
rect 11068 6373 11084 6407
rect 11022 6339 11084 6373
rect 11022 6305 11034 6339
rect 11068 6305 11084 6339
rect 11022 6271 11084 6305
rect 11022 6237 11034 6271
rect 11068 6237 11084 6271
rect 11022 6203 11084 6237
rect 11022 6169 11034 6203
rect 11068 6169 11084 6203
rect 11022 6135 11084 6169
rect 11022 6101 11034 6135
rect 11068 6101 11084 6135
rect 11022 6067 11084 6101
rect 11022 6033 11034 6067
rect 11068 6033 11084 6067
rect 11022 5999 11084 6033
rect 11022 5965 11034 5999
rect 11068 5965 11084 5999
rect 11022 5931 11084 5965
rect 11022 5897 11034 5931
rect 11068 5897 11084 5931
rect 11022 5863 11084 5897
rect 11022 5829 11034 5863
rect 11068 5829 11084 5863
rect 11022 5795 11084 5829
rect 11022 5761 11034 5795
rect 11068 5761 11084 5795
rect 11022 5727 11084 5761
rect 11022 5693 11034 5727
rect 11068 5693 11084 5727
rect 11022 5659 11084 5693
rect 11022 5625 11034 5659
rect 11068 5625 11084 5659
rect 11022 5584 11084 5625
rect 11114 6543 11180 6584
rect 11114 6509 11130 6543
rect 11164 6509 11180 6543
rect 11114 6475 11180 6509
rect 11114 6441 11130 6475
rect 11164 6441 11180 6475
rect 11114 6407 11180 6441
rect 11114 6373 11130 6407
rect 11164 6373 11180 6407
rect 11114 6339 11180 6373
rect 11114 6305 11130 6339
rect 11164 6305 11180 6339
rect 11114 6271 11180 6305
rect 11114 6237 11130 6271
rect 11164 6237 11180 6271
rect 11114 6203 11180 6237
rect 11114 6169 11130 6203
rect 11164 6169 11180 6203
rect 11114 6135 11180 6169
rect 11114 6101 11130 6135
rect 11164 6101 11180 6135
rect 11114 6067 11180 6101
rect 11114 6033 11130 6067
rect 11164 6033 11180 6067
rect 11114 5999 11180 6033
rect 11114 5965 11130 5999
rect 11164 5965 11180 5999
rect 11114 5931 11180 5965
rect 11114 5897 11130 5931
rect 11164 5897 11180 5931
rect 11114 5863 11180 5897
rect 11114 5829 11130 5863
rect 11164 5829 11180 5863
rect 11114 5795 11180 5829
rect 11114 5761 11130 5795
rect 11164 5761 11180 5795
rect 11114 5727 11180 5761
rect 11114 5693 11130 5727
rect 11164 5693 11180 5727
rect 11114 5659 11180 5693
rect 11114 5625 11130 5659
rect 11164 5625 11180 5659
rect 11114 5584 11180 5625
rect 11210 6543 11276 6584
rect 11210 6509 11226 6543
rect 11260 6509 11276 6543
rect 11210 6475 11276 6509
rect 11210 6441 11226 6475
rect 11260 6441 11276 6475
rect 11210 6407 11276 6441
rect 11210 6373 11226 6407
rect 11260 6373 11276 6407
rect 11210 6339 11276 6373
rect 11210 6305 11226 6339
rect 11260 6305 11276 6339
rect 11210 6271 11276 6305
rect 11210 6237 11226 6271
rect 11260 6237 11276 6271
rect 11210 6203 11276 6237
rect 11210 6169 11226 6203
rect 11260 6169 11276 6203
rect 11210 6135 11276 6169
rect 11210 6101 11226 6135
rect 11260 6101 11276 6135
rect 11210 6067 11276 6101
rect 11210 6033 11226 6067
rect 11260 6033 11276 6067
rect 11210 5999 11276 6033
rect 11210 5965 11226 5999
rect 11260 5965 11276 5999
rect 11210 5931 11276 5965
rect 11210 5897 11226 5931
rect 11260 5897 11276 5931
rect 11210 5863 11276 5897
rect 11210 5829 11226 5863
rect 11260 5829 11276 5863
rect 11210 5795 11276 5829
rect 11210 5761 11226 5795
rect 11260 5761 11276 5795
rect 11210 5727 11276 5761
rect 11210 5693 11226 5727
rect 11260 5693 11276 5727
rect 11210 5659 11276 5693
rect 11210 5625 11226 5659
rect 11260 5625 11276 5659
rect 11210 5584 11276 5625
rect 11306 6543 11372 6584
rect 11306 6509 11322 6543
rect 11356 6509 11372 6543
rect 11306 6475 11372 6509
rect 11306 6441 11322 6475
rect 11356 6441 11372 6475
rect 11306 6407 11372 6441
rect 11306 6373 11322 6407
rect 11356 6373 11372 6407
rect 11306 6339 11372 6373
rect 11306 6305 11322 6339
rect 11356 6305 11372 6339
rect 11306 6271 11372 6305
rect 11306 6237 11322 6271
rect 11356 6237 11372 6271
rect 11306 6203 11372 6237
rect 11306 6169 11322 6203
rect 11356 6169 11372 6203
rect 11306 6135 11372 6169
rect 11306 6101 11322 6135
rect 11356 6101 11372 6135
rect 11306 6067 11372 6101
rect 11306 6033 11322 6067
rect 11356 6033 11372 6067
rect 11306 5999 11372 6033
rect 11306 5965 11322 5999
rect 11356 5965 11372 5999
rect 11306 5931 11372 5965
rect 11306 5897 11322 5931
rect 11356 5897 11372 5931
rect 11306 5863 11372 5897
rect 11306 5829 11322 5863
rect 11356 5829 11372 5863
rect 11306 5795 11372 5829
rect 11306 5761 11322 5795
rect 11356 5761 11372 5795
rect 11306 5727 11372 5761
rect 11306 5693 11322 5727
rect 11356 5693 11372 5727
rect 11306 5659 11372 5693
rect 11306 5625 11322 5659
rect 11356 5625 11372 5659
rect 11306 5584 11372 5625
rect 11402 6543 11468 6584
rect 11402 6509 11418 6543
rect 11452 6509 11468 6543
rect 11402 6475 11468 6509
rect 11402 6441 11418 6475
rect 11452 6441 11468 6475
rect 11402 6407 11468 6441
rect 11402 6373 11418 6407
rect 11452 6373 11468 6407
rect 11402 6339 11468 6373
rect 11402 6305 11418 6339
rect 11452 6305 11468 6339
rect 11402 6271 11468 6305
rect 11402 6237 11418 6271
rect 11452 6237 11468 6271
rect 11402 6203 11468 6237
rect 11402 6169 11418 6203
rect 11452 6169 11468 6203
rect 11402 6135 11468 6169
rect 11402 6101 11418 6135
rect 11452 6101 11468 6135
rect 11402 6067 11468 6101
rect 11402 6033 11418 6067
rect 11452 6033 11468 6067
rect 11402 5999 11468 6033
rect 11402 5965 11418 5999
rect 11452 5965 11468 5999
rect 11402 5931 11468 5965
rect 11402 5897 11418 5931
rect 11452 5897 11468 5931
rect 11402 5863 11468 5897
rect 11402 5829 11418 5863
rect 11452 5829 11468 5863
rect 11402 5795 11468 5829
rect 11402 5761 11418 5795
rect 11452 5761 11468 5795
rect 11402 5727 11468 5761
rect 11402 5693 11418 5727
rect 11452 5693 11468 5727
rect 11402 5659 11468 5693
rect 11402 5625 11418 5659
rect 11452 5625 11468 5659
rect 11402 5584 11468 5625
rect 11498 6543 11564 6584
rect 11498 6509 11514 6543
rect 11548 6509 11564 6543
rect 11498 6475 11564 6509
rect 11498 6441 11514 6475
rect 11548 6441 11564 6475
rect 11498 6407 11564 6441
rect 11498 6373 11514 6407
rect 11548 6373 11564 6407
rect 11498 6339 11564 6373
rect 11498 6305 11514 6339
rect 11548 6305 11564 6339
rect 11498 6271 11564 6305
rect 11498 6237 11514 6271
rect 11548 6237 11564 6271
rect 11498 6203 11564 6237
rect 11498 6169 11514 6203
rect 11548 6169 11564 6203
rect 11498 6135 11564 6169
rect 11498 6101 11514 6135
rect 11548 6101 11564 6135
rect 11498 6067 11564 6101
rect 11498 6033 11514 6067
rect 11548 6033 11564 6067
rect 11498 5999 11564 6033
rect 11498 5965 11514 5999
rect 11548 5965 11564 5999
rect 11498 5931 11564 5965
rect 11498 5897 11514 5931
rect 11548 5897 11564 5931
rect 11498 5863 11564 5897
rect 11498 5829 11514 5863
rect 11548 5829 11564 5863
rect 11498 5795 11564 5829
rect 11498 5761 11514 5795
rect 11548 5761 11564 5795
rect 11498 5727 11564 5761
rect 11498 5693 11514 5727
rect 11548 5693 11564 5727
rect 11498 5659 11564 5693
rect 11498 5625 11514 5659
rect 11548 5625 11564 5659
rect 11498 5584 11564 5625
rect 11594 6543 11660 6584
rect 11594 6509 11610 6543
rect 11644 6509 11660 6543
rect 11594 6475 11660 6509
rect 11594 6441 11610 6475
rect 11644 6441 11660 6475
rect 11594 6407 11660 6441
rect 11594 6373 11610 6407
rect 11644 6373 11660 6407
rect 11594 6339 11660 6373
rect 11594 6305 11610 6339
rect 11644 6305 11660 6339
rect 11594 6271 11660 6305
rect 11594 6237 11610 6271
rect 11644 6237 11660 6271
rect 11594 6203 11660 6237
rect 11594 6169 11610 6203
rect 11644 6169 11660 6203
rect 11594 6135 11660 6169
rect 11594 6101 11610 6135
rect 11644 6101 11660 6135
rect 11594 6067 11660 6101
rect 11594 6033 11610 6067
rect 11644 6033 11660 6067
rect 11594 5999 11660 6033
rect 11594 5965 11610 5999
rect 11644 5965 11660 5999
rect 11594 5931 11660 5965
rect 11594 5897 11610 5931
rect 11644 5897 11660 5931
rect 11594 5863 11660 5897
rect 11594 5829 11610 5863
rect 11644 5829 11660 5863
rect 11594 5795 11660 5829
rect 11594 5761 11610 5795
rect 11644 5761 11660 5795
rect 11594 5727 11660 5761
rect 11594 5693 11610 5727
rect 11644 5693 11660 5727
rect 11594 5659 11660 5693
rect 11594 5625 11610 5659
rect 11644 5625 11660 5659
rect 11594 5584 11660 5625
rect 11690 6543 11756 6584
rect 11690 6509 11706 6543
rect 11740 6509 11756 6543
rect 11690 6475 11756 6509
rect 11690 6441 11706 6475
rect 11740 6441 11756 6475
rect 11690 6407 11756 6441
rect 11690 6373 11706 6407
rect 11740 6373 11756 6407
rect 11690 6339 11756 6373
rect 11690 6305 11706 6339
rect 11740 6305 11756 6339
rect 11690 6271 11756 6305
rect 11690 6237 11706 6271
rect 11740 6237 11756 6271
rect 11690 6203 11756 6237
rect 11690 6169 11706 6203
rect 11740 6169 11756 6203
rect 11690 6135 11756 6169
rect 11690 6101 11706 6135
rect 11740 6101 11756 6135
rect 11690 6067 11756 6101
rect 11690 6033 11706 6067
rect 11740 6033 11756 6067
rect 11690 5999 11756 6033
rect 11690 5965 11706 5999
rect 11740 5965 11756 5999
rect 11690 5931 11756 5965
rect 11690 5897 11706 5931
rect 11740 5897 11756 5931
rect 11690 5863 11756 5897
rect 11690 5829 11706 5863
rect 11740 5829 11756 5863
rect 11690 5795 11756 5829
rect 11690 5761 11706 5795
rect 11740 5761 11756 5795
rect 11690 5727 11756 5761
rect 11690 5693 11706 5727
rect 11740 5693 11756 5727
rect 11690 5659 11756 5693
rect 11690 5625 11706 5659
rect 11740 5625 11756 5659
rect 11690 5584 11756 5625
rect 11786 6543 11848 6584
rect 11786 6509 11802 6543
rect 11836 6509 11848 6543
rect 11786 6475 11848 6509
rect 11786 6441 11802 6475
rect 11836 6441 11848 6475
rect 11786 6407 11848 6441
rect 11786 6373 11802 6407
rect 11836 6373 11848 6407
rect 11786 6339 11848 6373
rect 11786 6305 11802 6339
rect 11836 6305 11848 6339
rect 11786 6271 11848 6305
rect 11786 6237 11802 6271
rect 11836 6237 11848 6271
rect 11786 6203 11848 6237
rect 11786 6169 11802 6203
rect 11836 6169 11848 6203
rect 11786 6135 11848 6169
rect 11786 6101 11802 6135
rect 11836 6101 11848 6135
rect 11786 6067 11848 6101
rect 11786 6033 11802 6067
rect 11836 6033 11848 6067
rect 11786 5999 11848 6033
rect 11786 5965 11802 5999
rect 11836 5965 11848 5999
rect 11786 5931 11848 5965
rect 11786 5897 11802 5931
rect 11836 5897 11848 5931
rect 11786 5863 11848 5897
rect 11786 5829 11802 5863
rect 11836 5829 11848 5863
rect 11786 5795 11848 5829
rect 11786 5761 11802 5795
rect 11836 5761 11848 5795
rect 11786 5727 11848 5761
rect 11786 5693 11802 5727
rect 11836 5693 11848 5727
rect 11786 5659 11848 5693
rect 11786 5625 11802 5659
rect 11836 5625 11848 5659
rect 11786 5584 11848 5625
rect 12412 6521 12474 6562
rect 12412 6487 12424 6521
rect 12458 6487 12474 6521
rect 12412 6453 12474 6487
rect 12412 6419 12424 6453
rect 12458 6419 12474 6453
rect 12412 6385 12474 6419
rect 12412 6351 12424 6385
rect 12458 6351 12474 6385
rect 12412 6317 12474 6351
rect 12412 6283 12424 6317
rect 12458 6283 12474 6317
rect 12412 6249 12474 6283
rect 12412 6215 12424 6249
rect 12458 6215 12474 6249
rect 12412 6181 12474 6215
rect 12412 6147 12424 6181
rect 12458 6147 12474 6181
rect 12412 6113 12474 6147
rect 12412 6079 12424 6113
rect 12458 6079 12474 6113
rect 12412 6045 12474 6079
rect 12412 6011 12424 6045
rect 12458 6011 12474 6045
rect 12412 5977 12474 6011
rect 12412 5943 12424 5977
rect 12458 5943 12474 5977
rect 12412 5909 12474 5943
rect 12412 5875 12424 5909
rect 12458 5875 12474 5909
rect 12412 5841 12474 5875
rect 12412 5807 12424 5841
rect 12458 5807 12474 5841
rect 12412 5773 12474 5807
rect 12412 5739 12424 5773
rect 12458 5739 12474 5773
rect 12412 5705 12474 5739
rect 12412 5671 12424 5705
rect 12458 5671 12474 5705
rect 12412 5637 12474 5671
rect 12412 5603 12424 5637
rect 12458 5603 12474 5637
rect 12412 5562 12474 5603
rect 12504 6521 12570 6562
rect 12504 6487 12520 6521
rect 12554 6487 12570 6521
rect 12504 6453 12570 6487
rect 12504 6419 12520 6453
rect 12554 6419 12570 6453
rect 12504 6385 12570 6419
rect 12504 6351 12520 6385
rect 12554 6351 12570 6385
rect 12504 6317 12570 6351
rect 12504 6283 12520 6317
rect 12554 6283 12570 6317
rect 12504 6249 12570 6283
rect 12504 6215 12520 6249
rect 12554 6215 12570 6249
rect 12504 6181 12570 6215
rect 12504 6147 12520 6181
rect 12554 6147 12570 6181
rect 12504 6113 12570 6147
rect 12504 6079 12520 6113
rect 12554 6079 12570 6113
rect 12504 6045 12570 6079
rect 12504 6011 12520 6045
rect 12554 6011 12570 6045
rect 12504 5977 12570 6011
rect 12504 5943 12520 5977
rect 12554 5943 12570 5977
rect 12504 5909 12570 5943
rect 12504 5875 12520 5909
rect 12554 5875 12570 5909
rect 12504 5841 12570 5875
rect 12504 5807 12520 5841
rect 12554 5807 12570 5841
rect 12504 5773 12570 5807
rect 12504 5739 12520 5773
rect 12554 5739 12570 5773
rect 12504 5705 12570 5739
rect 12504 5671 12520 5705
rect 12554 5671 12570 5705
rect 12504 5637 12570 5671
rect 12504 5603 12520 5637
rect 12554 5603 12570 5637
rect 12504 5562 12570 5603
rect 12600 6521 12666 6562
rect 12600 6487 12616 6521
rect 12650 6487 12666 6521
rect 12600 6453 12666 6487
rect 12600 6419 12616 6453
rect 12650 6419 12666 6453
rect 12600 6385 12666 6419
rect 12600 6351 12616 6385
rect 12650 6351 12666 6385
rect 12600 6317 12666 6351
rect 12600 6283 12616 6317
rect 12650 6283 12666 6317
rect 12600 6249 12666 6283
rect 12600 6215 12616 6249
rect 12650 6215 12666 6249
rect 12600 6181 12666 6215
rect 12600 6147 12616 6181
rect 12650 6147 12666 6181
rect 12600 6113 12666 6147
rect 12600 6079 12616 6113
rect 12650 6079 12666 6113
rect 12600 6045 12666 6079
rect 12600 6011 12616 6045
rect 12650 6011 12666 6045
rect 12600 5977 12666 6011
rect 12600 5943 12616 5977
rect 12650 5943 12666 5977
rect 12600 5909 12666 5943
rect 12600 5875 12616 5909
rect 12650 5875 12666 5909
rect 12600 5841 12666 5875
rect 12600 5807 12616 5841
rect 12650 5807 12666 5841
rect 12600 5773 12666 5807
rect 12600 5739 12616 5773
rect 12650 5739 12666 5773
rect 12600 5705 12666 5739
rect 12600 5671 12616 5705
rect 12650 5671 12666 5705
rect 12600 5637 12666 5671
rect 12600 5603 12616 5637
rect 12650 5603 12666 5637
rect 12600 5562 12666 5603
rect 12696 6521 12762 6562
rect 12696 6487 12712 6521
rect 12746 6487 12762 6521
rect 12696 6453 12762 6487
rect 12696 6419 12712 6453
rect 12746 6419 12762 6453
rect 12696 6385 12762 6419
rect 12696 6351 12712 6385
rect 12746 6351 12762 6385
rect 12696 6317 12762 6351
rect 12696 6283 12712 6317
rect 12746 6283 12762 6317
rect 12696 6249 12762 6283
rect 12696 6215 12712 6249
rect 12746 6215 12762 6249
rect 12696 6181 12762 6215
rect 12696 6147 12712 6181
rect 12746 6147 12762 6181
rect 12696 6113 12762 6147
rect 12696 6079 12712 6113
rect 12746 6079 12762 6113
rect 12696 6045 12762 6079
rect 12696 6011 12712 6045
rect 12746 6011 12762 6045
rect 12696 5977 12762 6011
rect 12696 5943 12712 5977
rect 12746 5943 12762 5977
rect 12696 5909 12762 5943
rect 12696 5875 12712 5909
rect 12746 5875 12762 5909
rect 12696 5841 12762 5875
rect 12696 5807 12712 5841
rect 12746 5807 12762 5841
rect 12696 5773 12762 5807
rect 12696 5739 12712 5773
rect 12746 5739 12762 5773
rect 12696 5705 12762 5739
rect 12696 5671 12712 5705
rect 12746 5671 12762 5705
rect 12696 5637 12762 5671
rect 12696 5603 12712 5637
rect 12746 5603 12762 5637
rect 12696 5562 12762 5603
rect 12792 6521 12858 6562
rect 12792 6487 12808 6521
rect 12842 6487 12858 6521
rect 12792 6453 12858 6487
rect 12792 6419 12808 6453
rect 12842 6419 12858 6453
rect 12792 6385 12858 6419
rect 12792 6351 12808 6385
rect 12842 6351 12858 6385
rect 12792 6317 12858 6351
rect 12792 6283 12808 6317
rect 12842 6283 12858 6317
rect 12792 6249 12858 6283
rect 12792 6215 12808 6249
rect 12842 6215 12858 6249
rect 12792 6181 12858 6215
rect 12792 6147 12808 6181
rect 12842 6147 12858 6181
rect 12792 6113 12858 6147
rect 12792 6079 12808 6113
rect 12842 6079 12858 6113
rect 12792 6045 12858 6079
rect 12792 6011 12808 6045
rect 12842 6011 12858 6045
rect 12792 5977 12858 6011
rect 12792 5943 12808 5977
rect 12842 5943 12858 5977
rect 12792 5909 12858 5943
rect 12792 5875 12808 5909
rect 12842 5875 12858 5909
rect 12792 5841 12858 5875
rect 12792 5807 12808 5841
rect 12842 5807 12858 5841
rect 12792 5773 12858 5807
rect 12792 5739 12808 5773
rect 12842 5739 12858 5773
rect 12792 5705 12858 5739
rect 12792 5671 12808 5705
rect 12842 5671 12858 5705
rect 12792 5637 12858 5671
rect 12792 5603 12808 5637
rect 12842 5603 12858 5637
rect 12792 5562 12858 5603
rect 12888 6521 12954 6562
rect 12888 6487 12904 6521
rect 12938 6487 12954 6521
rect 12888 6453 12954 6487
rect 12888 6419 12904 6453
rect 12938 6419 12954 6453
rect 12888 6385 12954 6419
rect 12888 6351 12904 6385
rect 12938 6351 12954 6385
rect 12888 6317 12954 6351
rect 12888 6283 12904 6317
rect 12938 6283 12954 6317
rect 12888 6249 12954 6283
rect 12888 6215 12904 6249
rect 12938 6215 12954 6249
rect 12888 6181 12954 6215
rect 12888 6147 12904 6181
rect 12938 6147 12954 6181
rect 12888 6113 12954 6147
rect 12888 6079 12904 6113
rect 12938 6079 12954 6113
rect 12888 6045 12954 6079
rect 12888 6011 12904 6045
rect 12938 6011 12954 6045
rect 12888 5977 12954 6011
rect 12888 5943 12904 5977
rect 12938 5943 12954 5977
rect 12888 5909 12954 5943
rect 12888 5875 12904 5909
rect 12938 5875 12954 5909
rect 12888 5841 12954 5875
rect 12888 5807 12904 5841
rect 12938 5807 12954 5841
rect 12888 5773 12954 5807
rect 12888 5739 12904 5773
rect 12938 5739 12954 5773
rect 12888 5705 12954 5739
rect 12888 5671 12904 5705
rect 12938 5671 12954 5705
rect 12888 5637 12954 5671
rect 12888 5603 12904 5637
rect 12938 5603 12954 5637
rect 12888 5562 12954 5603
rect 12984 6521 13050 6562
rect 12984 6487 13000 6521
rect 13034 6487 13050 6521
rect 12984 6453 13050 6487
rect 12984 6419 13000 6453
rect 13034 6419 13050 6453
rect 12984 6385 13050 6419
rect 12984 6351 13000 6385
rect 13034 6351 13050 6385
rect 12984 6317 13050 6351
rect 12984 6283 13000 6317
rect 13034 6283 13050 6317
rect 12984 6249 13050 6283
rect 12984 6215 13000 6249
rect 13034 6215 13050 6249
rect 12984 6181 13050 6215
rect 12984 6147 13000 6181
rect 13034 6147 13050 6181
rect 12984 6113 13050 6147
rect 12984 6079 13000 6113
rect 13034 6079 13050 6113
rect 12984 6045 13050 6079
rect 12984 6011 13000 6045
rect 13034 6011 13050 6045
rect 12984 5977 13050 6011
rect 12984 5943 13000 5977
rect 13034 5943 13050 5977
rect 12984 5909 13050 5943
rect 12984 5875 13000 5909
rect 13034 5875 13050 5909
rect 12984 5841 13050 5875
rect 12984 5807 13000 5841
rect 13034 5807 13050 5841
rect 12984 5773 13050 5807
rect 12984 5739 13000 5773
rect 13034 5739 13050 5773
rect 12984 5705 13050 5739
rect 12984 5671 13000 5705
rect 13034 5671 13050 5705
rect 12984 5637 13050 5671
rect 12984 5603 13000 5637
rect 13034 5603 13050 5637
rect 12984 5562 13050 5603
rect 13080 6521 13146 6562
rect 13080 6487 13096 6521
rect 13130 6487 13146 6521
rect 13080 6453 13146 6487
rect 13080 6419 13096 6453
rect 13130 6419 13146 6453
rect 13080 6385 13146 6419
rect 13080 6351 13096 6385
rect 13130 6351 13146 6385
rect 13080 6317 13146 6351
rect 13080 6283 13096 6317
rect 13130 6283 13146 6317
rect 13080 6249 13146 6283
rect 13080 6215 13096 6249
rect 13130 6215 13146 6249
rect 13080 6181 13146 6215
rect 13080 6147 13096 6181
rect 13130 6147 13146 6181
rect 13080 6113 13146 6147
rect 13080 6079 13096 6113
rect 13130 6079 13146 6113
rect 13080 6045 13146 6079
rect 13080 6011 13096 6045
rect 13130 6011 13146 6045
rect 13080 5977 13146 6011
rect 13080 5943 13096 5977
rect 13130 5943 13146 5977
rect 13080 5909 13146 5943
rect 13080 5875 13096 5909
rect 13130 5875 13146 5909
rect 13080 5841 13146 5875
rect 13080 5807 13096 5841
rect 13130 5807 13146 5841
rect 13080 5773 13146 5807
rect 13080 5739 13096 5773
rect 13130 5739 13146 5773
rect 13080 5705 13146 5739
rect 13080 5671 13096 5705
rect 13130 5671 13146 5705
rect 13080 5637 13146 5671
rect 13080 5603 13096 5637
rect 13130 5603 13146 5637
rect 13080 5562 13146 5603
rect 13176 6521 13242 6562
rect 13176 6487 13192 6521
rect 13226 6487 13242 6521
rect 13176 6453 13242 6487
rect 13176 6419 13192 6453
rect 13226 6419 13242 6453
rect 13176 6385 13242 6419
rect 13176 6351 13192 6385
rect 13226 6351 13242 6385
rect 13176 6317 13242 6351
rect 13176 6283 13192 6317
rect 13226 6283 13242 6317
rect 13176 6249 13242 6283
rect 13176 6215 13192 6249
rect 13226 6215 13242 6249
rect 13176 6181 13242 6215
rect 13176 6147 13192 6181
rect 13226 6147 13242 6181
rect 13176 6113 13242 6147
rect 13176 6079 13192 6113
rect 13226 6079 13242 6113
rect 13176 6045 13242 6079
rect 13176 6011 13192 6045
rect 13226 6011 13242 6045
rect 13176 5977 13242 6011
rect 13176 5943 13192 5977
rect 13226 5943 13242 5977
rect 13176 5909 13242 5943
rect 13176 5875 13192 5909
rect 13226 5875 13242 5909
rect 13176 5841 13242 5875
rect 13176 5807 13192 5841
rect 13226 5807 13242 5841
rect 13176 5773 13242 5807
rect 13176 5739 13192 5773
rect 13226 5739 13242 5773
rect 13176 5705 13242 5739
rect 13176 5671 13192 5705
rect 13226 5671 13242 5705
rect 13176 5637 13242 5671
rect 13176 5603 13192 5637
rect 13226 5603 13242 5637
rect 13176 5562 13242 5603
rect 13272 6521 13338 6562
rect 13272 6487 13288 6521
rect 13322 6487 13338 6521
rect 13272 6453 13338 6487
rect 13272 6419 13288 6453
rect 13322 6419 13338 6453
rect 13272 6385 13338 6419
rect 13272 6351 13288 6385
rect 13322 6351 13338 6385
rect 13272 6317 13338 6351
rect 13272 6283 13288 6317
rect 13322 6283 13338 6317
rect 13272 6249 13338 6283
rect 13272 6215 13288 6249
rect 13322 6215 13338 6249
rect 13272 6181 13338 6215
rect 13272 6147 13288 6181
rect 13322 6147 13338 6181
rect 13272 6113 13338 6147
rect 13272 6079 13288 6113
rect 13322 6079 13338 6113
rect 13272 6045 13338 6079
rect 13272 6011 13288 6045
rect 13322 6011 13338 6045
rect 13272 5977 13338 6011
rect 13272 5943 13288 5977
rect 13322 5943 13338 5977
rect 13272 5909 13338 5943
rect 13272 5875 13288 5909
rect 13322 5875 13338 5909
rect 13272 5841 13338 5875
rect 13272 5807 13288 5841
rect 13322 5807 13338 5841
rect 13272 5773 13338 5807
rect 13272 5739 13288 5773
rect 13322 5739 13338 5773
rect 13272 5705 13338 5739
rect 13272 5671 13288 5705
rect 13322 5671 13338 5705
rect 13272 5637 13338 5671
rect 13272 5603 13288 5637
rect 13322 5603 13338 5637
rect 13272 5562 13338 5603
rect 13368 6521 13434 6562
rect 13368 6487 13384 6521
rect 13418 6487 13434 6521
rect 13368 6453 13434 6487
rect 13368 6419 13384 6453
rect 13418 6419 13434 6453
rect 13368 6385 13434 6419
rect 13368 6351 13384 6385
rect 13418 6351 13434 6385
rect 13368 6317 13434 6351
rect 13368 6283 13384 6317
rect 13418 6283 13434 6317
rect 13368 6249 13434 6283
rect 13368 6215 13384 6249
rect 13418 6215 13434 6249
rect 13368 6181 13434 6215
rect 13368 6147 13384 6181
rect 13418 6147 13434 6181
rect 13368 6113 13434 6147
rect 13368 6079 13384 6113
rect 13418 6079 13434 6113
rect 13368 6045 13434 6079
rect 13368 6011 13384 6045
rect 13418 6011 13434 6045
rect 13368 5977 13434 6011
rect 13368 5943 13384 5977
rect 13418 5943 13434 5977
rect 13368 5909 13434 5943
rect 13368 5875 13384 5909
rect 13418 5875 13434 5909
rect 13368 5841 13434 5875
rect 13368 5807 13384 5841
rect 13418 5807 13434 5841
rect 13368 5773 13434 5807
rect 13368 5739 13384 5773
rect 13418 5739 13434 5773
rect 13368 5705 13434 5739
rect 13368 5671 13384 5705
rect 13418 5671 13434 5705
rect 13368 5637 13434 5671
rect 13368 5603 13384 5637
rect 13418 5603 13434 5637
rect 13368 5562 13434 5603
rect 13464 6521 13530 6562
rect 13464 6487 13480 6521
rect 13514 6487 13530 6521
rect 13464 6453 13530 6487
rect 13464 6419 13480 6453
rect 13514 6419 13530 6453
rect 13464 6385 13530 6419
rect 13464 6351 13480 6385
rect 13514 6351 13530 6385
rect 13464 6317 13530 6351
rect 13464 6283 13480 6317
rect 13514 6283 13530 6317
rect 13464 6249 13530 6283
rect 13464 6215 13480 6249
rect 13514 6215 13530 6249
rect 13464 6181 13530 6215
rect 13464 6147 13480 6181
rect 13514 6147 13530 6181
rect 13464 6113 13530 6147
rect 13464 6079 13480 6113
rect 13514 6079 13530 6113
rect 13464 6045 13530 6079
rect 13464 6011 13480 6045
rect 13514 6011 13530 6045
rect 13464 5977 13530 6011
rect 13464 5943 13480 5977
rect 13514 5943 13530 5977
rect 13464 5909 13530 5943
rect 13464 5875 13480 5909
rect 13514 5875 13530 5909
rect 13464 5841 13530 5875
rect 13464 5807 13480 5841
rect 13514 5807 13530 5841
rect 13464 5773 13530 5807
rect 13464 5739 13480 5773
rect 13514 5739 13530 5773
rect 13464 5705 13530 5739
rect 13464 5671 13480 5705
rect 13514 5671 13530 5705
rect 13464 5637 13530 5671
rect 13464 5603 13480 5637
rect 13514 5603 13530 5637
rect 13464 5562 13530 5603
rect 13560 6521 13622 6562
rect 13560 6487 13576 6521
rect 13610 6487 13622 6521
rect 13560 6453 13622 6487
rect 13560 6419 13576 6453
rect 13610 6419 13622 6453
rect 13560 6385 13622 6419
rect 13560 6351 13576 6385
rect 13610 6351 13622 6385
rect 13560 6317 13622 6351
rect 13560 6283 13576 6317
rect 13610 6283 13622 6317
rect 13560 6249 13622 6283
rect 13560 6215 13576 6249
rect 13610 6215 13622 6249
rect 13560 6181 13622 6215
rect 13560 6147 13576 6181
rect 13610 6147 13622 6181
rect 13560 6113 13622 6147
rect 13560 6079 13576 6113
rect 13610 6079 13622 6113
rect 13560 6045 13622 6079
rect 13560 6011 13576 6045
rect 13610 6011 13622 6045
rect 13560 5977 13622 6011
rect 13560 5943 13576 5977
rect 13610 5943 13622 5977
rect 13560 5909 13622 5943
rect 13560 5875 13576 5909
rect 13610 5875 13622 5909
rect 13560 5841 13622 5875
rect 13560 5807 13576 5841
rect 13610 5807 13622 5841
rect 13560 5773 13622 5807
rect 13560 5739 13576 5773
rect 13610 5739 13622 5773
rect 13560 5705 13622 5739
rect 13560 5671 13576 5705
rect 13610 5671 13622 5705
rect 13560 5637 13622 5671
rect 13560 5603 13576 5637
rect 13610 5603 13622 5637
rect 13560 5562 13622 5603
rect 14178 6517 14240 6558
rect 14178 6483 14190 6517
rect 14224 6483 14240 6517
rect 14178 6449 14240 6483
rect 14178 6415 14190 6449
rect 14224 6415 14240 6449
rect 14178 6381 14240 6415
rect 14178 6347 14190 6381
rect 14224 6347 14240 6381
rect 14178 6313 14240 6347
rect 14178 6279 14190 6313
rect 14224 6279 14240 6313
rect 14178 6245 14240 6279
rect 14178 6211 14190 6245
rect 14224 6211 14240 6245
rect 14178 6177 14240 6211
rect 14178 6143 14190 6177
rect 14224 6143 14240 6177
rect 14178 6109 14240 6143
rect 14178 6075 14190 6109
rect 14224 6075 14240 6109
rect 14178 6041 14240 6075
rect 14178 6007 14190 6041
rect 14224 6007 14240 6041
rect 14178 5973 14240 6007
rect 14178 5939 14190 5973
rect 14224 5939 14240 5973
rect 14178 5905 14240 5939
rect 14178 5871 14190 5905
rect 14224 5871 14240 5905
rect 14178 5837 14240 5871
rect 14178 5803 14190 5837
rect 14224 5803 14240 5837
rect 14178 5769 14240 5803
rect 14178 5735 14190 5769
rect 14224 5735 14240 5769
rect 14178 5701 14240 5735
rect 14178 5667 14190 5701
rect 14224 5667 14240 5701
rect 14178 5633 14240 5667
rect 14178 5599 14190 5633
rect 14224 5599 14240 5633
rect -880 5521 -868 5555
rect -834 5521 -822 5555
rect 14178 5558 14240 5599
rect 14270 6517 14336 6558
rect 14270 6483 14286 6517
rect 14320 6483 14336 6517
rect 14270 6449 14336 6483
rect 14270 6415 14286 6449
rect 14320 6415 14336 6449
rect 14270 6381 14336 6415
rect 14270 6347 14286 6381
rect 14320 6347 14336 6381
rect 14270 6313 14336 6347
rect 14270 6279 14286 6313
rect 14320 6279 14336 6313
rect 14270 6245 14336 6279
rect 14270 6211 14286 6245
rect 14320 6211 14336 6245
rect 14270 6177 14336 6211
rect 14270 6143 14286 6177
rect 14320 6143 14336 6177
rect 14270 6109 14336 6143
rect 14270 6075 14286 6109
rect 14320 6075 14336 6109
rect 14270 6041 14336 6075
rect 14270 6007 14286 6041
rect 14320 6007 14336 6041
rect 14270 5973 14336 6007
rect 14270 5939 14286 5973
rect 14320 5939 14336 5973
rect 14270 5905 14336 5939
rect 14270 5871 14286 5905
rect 14320 5871 14336 5905
rect 14270 5837 14336 5871
rect 14270 5803 14286 5837
rect 14320 5803 14336 5837
rect 14270 5769 14336 5803
rect 14270 5735 14286 5769
rect 14320 5735 14336 5769
rect 14270 5701 14336 5735
rect 14270 5667 14286 5701
rect 14320 5667 14336 5701
rect 14270 5633 14336 5667
rect 14270 5599 14286 5633
rect 14320 5599 14336 5633
rect 14270 5558 14336 5599
rect 14366 6517 14432 6558
rect 14366 6483 14382 6517
rect 14416 6483 14432 6517
rect 14366 6449 14432 6483
rect 14366 6415 14382 6449
rect 14416 6415 14432 6449
rect 14366 6381 14432 6415
rect 14366 6347 14382 6381
rect 14416 6347 14432 6381
rect 14366 6313 14432 6347
rect 14366 6279 14382 6313
rect 14416 6279 14432 6313
rect 14366 6245 14432 6279
rect 14366 6211 14382 6245
rect 14416 6211 14432 6245
rect 14366 6177 14432 6211
rect 14366 6143 14382 6177
rect 14416 6143 14432 6177
rect 14366 6109 14432 6143
rect 14366 6075 14382 6109
rect 14416 6075 14432 6109
rect 14366 6041 14432 6075
rect 14366 6007 14382 6041
rect 14416 6007 14432 6041
rect 14366 5973 14432 6007
rect 14366 5939 14382 5973
rect 14416 5939 14432 5973
rect 14366 5905 14432 5939
rect 14366 5871 14382 5905
rect 14416 5871 14432 5905
rect 14366 5837 14432 5871
rect 14366 5803 14382 5837
rect 14416 5803 14432 5837
rect 14366 5769 14432 5803
rect 14366 5735 14382 5769
rect 14416 5735 14432 5769
rect 14366 5701 14432 5735
rect 14366 5667 14382 5701
rect 14416 5667 14432 5701
rect 14366 5633 14432 5667
rect 14366 5599 14382 5633
rect 14416 5599 14432 5633
rect 14366 5558 14432 5599
rect 14462 6517 14528 6558
rect 14462 6483 14478 6517
rect 14512 6483 14528 6517
rect 14462 6449 14528 6483
rect 14462 6415 14478 6449
rect 14512 6415 14528 6449
rect 14462 6381 14528 6415
rect 14462 6347 14478 6381
rect 14512 6347 14528 6381
rect 14462 6313 14528 6347
rect 14462 6279 14478 6313
rect 14512 6279 14528 6313
rect 14462 6245 14528 6279
rect 14462 6211 14478 6245
rect 14512 6211 14528 6245
rect 14462 6177 14528 6211
rect 14462 6143 14478 6177
rect 14512 6143 14528 6177
rect 14462 6109 14528 6143
rect 14462 6075 14478 6109
rect 14512 6075 14528 6109
rect 14462 6041 14528 6075
rect 14462 6007 14478 6041
rect 14512 6007 14528 6041
rect 14462 5973 14528 6007
rect 14462 5939 14478 5973
rect 14512 5939 14528 5973
rect 14462 5905 14528 5939
rect 14462 5871 14478 5905
rect 14512 5871 14528 5905
rect 14462 5837 14528 5871
rect 14462 5803 14478 5837
rect 14512 5803 14528 5837
rect 14462 5769 14528 5803
rect 14462 5735 14478 5769
rect 14512 5735 14528 5769
rect 14462 5701 14528 5735
rect 14462 5667 14478 5701
rect 14512 5667 14528 5701
rect 14462 5633 14528 5667
rect 14462 5599 14478 5633
rect 14512 5599 14528 5633
rect 14462 5558 14528 5599
rect 14558 6517 14624 6558
rect 14558 6483 14574 6517
rect 14608 6483 14624 6517
rect 14558 6449 14624 6483
rect 14558 6415 14574 6449
rect 14608 6415 14624 6449
rect 14558 6381 14624 6415
rect 14558 6347 14574 6381
rect 14608 6347 14624 6381
rect 14558 6313 14624 6347
rect 14558 6279 14574 6313
rect 14608 6279 14624 6313
rect 14558 6245 14624 6279
rect 14558 6211 14574 6245
rect 14608 6211 14624 6245
rect 14558 6177 14624 6211
rect 14558 6143 14574 6177
rect 14608 6143 14624 6177
rect 14558 6109 14624 6143
rect 14558 6075 14574 6109
rect 14608 6075 14624 6109
rect 14558 6041 14624 6075
rect 14558 6007 14574 6041
rect 14608 6007 14624 6041
rect 14558 5973 14624 6007
rect 14558 5939 14574 5973
rect 14608 5939 14624 5973
rect 14558 5905 14624 5939
rect 14558 5871 14574 5905
rect 14608 5871 14624 5905
rect 14558 5837 14624 5871
rect 14558 5803 14574 5837
rect 14608 5803 14624 5837
rect 14558 5769 14624 5803
rect 14558 5735 14574 5769
rect 14608 5735 14624 5769
rect 14558 5701 14624 5735
rect 14558 5667 14574 5701
rect 14608 5667 14624 5701
rect 14558 5633 14624 5667
rect 14558 5599 14574 5633
rect 14608 5599 14624 5633
rect 14558 5558 14624 5599
rect 14654 6517 14720 6558
rect 14654 6483 14670 6517
rect 14704 6483 14720 6517
rect 14654 6449 14720 6483
rect 14654 6415 14670 6449
rect 14704 6415 14720 6449
rect 14654 6381 14720 6415
rect 14654 6347 14670 6381
rect 14704 6347 14720 6381
rect 14654 6313 14720 6347
rect 14654 6279 14670 6313
rect 14704 6279 14720 6313
rect 14654 6245 14720 6279
rect 14654 6211 14670 6245
rect 14704 6211 14720 6245
rect 14654 6177 14720 6211
rect 14654 6143 14670 6177
rect 14704 6143 14720 6177
rect 14654 6109 14720 6143
rect 14654 6075 14670 6109
rect 14704 6075 14720 6109
rect 14654 6041 14720 6075
rect 14654 6007 14670 6041
rect 14704 6007 14720 6041
rect 14654 5973 14720 6007
rect 14654 5939 14670 5973
rect 14704 5939 14720 5973
rect 14654 5905 14720 5939
rect 14654 5871 14670 5905
rect 14704 5871 14720 5905
rect 14654 5837 14720 5871
rect 14654 5803 14670 5837
rect 14704 5803 14720 5837
rect 14654 5769 14720 5803
rect 14654 5735 14670 5769
rect 14704 5735 14720 5769
rect 14654 5701 14720 5735
rect 14654 5667 14670 5701
rect 14704 5667 14720 5701
rect 14654 5633 14720 5667
rect 14654 5599 14670 5633
rect 14704 5599 14720 5633
rect 14654 5558 14720 5599
rect 14750 6517 14816 6558
rect 14750 6483 14766 6517
rect 14800 6483 14816 6517
rect 14750 6449 14816 6483
rect 14750 6415 14766 6449
rect 14800 6415 14816 6449
rect 14750 6381 14816 6415
rect 14750 6347 14766 6381
rect 14800 6347 14816 6381
rect 14750 6313 14816 6347
rect 14750 6279 14766 6313
rect 14800 6279 14816 6313
rect 14750 6245 14816 6279
rect 14750 6211 14766 6245
rect 14800 6211 14816 6245
rect 14750 6177 14816 6211
rect 14750 6143 14766 6177
rect 14800 6143 14816 6177
rect 14750 6109 14816 6143
rect 14750 6075 14766 6109
rect 14800 6075 14816 6109
rect 14750 6041 14816 6075
rect 14750 6007 14766 6041
rect 14800 6007 14816 6041
rect 14750 5973 14816 6007
rect 14750 5939 14766 5973
rect 14800 5939 14816 5973
rect 14750 5905 14816 5939
rect 14750 5871 14766 5905
rect 14800 5871 14816 5905
rect 14750 5837 14816 5871
rect 14750 5803 14766 5837
rect 14800 5803 14816 5837
rect 14750 5769 14816 5803
rect 14750 5735 14766 5769
rect 14800 5735 14816 5769
rect 14750 5701 14816 5735
rect 14750 5667 14766 5701
rect 14800 5667 14816 5701
rect 14750 5633 14816 5667
rect 14750 5599 14766 5633
rect 14800 5599 14816 5633
rect 14750 5558 14816 5599
rect 14846 6517 14912 6558
rect 14846 6483 14862 6517
rect 14896 6483 14912 6517
rect 14846 6449 14912 6483
rect 14846 6415 14862 6449
rect 14896 6415 14912 6449
rect 14846 6381 14912 6415
rect 14846 6347 14862 6381
rect 14896 6347 14912 6381
rect 14846 6313 14912 6347
rect 14846 6279 14862 6313
rect 14896 6279 14912 6313
rect 14846 6245 14912 6279
rect 14846 6211 14862 6245
rect 14896 6211 14912 6245
rect 14846 6177 14912 6211
rect 14846 6143 14862 6177
rect 14896 6143 14912 6177
rect 14846 6109 14912 6143
rect 14846 6075 14862 6109
rect 14896 6075 14912 6109
rect 14846 6041 14912 6075
rect 14846 6007 14862 6041
rect 14896 6007 14912 6041
rect 14846 5973 14912 6007
rect 14846 5939 14862 5973
rect 14896 5939 14912 5973
rect 14846 5905 14912 5939
rect 14846 5871 14862 5905
rect 14896 5871 14912 5905
rect 14846 5837 14912 5871
rect 14846 5803 14862 5837
rect 14896 5803 14912 5837
rect 14846 5769 14912 5803
rect 14846 5735 14862 5769
rect 14896 5735 14912 5769
rect 14846 5701 14912 5735
rect 14846 5667 14862 5701
rect 14896 5667 14912 5701
rect 14846 5633 14912 5667
rect 14846 5599 14862 5633
rect 14896 5599 14912 5633
rect 14846 5558 14912 5599
rect 14942 6517 15004 6558
rect 14942 6483 14958 6517
rect 14992 6483 15004 6517
rect 14942 6449 15004 6483
rect 14942 6415 14958 6449
rect 14992 6415 15004 6449
rect 14942 6381 15004 6415
rect 14942 6347 14958 6381
rect 14992 6347 15004 6381
rect 14942 6313 15004 6347
rect 14942 6279 14958 6313
rect 14992 6279 15004 6313
rect 14942 6245 15004 6279
rect 14942 6211 14958 6245
rect 14992 6211 15004 6245
rect 14942 6177 15004 6211
rect 14942 6143 14958 6177
rect 14992 6143 15004 6177
rect 14942 6109 15004 6143
rect 14942 6075 14958 6109
rect 14992 6075 15004 6109
rect 14942 6041 15004 6075
rect 14942 6007 14958 6041
rect 14992 6007 15004 6041
rect 14942 5973 15004 6007
rect 14942 5939 14958 5973
rect 14992 5939 15004 5973
rect 14942 5905 15004 5939
rect 14942 5871 14958 5905
rect 14992 5871 15004 5905
rect 14942 5837 15004 5871
rect 14942 5803 14958 5837
rect 14992 5803 15004 5837
rect 14942 5769 15004 5803
rect 14942 5735 14958 5769
rect 14992 5735 15004 5769
rect 14942 5701 15004 5735
rect 14942 5667 14958 5701
rect 14992 5667 15004 5701
rect 14942 5633 15004 5667
rect 14942 5599 14958 5633
rect 14992 5599 15004 5633
rect 14942 5558 15004 5599
rect 15506 5895 15568 5926
rect 15506 5861 15518 5895
rect 15552 5861 15568 5895
rect 15506 5827 15568 5861
rect 15506 5793 15518 5827
rect 15552 5793 15568 5827
rect 15506 5759 15568 5793
rect 15506 5725 15518 5759
rect 15552 5725 15568 5759
rect 15506 5691 15568 5725
rect 15506 5657 15518 5691
rect 15552 5657 15568 5691
rect 15506 5623 15568 5657
rect 15506 5589 15518 5623
rect 15552 5589 15568 5623
rect 15506 5555 15568 5589
rect -880 5487 -822 5521
rect -880 5453 -868 5487
rect -834 5453 -822 5487
rect -880 5419 -822 5453
rect -880 5385 -868 5419
rect -834 5385 -822 5419
rect -880 5351 -822 5385
rect -880 5317 -868 5351
rect -834 5317 -822 5351
rect -880 5283 -822 5317
rect -880 5249 -868 5283
rect -834 5249 -822 5283
rect -880 5215 -822 5249
rect -880 5181 -868 5215
rect -834 5181 -822 5215
rect -880 5147 -822 5181
rect -880 5113 -868 5147
rect -834 5113 -822 5147
rect -880 5079 -822 5113
rect -880 5045 -868 5079
rect -834 5045 -822 5079
rect -880 5011 -822 5045
rect 15506 5521 15518 5555
rect 15552 5521 15568 5555
rect 15506 5487 15568 5521
rect 15506 5453 15518 5487
rect 15552 5453 15568 5487
rect 15506 5419 15568 5453
rect 15506 5385 15518 5419
rect 15552 5385 15568 5419
rect 15506 5351 15568 5385
rect 15506 5317 15518 5351
rect 15552 5317 15568 5351
rect 15506 5283 15568 5317
rect 15506 5249 15518 5283
rect 15552 5249 15568 5283
rect 15506 5215 15568 5249
rect 15506 5181 15518 5215
rect 15552 5181 15568 5215
rect 15506 5147 15568 5181
rect 15506 5113 15518 5147
rect 15552 5113 15568 5147
rect 15506 5079 15568 5113
rect 15506 5045 15518 5079
rect 15552 5045 15568 5079
rect -880 4977 -868 5011
rect -834 4977 -822 5011
rect -880 4936 -822 4977
rect 15506 5011 15568 5045
rect 1472 4903 1534 4944
rect 1472 4869 1484 4903
rect 1518 4869 1534 4903
rect 1472 4835 1534 4869
rect 1472 4801 1484 4835
rect 1518 4801 1534 4835
rect 1472 4767 1534 4801
rect 1472 4733 1484 4767
rect 1518 4733 1534 4767
rect 1472 4699 1534 4733
rect 1472 4665 1484 4699
rect 1518 4665 1534 4699
rect 1472 4631 1534 4665
rect 1472 4597 1484 4631
rect 1518 4597 1534 4631
rect 1472 4563 1534 4597
rect 1472 4529 1484 4563
rect 1518 4529 1534 4563
rect -23598 4401 -23536 4442
rect -23598 4367 -23586 4401
rect -23552 4367 -23536 4401
rect -23598 4333 -23536 4367
rect -23598 4299 -23586 4333
rect -23552 4299 -23536 4333
rect -23598 4265 -23536 4299
rect -23598 4231 -23586 4265
rect -23552 4231 -23536 4265
rect -23598 4197 -23536 4231
rect -23598 4163 -23586 4197
rect -23552 4163 -23536 4197
rect -23598 4129 -23536 4163
rect -23598 4095 -23586 4129
rect -23552 4095 -23536 4129
rect -23598 4061 -23536 4095
rect -23598 4027 -23586 4061
rect -23552 4027 -23536 4061
rect -23598 3993 -23536 4027
rect -23598 3959 -23586 3993
rect -23552 3959 -23536 3993
rect -23598 3925 -23536 3959
rect -23598 3891 -23586 3925
rect -23552 3891 -23536 3925
rect -23598 3857 -23536 3891
rect -23598 3823 -23586 3857
rect -23552 3823 -23536 3857
rect -23598 3789 -23536 3823
rect -23598 3755 -23586 3789
rect -23552 3755 -23536 3789
rect -23598 3721 -23536 3755
rect -23598 3687 -23586 3721
rect -23552 3687 -23536 3721
rect -23598 3653 -23536 3687
rect -23598 3619 -23586 3653
rect -23552 3619 -23536 3653
rect -23598 3585 -23536 3619
rect -23598 3551 -23586 3585
rect -23552 3551 -23536 3585
rect -23598 3517 -23536 3551
rect -23598 3483 -23586 3517
rect -23552 3483 -23536 3517
rect -23598 3442 -23536 3483
rect -23506 4401 -23440 4442
rect -23506 4367 -23490 4401
rect -23456 4367 -23440 4401
rect -23506 4333 -23440 4367
rect -23506 4299 -23490 4333
rect -23456 4299 -23440 4333
rect -23506 4265 -23440 4299
rect -23506 4231 -23490 4265
rect -23456 4231 -23440 4265
rect -23506 4197 -23440 4231
rect -23506 4163 -23490 4197
rect -23456 4163 -23440 4197
rect -23506 4129 -23440 4163
rect -23506 4095 -23490 4129
rect -23456 4095 -23440 4129
rect -23506 4061 -23440 4095
rect -23506 4027 -23490 4061
rect -23456 4027 -23440 4061
rect -23506 3993 -23440 4027
rect -23506 3959 -23490 3993
rect -23456 3959 -23440 3993
rect -23506 3925 -23440 3959
rect -23506 3891 -23490 3925
rect -23456 3891 -23440 3925
rect -23506 3857 -23440 3891
rect -23506 3823 -23490 3857
rect -23456 3823 -23440 3857
rect -23506 3789 -23440 3823
rect -23506 3755 -23490 3789
rect -23456 3755 -23440 3789
rect -23506 3721 -23440 3755
rect -23506 3687 -23490 3721
rect -23456 3687 -23440 3721
rect -23506 3653 -23440 3687
rect -23506 3619 -23490 3653
rect -23456 3619 -23440 3653
rect -23506 3585 -23440 3619
rect -23506 3551 -23490 3585
rect -23456 3551 -23440 3585
rect -23506 3517 -23440 3551
rect -23506 3483 -23490 3517
rect -23456 3483 -23440 3517
rect -23506 3442 -23440 3483
rect -23410 4401 -23344 4442
rect -23410 4367 -23394 4401
rect -23360 4367 -23344 4401
rect -23410 4333 -23344 4367
rect -23410 4299 -23394 4333
rect -23360 4299 -23344 4333
rect -23410 4265 -23344 4299
rect -23410 4231 -23394 4265
rect -23360 4231 -23344 4265
rect -23410 4197 -23344 4231
rect -23410 4163 -23394 4197
rect -23360 4163 -23344 4197
rect -23410 4129 -23344 4163
rect -23410 4095 -23394 4129
rect -23360 4095 -23344 4129
rect -23410 4061 -23344 4095
rect -23410 4027 -23394 4061
rect -23360 4027 -23344 4061
rect -23410 3993 -23344 4027
rect -23410 3959 -23394 3993
rect -23360 3959 -23344 3993
rect -23410 3925 -23344 3959
rect -23410 3891 -23394 3925
rect -23360 3891 -23344 3925
rect -23410 3857 -23344 3891
rect -23410 3823 -23394 3857
rect -23360 3823 -23344 3857
rect -23410 3789 -23344 3823
rect -23410 3755 -23394 3789
rect -23360 3755 -23344 3789
rect -23410 3721 -23344 3755
rect -23410 3687 -23394 3721
rect -23360 3687 -23344 3721
rect -23410 3653 -23344 3687
rect -23410 3619 -23394 3653
rect -23360 3619 -23344 3653
rect -23410 3585 -23344 3619
rect -23410 3551 -23394 3585
rect -23360 3551 -23344 3585
rect -23410 3517 -23344 3551
rect -23410 3483 -23394 3517
rect -23360 3483 -23344 3517
rect -23410 3442 -23344 3483
rect -23314 4401 -23248 4442
rect -23314 4367 -23298 4401
rect -23264 4367 -23248 4401
rect -23314 4333 -23248 4367
rect -23314 4299 -23298 4333
rect -23264 4299 -23248 4333
rect -23314 4265 -23248 4299
rect -23314 4231 -23298 4265
rect -23264 4231 -23248 4265
rect -23314 4197 -23248 4231
rect -23314 4163 -23298 4197
rect -23264 4163 -23248 4197
rect -23314 4129 -23248 4163
rect -23314 4095 -23298 4129
rect -23264 4095 -23248 4129
rect -23314 4061 -23248 4095
rect -23314 4027 -23298 4061
rect -23264 4027 -23248 4061
rect -23314 3993 -23248 4027
rect -23314 3959 -23298 3993
rect -23264 3959 -23248 3993
rect -23314 3925 -23248 3959
rect -23314 3891 -23298 3925
rect -23264 3891 -23248 3925
rect -23314 3857 -23248 3891
rect -23314 3823 -23298 3857
rect -23264 3823 -23248 3857
rect -23314 3789 -23248 3823
rect -23314 3755 -23298 3789
rect -23264 3755 -23248 3789
rect -23314 3721 -23248 3755
rect -23314 3687 -23298 3721
rect -23264 3687 -23248 3721
rect -23314 3653 -23248 3687
rect -23314 3619 -23298 3653
rect -23264 3619 -23248 3653
rect -23314 3585 -23248 3619
rect -23314 3551 -23298 3585
rect -23264 3551 -23248 3585
rect -23314 3517 -23248 3551
rect -23314 3483 -23298 3517
rect -23264 3483 -23248 3517
rect -23314 3442 -23248 3483
rect -23218 4401 -23152 4442
rect -23218 4367 -23202 4401
rect -23168 4367 -23152 4401
rect -23218 4333 -23152 4367
rect -23218 4299 -23202 4333
rect -23168 4299 -23152 4333
rect -23218 4265 -23152 4299
rect -23218 4231 -23202 4265
rect -23168 4231 -23152 4265
rect -23218 4197 -23152 4231
rect -23218 4163 -23202 4197
rect -23168 4163 -23152 4197
rect -23218 4129 -23152 4163
rect -23218 4095 -23202 4129
rect -23168 4095 -23152 4129
rect -23218 4061 -23152 4095
rect -23218 4027 -23202 4061
rect -23168 4027 -23152 4061
rect -23218 3993 -23152 4027
rect -23218 3959 -23202 3993
rect -23168 3959 -23152 3993
rect -23218 3925 -23152 3959
rect -23218 3891 -23202 3925
rect -23168 3891 -23152 3925
rect -23218 3857 -23152 3891
rect -23218 3823 -23202 3857
rect -23168 3823 -23152 3857
rect -23218 3789 -23152 3823
rect -23218 3755 -23202 3789
rect -23168 3755 -23152 3789
rect -23218 3721 -23152 3755
rect -23218 3687 -23202 3721
rect -23168 3687 -23152 3721
rect -23218 3653 -23152 3687
rect -23218 3619 -23202 3653
rect -23168 3619 -23152 3653
rect -23218 3585 -23152 3619
rect -23218 3551 -23202 3585
rect -23168 3551 -23152 3585
rect -23218 3517 -23152 3551
rect -23218 3483 -23202 3517
rect -23168 3483 -23152 3517
rect -23218 3442 -23152 3483
rect -23122 4401 -23056 4442
rect -23122 4367 -23106 4401
rect -23072 4367 -23056 4401
rect -23122 4333 -23056 4367
rect -23122 4299 -23106 4333
rect -23072 4299 -23056 4333
rect -23122 4265 -23056 4299
rect -23122 4231 -23106 4265
rect -23072 4231 -23056 4265
rect -23122 4197 -23056 4231
rect -23122 4163 -23106 4197
rect -23072 4163 -23056 4197
rect -23122 4129 -23056 4163
rect -23122 4095 -23106 4129
rect -23072 4095 -23056 4129
rect -23122 4061 -23056 4095
rect -23122 4027 -23106 4061
rect -23072 4027 -23056 4061
rect -23122 3993 -23056 4027
rect -23122 3959 -23106 3993
rect -23072 3959 -23056 3993
rect -23122 3925 -23056 3959
rect -23122 3891 -23106 3925
rect -23072 3891 -23056 3925
rect -23122 3857 -23056 3891
rect -23122 3823 -23106 3857
rect -23072 3823 -23056 3857
rect -23122 3789 -23056 3823
rect -23122 3755 -23106 3789
rect -23072 3755 -23056 3789
rect -23122 3721 -23056 3755
rect -23122 3687 -23106 3721
rect -23072 3687 -23056 3721
rect -23122 3653 -23056 3687
rect -23122 3619 -23106 3653
rect -23072 3619 -23056 3653
rect -23122 3585 -23056 3619
rect -23122 3551 -23106 3585
rect -23072 3551 -23056 3585
rect -23122 3517 -23056 3551
rect -23122 3483 -23106 3517
rect -23072 3483 -23056 3517
rect -23122 3442 -23056 3483
rect -23026 4401 -22960 4442
rect -23026 4367 -23010 4401
rect -22976 4367 -22960 4401
rect -23026 4333 -22960 4367
rect -23026 4299 -23010 4333
rect -22976 4299 -22960 4333
rect -23026 4265 -22960 4299
rect -23026 4231 -23010 4265
rect -22976 4231 -22960 4265
rect -23026 4197 -22960 4231
rect -23026 4163 -23010 4197
rect -22976 4163 -22960 4197
rect -23026 4129 -22960 4163
rect -23026 4095 -23010 4129
rect -22976 4095 -22960 4129
rect -23026 4061 -22960 4095
rect -23026 4027 -23010 4061
rect -22976 4027 -22960 4061
rect -23026 3993 -22960 4027
rect -23026 3959 -23010 3993
rect -22976 3959 -22960 3993
rect -23026 3925 -22960 3959
rect -23026 3891 -23010 3925
rect -22976 3891 -22960 3925
rect -23026 3857 -22960 3891
rect -23026 3823 -23010 3857
rect -22976 3823 -22960 3857
rect -23026 3789 -22960 3823
rect -23026 3755 -23010 3789
rect -22976 3755 -22960 3789
rect -23026 3721 -22960 3755
rect -23026 3687 -23010 3721
rect -22976 3687 -22960 3721
rect -23026 3653 -22960 3687
rect -23026 3619 -23010 3653
rect -22976 3619 -22960 3653
rect -23026 3585 -22960 3619
rect -23026 3551 -23010 3585
rect -22976 3551 -22960 3585
rect -23026 3517 -22960 3551
rect -23026 3483 -23010 3517
rect -22976 3483 -22960 3517
rect -23026 3442 -22960 3483
rect -22930 4401 -22864 4442
rect -22930 4367 -22914 4401
rect -22880 4367 -22864 4401
rect -22930 4333 -22864 4367
rect -22930 4299 -22914 4333
rect -22880 4299 -22864 4333
rect -22930 4265 -22864 4299
rect -22930 4231 -22914 4265
rect -22880 4231 -22864 4265
rect -22930 4197 -22864 4231
rect -22930 4163 -22914 4197
rect -22880 4163 -22864 4197
rect -22930 4129 -22864 4163
rect -22930 4095 -22914 4129
rect -22880 4095 -22864 4129
rect -22930 4061 -22864 4095
rect -22930 4027 -22914 4061
rect -22880 4027 -22864 4061
rect -22930 3993 -22864 4027
rect -22930 3959 -22914 3993
rect -22880 3959 -22864 3993
rect -22930 3925 -22864 3959
rect -22930 3891 -22914 3925
rect -22880 3891 -22864 3925
rect -22930 3857 -22864 3891
rect -22930 3823 -22914 3857
rect -22880 3823 -22864 3857
rect -22930 3789 -22864 3823
rect -22930 3755 -22914 3789
rect -22880 3755 -22864 3789
rect -22930 3721 -22864 3755
rect -22930 3687 -22914 3721
rect -22880 3687 -22864 3721
rect -22930 3653 -22864 3687
rect -22930 3619 -22914 3653
rect -22880 3619 -22864 3653
rect -22930 3585 -22864 3619
rect -22930 3551 -22914 3585
rect -22880 3551 -22864 3585
rect -22930 3517 -22864 3551
rect -22930 3483 -22914 3517
rect -22880 3483 -22864 3517
rect -22930 3442 -22864 3483
rect -22834 4401 -22768 4442
rect -22834 4367 -22818 4401
rect -22784 4367 -22768 4401
rect -22834 4333 -22768 4367
rect -22834 4299 -22818 4333
rect -22784 4299 -22768 4333
rect -22834 4265 -22768 4299
rect -22834 4231 -22818 4265
rect -22784 4231 -22768 4265
rect -22834 4197 -22768 4231
rect -22834 4163 -22818 4197
rect -22784 4163 -22768 4197
rect -22834 4129 -22768 4163
rect -22834 4095 -22818 4129
rect -22784 4095 -22768 4129
rect -22834 4061 -22768 4095
rect -22834 4027 -22818 4061
rect -22784 4027 -22768 4061
rect -22834 3993 -22768 4027
rect -22834 3959 -22818 3993
rect -22784 3959 -22768 3993
rect -22834 3925 -22768 3959
rect -22834 3891 -22818 3925
rect -22784 3891 -22768 3925
rect -22834 3857 -22768 3891
rect -22834 3823 -22818 3857
rect -22784 3823 -22768 3857
rect -22834 3789 -22768 3823
rect -22834 3755 -22818 3789
rect -22784 3755 -22768 3789
rect -22834 3721 -22768 3755
rect -22834 3687 -22818 3721
rect -22784 3687 -22768 3721
rect -22834 3653 -22768 3687
rect -22834 3619 -22818 3653
rect -22784 3619 -22768 3653
rect -22834 3585 -22768 3619
rect -22834 3551 -22818 3585
rect -22784 3551 -22768 3585
rect -22834 3517 -22768 3551
rect -22834 3483 -22818 3517
rect -22784 3483 -22768 3517
rect -22834 3442 -22768 3483
rect -22738 4401 -22672 4442
rect -22738 4367 -22722 4401
rect -22688 4367 -22672 4401
rect -22738 4333 -22672 4367
rect -22738 4299 -22722 4333
rect -22688 4299 -22672 4333
rect -22738 4265 -22672 4299
rect -22738 4231 -22722 4265
rect -22688 4231 -22672 4265
rect -22738 4197 -22672 4231
rect -22738 4163 -22722 4197
rect -22688 4163 -22672 4197
rect -22738 4129 -22672 4163
rect -22738 4095 -22722 4129
rect -22688 4095 -22672 4129
rect -22738 4061 -22672 4095
rect -22738 4027 -22722 4061
rect -22688 4027 -22672 4061
rect -22738 3993 -22672 4027
rect -22738 3959 -22722 3993
rect -22688 3959 -22672 3993
rect -22738 3925 -22672 3959
rect -22738 3891 -22722 3925
rect -22688 3891 -22672 3925
rect -22738 3857 -22672 3891
rect -22738 3823 -22722 3857
rect -22688 3823 -22672 3857
rect -22738 3789 -22672 3823
rect -22738 3755 -22722 3789
rect -22688 3755 -22672 3789
rect -22738 3721 -22672 3755
rect -22738 3687 -22722 3721
rect -22688 3687 -22672 3721
rect -22738 3653 -22672 3687
rect -22738 3619 -22722 3653
rect -22688 3619 -22672 3653
rect -22738 3585 -22672 3619
rect -22738 3551 -22722 3585
rect -22688 3551 -22672 3585
rect -22738 3517 -22672 3551
rect -22738 3483 -22722 3517
rect -22688 3483 -22672 3517
rect -22738 3442 -22672 3483
rect -22642 4401 -22576 4442
rect -22642 4367 -22626 4401
rect -22592 4367 -22576 4401
rect -22642 4333 -22576 4367
rect -22642 4299 -22626 4333
rect -22592 4299 -22576 4333
rect -22642 4265 -22576 4299
rect -22642 4231 -22626 4265
rect -22592 4231 -22576 4265
rect -22642 4197 -22576 4231
rect -22642 4163 -22626 4197
rect -22592 4163 -22576 4197
rect -22642 4129 -22576 4163
rect -22642 4095 -22626 4129
rect -22592 4095 -22576 4129
rect -22642 4061 -22576 4095
rect -22642 4027 -22626 4061
rect -22592 4027 -22576 4061
rect -22642 3993 -22576 4027
rect -22642 3959 -22626 3993
rect -22592 3959 -22576 3993
rect -22642 3925 -22576 3959
rect -22642 3891 -22626 3925
rect -22592 3891 -22576 3925
rect -22642 3857 -22576 3891
rect -22642 3823 -22626 3857
rect -22592 3823 -22576 3857
rect -22642 3789 -22576 3823
rect -22642 3755 -22626 3789
rect -22592 3755 -22576 3789
rect -22642 3721 -22576 3755
rect -22642 3687 -22626 3721
rect -22592 3687 -22576 3721
rect -22642 3653 -22576 3687
rect -22642 3619 -22626 3653
rect -22592 3619 -22576 3653
rect -22642 3585 -22576 3619
rect -22642 3551 -22626 3585
rect -22592 3551 -22576 3585
rect -22642 3517 -22576 3551
rect -22642 3483 -22626 3517
rect -22592 3483 -22576 3517
rect -22642 3442 -22576 3483
rect -22546 4401 -22480 4442
rect -22546 4367 -22530 4401
rect -22496 4367 -22480 4401
rect -22546 4333 -22480 4367
rect -22546 4299 -22530 4333
rect -22496 4299 -22480 4333
rect -22546 4265 -22480 4299
rect -22546 4231 -22530 4265
rect -22496 4231 -22480 4265
rect -22546 4197 -22480 4231
rect -22546 4163 -22530 4197
rect -22496 4163 -22480 4197
rect -22546 4129 -22480 4163
rect -22546 4095 -22530 4129
rect -22496 4095 -22480 4129
rect -22546 4061 -22480 4095
rect -22546 4027 -22530 4061
rect -22496 4027 -22480 4061
rect -22546 3993 -22480 4027
rect -22546 3959 -22530 3993
rect -22496 3959 -22480 3993
rect -22546 3925 -22480 3959
rect -22546 3891 -22530 3925
rect -22496 3891 -22480 3925
rect -22546 3857 -22480 3891
rect -22546 3823 -22530 3857
rect -22496 3823 -22480 3857
rect -22546 3789 -22480 3823
rect -22546 3755 -22530 3789
rect -22496 3755 -22480 3789
rect -22546 3721 -22480 3755
rect -22546 3687 -22530 3721
rect -22496 3687 -22480 3721
rect -22546 3653 -22480 3687
rect -22546 3619 -22530 3653
rect -22496 3619 -22480 3653
rect -22546 3585 -22480 3619
rect -22546 3551 -22530 3585
rect -22496 3551 -22480 3585
rect -22546 3517 -22480 3551
rect -22546 3483 -22530 3517
rect -22496 3483 -22480 3517
rect -22546 3442 -22480 3483
rect -22450 4401 -22384 4442
rect -22450 4367 -22434 4401
rect -22400 4367 -22384 4401
rect -22450 4333 -22384 4367
rect -22450 4299 -22434 4333
rect -22400 4299 -22384 4333
rect -22450 4265 -22384 4299
rect -22450 4231 -22434 4265
rect -22400 4231 -22384 4265
rect -22450 4197 -22384 4231
rect -22450 4163 -22434 4197
rect -22400 4163 -22384 4197
rect -22450 4129 -22384 4163
rect -22450 4095 -22434 4129
rect -22400 4095 -22384 4129
rect -22450 4061 -22384 4095
rect -22450 4027 -22434 4061
rect -22400 4027 -22384 4061
rect -22450 3993 -22384 4027
rect -22450 3959 -22434 3993
rect -22400 3959 -22384 3993
rect -22450 3925 -22384 3959
rect -22450 3891 -22434 3925
rect -22400 3891 -22384 3925
rect -22450 3857 -22384 3891
rect -22450 3823 -22434 3857
rect -22400 3823 -22384 3857
rect -22450 3789 -22384 3823
rect -22450 3755 -22434 3789
rect -22400 3755 -22384 3789
rect -22450 3721 -22384 3755
rect -22450 3687 -22434 3721
rect -22400 3687 -22384 3721
rect -22450 3653 -22384 3687
rect -22450 3619 -22434 3653
rect -22400 3619 -22384 3653
rect -22450 3585 -22384 3619
rect -22450 3551 -22434 3585
rect -22400 3551 -22384 3585
rect -22450 3517 -22384 3551
rect -22450 3483 -22434 3517
rect -22400 3483 -22384 3517
rect -22450 3442 -22384 3483
rect -22354 4401 -22288 4442
rect -22354 4367 -22338 4401
rect -22304 4367 -22288 4401
rect -22354 4333 -22288 4367
rect -22354 4299 -22338 4333
rect -22304 4299 -22288 4333
rect -22354 4265 -22288 4299
rect -22354 4231 -22338 4265
rect -22304 4231 -22288 4265
rect -22354 4197 -22288 4231
rect -22354 4163 -22338 4197
rect -22304 4163 -22288 4197
rect -22354 4129 -22288 4163
rect -22354 4095 -22338 4129
rect -22304 4095 -22288 4129
rect -22354 4061 -22288 4095
rect -22354 4027 -22338 4061
rect -22304 4027 -22288 4061
rect -22354 3993 -22288 4027
rect -22354 3959 -22338 3993
rect -22304 3959 -22288 3993
rect -22354 3925 -22288 3959
rect -22354 3891 -22338 3925
rect -22304 3891 -22288 3925
rect -22354 3857 -22288 3891
rect -22354 3823 -22338 3857
rect -22304 3823 -22288 3857
rect -22354 3789 -22288 3823
rect -22354 3755 -22338 3789
rect -22304 3755 -22288 3789
rect -22354 3721 -22288 3755
rect -22354 3687 -22338 3721
rect -22304 3687 -22288 3721
rect -22354 3653 -22288 3687
rect -22354 3619 -22338 3653
rect -22304 3619 -22288 3653
rect -22354 3585 -22288 3619
rect -22354 3551 -22338 3585
rect -22304 3551 -22288 3585
rect -22354 3517 -22288 3551
rect -22354 3483 -22338 3517
rect -22304 3483 -22288 3517
rect -22354 3442 -22288 3483
rect -22258 4401 -22192 4442
rect -22258 4367 -22242 4401
rect -22208 4367 -22192 4401
rect -22258 4333 -22192 4367
rect -22258 4299 -22242 4333
rect -22208 4299 -22192 4333
rect -22258 4265 -22192 4299
rect -22258 4231 -22242 4265
rect -22208 4231 -22192 4265
rect -22258 4197 -22192 4231
rect -22258 4163 -22242 4197
rect -22208 4163 -22192 4197
rect -22258 4129 -22192 4163
rect -22258 4095 -22242 4129
rect -22208 4095 -22192 4129
rect -22258 4061 -22192 4095
rect -22258 4027 -22242 4061
rect -22208 4027 -22192 4061
rect -22258 3993 -22192 4027
rect -22258 3959 -22242 3993
rect -22208 3959 -22192 3993
rect -22258 3925 -22192 3959
rect -22258 3891 -22242 3925
rect -22208 3891 -22192 3925
rect -22258 3857 -22192 3891
rect -22258 3823 -22242 3857
rect -22208 3823 -22192 3857
rect -22258 3789 -22192 3823
rect -22258 3755 -22242 3789
rect -22208 3755 -22192 3789
rect -22258 3721 -22192 3755
rect -22258 3687 -22242 3721
rect -22208 3687 -22192 3721
rect -22258 3653 -22192 3687
rect -22258 3619 -22242 3653
rect -22208 3619 -22192 3653
rect -22258 3585 -22192 3619
rect -22258 3551 -22242 3585
rect -22208 3551 -22192 3585
rect -22258 3517 -22192 3551
rect -22258 3483 -22242 3517
rect -22208 3483 -22192 3517
rect -22258 3442 -22192 3483
rect -22162 4401 -22096 4442
rect -22162 4367 -22146 4401
rect -22112 4367 -22096 4401
rect -22162 4333 -22096 4367
rect -22162 4299 -22146 4333
rect -22112 4299 -22096 4333
rect -22162 4265 -22096 4299
rect -22162 4231 -22146 4265
rect -22112 4231 -22096 4265
rect -22162 4197 -22096 4231
rect -22162 4163 -22146 4197
rect -22112 4163 -22096 4197
rect -22162 4129 -22096 4163
rect -22162 4095 -22146 4129
rect -22112 4095 -22096 4129
rect -22162 4061 -22096 4095
rect -22162 4027 -22146 4061
rect -22112 4027 -22096 4061
rect -22162 3993 -22096 4027
rect -22162 3959 -22146 3993
rect -22112 3959 -22096 3993
rect -22162 3925 -22096 3959
rect -22162 3891 -22146 3925
rect -22112 3891 -22096 3925
rect -22162 3857 -22096 3891
rect -22162 3823 -22146 3857
rect -22112 3823 -22096 3857
rect -22162 3789 -22096 3823
rect -22162 3755 -22146 3789
rect -22112 3755 -22096 3789
rect -22162 3721 -22096 3755
rect -22162 3687 -22146 3721
rect -22112 3687 -22096 3721
rect -22162 3653 -22096 3687
rect -22162 3619 -22146 3653
rect -22112 3619 -22096 3653
rect -22162 3585 -22096 3619
rect -22162 3551 -22146 3585
rect -22112 3551 -22096 3585
rect -22162 3517 -22096 3551
rect -22162 3483 -22146 3517
rect -22112 3483 -22096 3517
rect -22162 3442 -22096 3483
rect -22066 4401 -22000 4442
rect -22066 4367 -22050 4401
rect -22016 4367 -22000 4401
rect -22066 4333 -22000 4367
rect -22066 4299 -22050 4333
rect -22016 4299 -22000 4333
rect -22066 4265 -22000 4299
rect -22066 4231 -22050 4265
rect -22016 4231 -22000 4265
rect -22066 4197 -22000 4231
rect -22066 4163 -22050 4197
rect -22016 4163 -22000 4197
rect -22066 4129 -22000 4163
rect -22066 4095 -22050 4129
rect -22016 4095 -22000 4129
rect -22066 4061 -22000 4095
rect -22066 4027 -22050 4061
rect -22016 4027 -22000 4061
rect -22066 3993 -22000 4027
rect -22066 3959 -22050 3993
rect -22016 3959 -22000 3993
rect -22066 3925 -22000 3959
rect -22066 3891 -22050 3925
rect -22016 3891 -22000 3925
rect -22066 3857 -22000 3891
rect -22066 3823 -22050 3857
rect -22016 3823 -22000 3857
rect -22066 3789 -22000 3823
rect -22066 3755 -22050 3789
rect -22016 3755 -22000 3789
rect -22066 3721 -22000 3755
rect -22066 3687 -22050 3721
rect -22016 3687 -22000 3721
rect -22066 3653 -22000 3687
rect -22066 3619 -22050 3653
rect -22016 3619 -22000 3653
rect -22066 3585 -22000 3619
rect -22066 3551 -22050 3585
rect -22016 3551 -22000 3585
rect -22066 3517 -22000 3551
rect -22066 3483 -22050 3517
rect -22016 3483 -22000 3517
rect -22066 3442 -22000 3483
rect -21970 4401 -21904 4442
rect -21970 4367 -21954 4401
rect -21920 4367 -21904 4401
rect -21970 4333 -21904 4367
rect -21970 4299 -21954 4333
rect -21920 4299 -21904 4333
rect -21970 4265 -21904 4299
rect -21970 4231 -21954 4265
rect -21920 4231 -21904 4265
rect -21970 4197 -21904 4231
rect -21970 4163 -21954 4197
rect -21920 4163 -21904 4197
rect -21970 4129 -21904 4163
rect -21970 4095 -21954 4129
rect -21920 4095 -21904 4129
rect -21970 4061 -21904 4095
rect -21970 4027 -21954 4061
rect -21920 4027 -21904 4061
rect -21970 3993 -21904 4027
rect -21970 3959 -21954 3993
rect -21920 3959 -21904 3993
rect -21970 3925 -21904 3959
rect -21970 3891 -21954 3925
rect -21920 3891 -21904 3925
rect -21970 3857 -21904 3891
rect -21970 3823 -21954 3857
rect -21920 3823 -21904 3857
rect -21970 3789 -21904 3823
rect -21970 3755 -21954 3789
rect -21920 3755 -21904 3789
rect -21970 3721 -21904 3755
rect -21970 3687 -21954 3721
rect -21920 3687 -21904 3721
rect -21970 3653 -21904 3687
rect -21970 3619 -21954 3653
rect -21920 3619 -21904 3653
rect -21970 3585 -21904 3619
rect -21970 3551 -21954 3585
rect -21920 3551 -21904 3585
rect -21970 3517 -21904 3551
rect -21970 3483 -21954 3517
rect -21920 3483 -21904 3517
rect -21970 3442 -21904 3483
rect -21874 4401 -21808 4442
rect -21874 4367 -21858 4401
rect -21824 4367 -21808 4401
rect -21874 4333 -21808 4367
rect -21874 4299 -21858 4333
rect -21824 4299 -21808 4333
rect -21874 4265 -21808 4299
rect -21874 4231 -21858 4265
rect -21824 4231 -21808 4265
rect -21874 4197 -21808 4231
rect -21874 4163 -21858 4197
rect -21824 4163 -21808 4197
rect -21874 4129 -21808 4163
rect -21874 4095 -21858 4129
rect -21824 4095 -21808 4129
rect -21874 4061 -21808 4095
rect -21874 4027 -21858 4061
rect -21824 4027 -21808 4061
rect -21874 3993 -21808 4027
rect -21874 3959 -21858 3993
rect -21824 3959 -21808 3993
rect -21874 3925 -21808 3959
rect -21874 3891 -21858 3925
rect -21824 3891 -21808 3925
rect -21874 3857 -21808 3891
rect -21874 3823 -21858 3857
rect -21824 3823 -21808 3857
rect -21874 3789 -21808 3823
rect -21874 3755 -21858 3789
rect -21824 3755 -21808 3789
rect -21874 3721 -21808 3755
rect -21874 3687 -21858 3721
rect -21824 3687 -21808 3721
rect -21874 3653 -21808 3687
rect -21874 3619 -21858 3653
rect -21824 3619 -21808 3653
rect -21874 3585 -21808 3619
rect -21874 3551 -21858 3585
rect -21824 3551 -21808 3585
rect -21874 3517 -21808 3551
rect -21874 3483 -21858 3517
rect -21824 3483 -21808 3517
rect -21874 3442 -21808 3483
rect -21778 4401 -21712 4442
rect -21778 4367 -21762 4401
rect -21728 4367 -21712 4401
rect -21778 4333 -21712 4367
rect -21778 4299 -21762 4333
rect -21728 4299 -21712 4333
rect -21778 4265 -21712 4299
rect -21778 4231 -21762 4265
rect -21728 4231 -21712 4265
rect -21778 4197 -21712 4231
rect -21778 4163 -21762 4197
rect -21728 4163 -21712 4197
rect -21778 4129 -21712 4163
rect -21778 4095 -21762 4129
rect -21728 4095 -21712 4129
rect -21778 4061 -21712 4095
rect -21778 4027 -21762 4061
rect -21728 4027 -21712 4061
rect -21778 3993 -21712 4027
rect -21778 3959 -21762 3993
rect -21728 3959 -21712 3993
rect -21778 3925 -21712 3959
rect -21778 3891 -21762 3925
rect -21728 3891 -21712 3925
rect -21778 3857 -21712 3891
rect -21778 3823 -21762 3857
rect -21728 3823 -21712 3857
rect -21778 3789 -21712 3823
rect -21778 3755 -21762 3789
rect -21728 3755 -21712 3789
rect -21778 3721 -21712 3755
rect -21778 3687 -21762 3721
rect -21728 3687 -21712 3721
rect -21778 3653 -21712 3687
rect -21778 3619 -21762 3653
rect -21728 3619 -21712 3653
rect -21778 3585 -21712 3619
rect -21778 3551 -21762 3585
rect -21728 3551 -21712 3585
rect -21778 3517 -21712 3551
rect -21778 3483 -21762 3517
rect -21728 3483 -21712 3517
rect -21778 3442 -21712 3483
rect -21682 4401 -21620 4442
rect -21682 4367 -21666 4401
rect -21632 4367 -21620 4401
rect -21682 4333 -21620 4367
rect -21682 4299 -21666 4333
rect -21632 4299 -21620 4333
rect -21682 4265 -21620 4299
rect -21682 4231 -21666 4265
rect -21632 4231 -21620 4265
rect -21682 4197 -21620 4231
rect -21682 4163 -21666 4197
rect -21632 4163 -21620 4197
rect -21682 4129 -21620 4163
rect -21682 4095 -21666 4129
rect -21632 4095 -21620 4129
rect -21682 4061 -21620 4095
rect -21682 4027 -21666 4061
rect -21632 4027 -21620 4061
rect -21682 3993 -21620 4027
rect -21682 3959 -21666 3993
rect -21632 3959 -21620 3993
rect -21682 3925 -21620 3959
rect -21682 3891 -21666 3925
rect -21632 3891 -21620 3925
rect -21682 3857 -21620 3891
rect -21682 3823 -21666 3857
rect -21632 3823 -21620 3857
rect -21682 3789 -21620 3823
rect -21682 3755 -21666 3789
rect -21632 3755 -21620 3789
rect -21682 3721 -21620 3755
rect -21682 3687 -21666 3721
rect -21632 3687 -21620 3721
rect -21682 3653 -21620 3687
rect -21682 3619 -21666 3653
rect -21632 3619 -21620 3653
rect -21682 3585 -21620 3619
rect -21682 3551 -21666 3585
rect -21632 3551 -21620 3585
rect -21682 3517 -21620 3551
rect -21682 3483 -21666 3517
rect -21632 3483 -21620 3517
rect -21682 3442 -21620 3483
rect -21454 4407 -21392 4448
rect -21454 4373 -21442 4407
rect -21408 4373 -21392 4407
rect -21454 4339 -21392 4373
rect -21454 4305 -21442 4339
rect -21408 4305 -21392 4339
rect -21454 4271 -21392 4305
rect -21454 4237 -21442 4271
rect -21408 4237 -21392 4271
rect -21454 4203 -21392 4237
rect -21454 4169 -21442 4203
rect -21408 4169 -21392 4203
rect -21454 4135 -21392 4169
rect -21454 4101 -21442 4135
rect -21408 4101 -21392 4135
rect -21454 4067 -21392 4101
rect -21454 4033 -21442 4067
rect -21408 4033 -21392 4067
rect -21454 3999 -21392 4033
rect -21454 3965 -21442 3999
rect -21408 3965 -21392 3999
rect -21454 3931 -21392 3965
rect -21454 3897 -21442 3931
rect -21408 3897 -21392 3931
rect -21454 3863 -21392 3897
rect -21454 3829 -21442 3863
rect -21408 3829 -21392 3863
rect -21454 3795 -21392 3829
rect -21454 3761 -21442 3795
rect -21408 3761 -21392 3795
rect -21454 3727 -21392 3761
rect -21454 3693 -21442 3727
rect -21408 3693 -21392 3727
rect -21454 3659 -21392 3693
rect -21454 3625 -21442 3659
rect -21408 3625 -21392 3659
rect -21454 3591 -21392 3625
rect -21454 3557 -21442 3591
rect -21408 3557 -21392 3591
rect -21454 3523 -21392 3557
rect -21454 3489 -21442 3523
rect -21408 3489 -21392 3523
rect -21454 3448 -21392 3489
rect -21362 4407 -21296 4448
rect -21362 4373 -21346 4407
rect -21312 4373 -21296 4407
rect -21362 4339 -21296 4373
rect -21362 4305 -21346 4339
rect -21312 4305 -21296 4339
rect -21362 4271 -21296 4305
rect -21362 4237 -21346 4271
rect -21312 4237 -21296 4271
rect -21362 4203 -21296 4237
rect -21362 4169 -21346 4203
rect -21312 4169 -21296 4203
rect -21362 4135 -21296 4169
rect -21362 4101 -21346 4135
rect -21312 4101 -21296 4135
rect -21362 4067 -21296 4101
rect -21362 4033 -21346 4067
rect -21312 4033 -21296 4067
rect -21362 3999 -21296 4033
rect -21362 3965 -21346 3999
rect -21312 3965 -21296 3999
rect -21362 3931 -21296 3965
rect -21362 3897 -21346 3931
rect -21312 3897 -21296 3931
rect -21362 3863 -21296 3897
rect -21362 3829 -21346 3863
rect -21312 3829 -21296 3863
rect -21362 3795 -21296 3829
rect -21362 3761 -21346 3795
rect -21312 3761 -21296 3795
rect -21362 3727 -21296 3761
rect -21362 3693 -21346 3727
rect -21312 3693 -21296 3727
rect -21362 3659 -21296 3693
rect -21362 3625 -21346 3659
rect -21312 3625 -21296 3659
rect -21362 3591 -21296 3625
rect -21362 3557 -21346 3591
rect -21312 3557 -21296 3591
rect -21362 3523 -21296 3557
rect -21362 3489 -21346 3523
rect -21312 3489 -21296 3523
rect -21362 3448 -21296 3489
rect -21266 4407 -21200 4448
rect -21266 4373 -21250 4407
rect -21216 4373 -21200 4407
rect -21266 4339 -21200 4373
rect -21266 4305 -21250 4339
rect -21216 4305 -21200 4339
rect -21266 4271 -21200 4305
rect -21266 4237 -21250 4271
rect -21216 4237 -21200 4271
rect -21266 4203 -21200 4237
rect -21266 4169 -21250 4203
rect -21216 4169 -21200 4203
rect -21266 4135 -21200 4169
rect -21266 4101 -21250 4135
rect -21216 4101 -21200 4135
rect -21266 4067 -21200 4101
rect -21266 4033 -21250 4067
rect -21216 4033 -21200 4067
rect -21266 3999 -21200 4033
rect -21266 3965 -21250 3999
rect -21216 3965 -21200 3999
rect -21266 3931 -21200 3965
rect -21266 3897 -21250 3931
rect -21216 3897 -21200 3931
rect -21266 3863 -21200 3897
rect -21266 3829 -21250 3863
rect -21216 3829 -21200 3863
rect -21266 3795 -21200 3829
rect -21266 3761 -21250 3795
rect -21216 3761 -21200 3795
rect -21266 3727 -21200 3761
rect -21266 3693 -21250 3727
rect -21216 3693 -21200 3727
rect -21266 3659 -21200 3693
rect -21266 3625 -21250 3659
rect -21216 3625 -21200 3659
rect -21266 3591 -21200 3625
rect -21266 3557 -21250 3591
rect -21216 3557 -21200 3591
rect -21266 3523 -21200 3557
rect -21266 3489 -21250 3523
rect -21216 3489 -21200 3523
rect -21266 3448 -21200 3489
rect -21170 4407 -21104 4448
rect -21170 4373 -21154 4407
rect -21120 4373 -21104 4407
rect -21170 4339 -21104 4373
rect -21170 4305 -21154 4339
rect -21120 4305 -21104 4339
rect -21170 4271 -21104 4305
rect -21170 4237 -21154 4271
rect -21120 4237 -21104 4271
rect -21170 4203 -21104 4237
rect -21170 4169 -21154 4203
rect -21120 4169 -21104 4203
rect -21170 4135 -21104 4169
rect -21170 4101 -21154 4135
rect -21120 4101 -21104 4135
rect -21170 4067 -21104 4101
rect -21170 4033 -21154 4067
rect -21120 4033 -21104 4067
rect -21170 3999 -21104 4033
rect -21170 3965 -21154 3999
rect -21120 3965 -21104 3999
rect -21170 3931 -21104 3965
rect -21170 3897 -21154 3931
rect -21120 3897 -21104 3931
rect -21170 3863 -21104 3897
rect -21170 3829 -21154 3863
rect -21120 3829 -21104 3863
rect -21170 3795 -21104 3829
rect -21170 3761 -21154 3795
rect -21120 3761 -21104 3795
rect -21170 3727 -21104 3761
rect -21170 3693 -21154 3727
rect -21120 3693 -21104 3727
rect -21170 3659 -21104 3693
rect -21170 3625 -21154 3659
rect -21120 3625 -21104 3659
rect -21170 3591 -21104 3625
rect -21170 3557 -21154 3591
rect -21120 3557 -21104 3591
rect -21170 3523 -21104 3557
rect -21170 3489 -21154 3523
rect -21120 3489 -21104 3523
rect -21170 3448 -21104 3489
rect -21074 4407 -21008 4448
rect -21074 4373 -21058 4407
rect -21024 4373 -21008 4407
rect -21074 4339 -21008 4373
rect -21074 4305 -21058 4339
rect -21024 4305 -21008 4339
rect -21074 4271 -21008 4305
rect -21074 4237 -21058 4271
rect -21024 4237 -21008 4271
rect -21074 4203 -21008 4237
rect -21074 4169 -21058 4203
rect -21024 4169 -21008 4203
rect -21074 4135 -21008 4169
rect -21074 4101 -21058 4135
rect -21024 4101 -21008 4135
rect -21074 4067 -21008 4101
rect -21074 4033 -21058 4067
rect -21024 4033 -21008 4067
rect -21074 3999 -21008 4033
rect -21074 3965 -21058 3999
rect -21024 3965 -21008 3999
rect -21074 3931 -21008 3965
rect -21074 3897 -21058 3931
rect -21024 3897 -21008 3931
rect -21074 3863 -21008 3897
rect -21074 3829 -21058 3863
rect -21024 3829 -21008 3863
rect -21074 3795 -21008 3829
rect -21074 3761 -21058 3795
rect -21024 3761 -21008 3795
rect -21074 3727 -21008 3761
rect -21074 3693 -21058 3727
rect -21024 3693 -21008 3727
rect -21074 3659 -21008 3693
rect -21074 3625 -21058 3659
rect -21024 3625 -21008 3659
rect -21074 3591 -21008 3625
rect -21074 3557 -21058 3591
rect -21024 3557 -21008 3591
rect -21074 3523 -21008 3557
rect -21074 3489 -21058 3523
rect -21024 3489 -21008 3523
rect -21074 3448 -21008 3489
rect -20978 4407 -20912 4448
rect -20978 4373 -20962 4407
rect -20928 4373 -20912 4407
rect -20978 4339 -20912 4373
rect -20978 4305 -20962 4339
rect -20928 4305 -20912 4339
rect -20978 4271 -20912 4305
rect -20978 4237 -20962 4271
rect -20928 4237 -20912 4271
rect -20978 4203 -20912 4237
rect -20978 4169 -20962 4203
rect -20928 4169 -20912 4203
rect -20978 4135 -20912 4169
rect -20978 4101 -20962 4135
rect -20928 4101 -20912 4135
rect -20978 4067 -20912 4101
rect -20978 4033 -20962 4067
rect -20928 4033 -20912 4067
rect -20978 3999 -20912 4033
rect -20978 3965 -20962 3999
rect -20928 3965 -20912 3999
rect -20978 3931 -20912 3965
rect -20978 3897 -20962 3931
rect -20928 3897 -20912 3931
rect -20978 3863 -20912 3897
rect -20978 3829 -20962 3863
rect -20928 3829 -20912 3863
rect -20978 3795 -20912 3829
rect -20978 3761 -20962 3795
rect -20928 3761 -20912 3795
rect -20978 3727 -20912 3761
rect -20978 3693 -20962 3727
rect -20928 3693 -20912 3727
rect -20978 3659 -20912 3693
rect -20978 3625 -20962 3659
rect -20928 3625 -20912 3659
rect -20978 3591 -20912 3625
rect -20978 3557 -20962 3591
rect -20928 3557 -20912 3591
rect -20978 3523 -20912 3557
rect -20978 3489 -20962 3523
rect -20928 3489 -20912 3523
rect -20978 3448 -20912 3489
rect -20882 4407 -20816 4448
rect -20882 4373 -20866 4407
rect -20832 4373 -20816 4407
rect -20882 4339 -20816 4373
rect -20882 4305 -20866 4339
rect -20832 4305 -20816 4339
rect -20882 4271 -20816 4305
rect -20882 4237 -20866 4271
rect -20832 4237 -20816 4271
rect -20882 4203 -20816 4237
rect -20882 4169 -20866 4203
rect -20832 4169 -20816 4203
rect -20882 4135 -20816 4169
rect -20882 4101 -20866 4135
rect -20832 4101 -20816 4135
rect -20882 4067 -20816 4101
rect -20882 4033 -20866 4067
rect -20832 4033 -20816 4067
rect -20882 3999 -20816 4033
rect -20882 3965 -20866 3999
rect -20832 3965 -20816 3999
rect -20882 3931 -20816 3965
rect -20882 3897 -20866 3931
rect -20832 3897 -20816 3931
rect -20882 3863 -20816 3897
rect -20882 3829 -20866 3863
rect -20832 3829 -20816 3863
rect -20882 3795 -20816 3829
rect -20882 3761 -20866 3795
rect -20832 3761 -20816 3795
rect -20882 3727 -20816 3761
rect -20882 3693 -20866 3727
rect -20832 3693 -20816 3727
rect -20882 3659 -20816 3693
rect -20882 3625 -20866 3659
rect -20832 3625 -20816 3659
rect -20882 3591 -20816 3625
rect -20882 3557 -20866 3591
rect -20832 3557 -20816 3591
rect -20882 3523 -20816 3557
rect -20882 3489 -20866 3523
rect -20832 3489 -20816 3523
rect -20882 3448 -20816 3489
rect -20786 4407 -20720 4448
rect -20786 4373 -20770 4407
rect -20736 4373 -20720 4407
rect -20786 4339 -20720 4373
rect -20786 4305 -20770 4339
rect -20736 4305 -20720 4339
rect -20786 4271 -20720 4305
rect -20786 4237 -20770 4271
rect -20736 4237 -20720 4271
rect -20786 4203 -20720 4237
rect -20786 4169 -20770 4203
rect -20736 4169 -20720 4203
rect -20786 4135 -20720 4169
rect -20786 4101 -20770 4135
rect -20736 4101 -20720 4135
rect -20786 4067 -20720 4101
rect -20786 4033 -20770 4067
rect -20736 4033 -20720 4067
rect -20786 3999 -20720 4033
rect -20786 3965 -20770 3999
rect -20736 3965 -20720 3999
rect -20786 3931 -20720 3965
rect -20786 3897 -20770 3931
rect -20736 3897 -20720 3931
rect -20786 3863 -20720 3897
rect -20786 3829 -20770 3863
rect -20736 3829 -20720 3863
rect -20786 3795 -20720 3829
rect -20786 3761 -20770 3795
rect -20736 3761 -20720 3795
rect -20786 3727 -20720 3761
rect -20786 3693 -20770 3727
rect -20736 3693 -20720 3727
rect -20786 3659 -20720 3693
rect -20786 3625 -20770 3659
rect -20736 3625 -20720 3659
rect -20786 3591 -20720 3625
rect -20786 3557 -20770 3591
rect -20736 3557 -20720 3591
rect -20786 3523 -20720 3557
rect -20786 3489 -20770 3523
rect -20736 3489 -20720 3523
rect -20786 3448 -20720 3489
rect -20690 4407 -20624 4448
rect -20690 4373 -20674 4407
rect -20640 4373 -20624 4407
rect -20690 4339 -20624 4373
rect -20690 4305 -20674 4339
rect -20640 4305 -20624 4339
rect -20690 4271 -20624 4305
rect -20690 4237 -20674 4271
rect -20640 4237 -20624 4271
rect -20690 4203 -20624 4237
rect -20690 4169 -20674 4203
rect -20640 4169 -20624 4203
rect -20690 4135 -20624 4169
rect -20690 4101 -20674 4135
rect -20640 4101 -20624 4135
rect -20690 4067 -20624 4101
rect -20690 4033 -20674 4067
rect -20640 4033 -20624 4067
rect -20690 3999 -20624 4033
rect -20690 3965 -20674 3999
rect -20640 3965 -20624 3999
rect -20690 3931 -20624 3965
rect -20690 3897 -20674 3931
rect -20640 3897 -20624 3931
rect -20690 3863 -20624 3897
rect -20690 3829 -20674 3863
rect -20640 3829 -20624 3863
rect -20690 3795 -20624 3829
rect -20690 3761 -20674 3795
rect -20640 3761 -20624 3795
rect -20690 3727 -20624 3761
rect -20690 3693 -20674 3727
rect -20640 3693 -20624 3727
rect -20690 3659 -20624 3693
rect -20690 3625 -20674 3659
rect -20640 3625 -20624 3659
rect -20690 3591 -20624 3625
rect -20690 3557 -20674 3591
rect -20640 3557 -20624 3591
rect -20690 3523 -20624 3557
rect -20690 3489 -20674 3523
rect -20640 3489 -20624 3523
rect -20690 3448 -20624 3489
rect -20594 4407 -20528 4448
rect -20594 4373 -20578 4407
rect -20544 4373 -20528 4407
rect -20594 4339 -20528 4373
rect -20594 4305 -20578 4339
rect -20544 4305 -20528 4339
rect -20594 4271 -20528 4305
rect -20594 4237 -20578 4271
rect -20544 4237 -20528 4271
rect -20594 4203 -20528 4237
rect -20594 4169 -20578 4203
rect -20544 4169 -20528 4203
rect -20594 4135 -20528 4169
rect -20594 4101 -20578 4135
rect -20544 4101 -20528 4135
rect -20594 4067 -20528 4101
rect -20594 4033 -20578 4067
rect -20544 4033 -20528 4067
rect -20594 3999 -20528 4033
rect -20594 3965 -20578 3999
rect -20544 3965 -20528 3999
rect -20594 3931 -20528 3965
rect -20594 3897 -20578 3931
rect -20544 3897 -20528 3931
rect -20594 3863 -20528 3897
rect -20594 3829 -20578 3863
rect -20544 3829 -20528 3863
rect -20594 3795 -20528 3829
rect -20594 3761 -20578 3795
rect -20544 3761 -20528 3795
rect -20594 3727 -20528 3761
rect -20594 3693 -20578 3727
rect -20544 3693 -20528 3727
rect -20594 3659 -20528 3693
rect -20594 3625 -20578 3659
rect -20544 3625 -20528 3659
rect -20594 3591 -20528 3625
rect -20594 3557 -20578 3591
rect -20544 3557 -20528 3591
rect -20594 3523 -20528 3557
rect -20594 3489 -20578 3523
rect -20544 3489 -20528 3523
rect -20594 3448 -20528 3489
rect -20498 4407 -20432 4448
rect -20498 4373 -20482 4407
rect -20448 4373 -20432 4407
rect -20498 4339 -20432 4373
rect -20498 4305 -20482 4339
rect -20448 4305 -20432 4339
rect -20498 4271 -20432 4305
rect -20498 4237 -20482 4271
rect -20448 4237 -20432 4271
rect -20498 4203 -20432 4237
rect -20498 4169 -20482 4203
rect -20448 4169 -20432 4203
rect -20498 4135 -20432 4169
rect -20498 4101 -20482 4135
rect -20448 4101 -20432 4135
rect -20498 4067 -20432 4101
rect -20498 4033 -20482 4067
rect -20448 4033 -20432 4067
rect -20498 3999 -20432 4033
rect -20498 3965 -20482 3999
rect -20448 3965 -20432 3999
rect -20498 3931 -20432 3965
rect -20498 3897 -20482 3931
rect -20448 3897 -20432 3931
rect -20498 3863 -20432 3897
rect -20498 3829 -20482 3863
rect -20448 3829 -20432 3863
rect -20498 3795 -20432 3829
rect -20498 3761 -20482 3795
rect -20448 3761 -20432 3795
rect -20498 3727 -20432 3761
rect -20498 3693 -20482 3727
rect -20448 3693 -20432 3727
rect -20498 3659 -20432 3693
rect -20498 3625 -20482 3659
rect -20448 3625 -20432 3659
rect -20498 3591 -20432 3625
rect -20498 3557 -20482 3591
rect -20448 3557 -20432 3591
rect -20498 3523 -20432 3557
rect -20498 3489 -20482 3523
rect -20448 3489 -20432 3523
rect -20498 3448 -20432 3489
rect -20402 4407 -20336 4448
rect -20402 4373 -20386 4407
rect -20352 4373 -20336 4407
rect -20402 4339 -20336 4373
rect -20402 4305 -20386 4339
rect -20352 4305 -20336 4339
rect -20402 4271 -20336 4305
rect -20402 4237 -20386 4271
rect -20352 4237 -20336 4271
rect -20402 4203 -20336 4237
rect -20402 4169 -20386 4203
rect -20352 4169 -20336 4203
rect -20402 4135 -20336 4169
rect -20402 4101 -20386 4135
rect -20352 4101 -20336 4135
rect -20402 4067 -20336 4101
rect -20402 4033 -20386 4067
rect -20352 4033 -20336 4067
rect -20402 3999 -20336 4033
rect -20402 3965 -20386 3999
rect -20352 3965 -20336 3999
rect -20402 3931 -20336 3965
rect -20402 3897 -20386 3931
rect -20352 3897 -20336 3931
rect -20402 3863 -20336 3897
rect -20402 3829 -20386 3863
rect -20352 3829 -20336 3863
rect -20402 3795 -20336 3829
rect -20402 3761 -20386 3795
rect -20352 3761 -20336 3795
rect -20402 3727 -20336 3761
rect -20402 3693 -20386 3727
rect -20352 3693 -20336 3727
rect -20402 3659 -20336 3693
rect -20402 3625 -20386 3659
rect -20352 3625 -20336 3659
rect -20402 3591 -20336 3625
rect -20402 3557 -20386 3591
rect -20352 3557 -20336 3591
rect -20402 3523 -20336 3557
rect -20402 3489 -20386 3523
rect -20352 3489 -20336 3523
rect -20402 3448 -20336 3489
rect -20306 4407 -20240 4448
rect -20306 4373 -20290 4407
rect -20256 4373 -20240 4407
rect -20306 4339 -20240 4373
rect -20306 4305 -20290 4339
rect -20256 4305 -20240 4339
rect -20306 4271 -20240 4305
rect -20306 4237 -20290 4271
rect -20256 4237 -20240 4271
rect -20306 4203 -20240 4237
rect -20306 4169 -20290 4203
rect -20256 4169 -20240 4203
rect -20306 4135 -20240 4169
rect -20306 4101 -20290 4135
rect -20256 4101 -20240 4135
rect -20306 4067 -20240 4101
rect -20306 4033 -20290 4067
rect -20256 4033 -20240 4067
rect -20306 3999 -20240 4033
rect -20306 3965 -20290 3999
rect -20256 3965 -20240 3999
rect -20306 3931 -20240 3965
rect -20306 3897 -20290 3931
rect -20256 3897 -20240 3931
rect -20306 3863 -20240 3897
rect -20306 3829 -20290 3863
rect -20256 3829 -20240 3863
rect -20306 3795 -20240 3829
rect -20306 3761 -20290 3795
rect -20256 3761 -20240 3795
rect -20306 3727 -20240 3761
rect -20306 3693 -20290 3727
rect -20256 3693 -20240 3727
rect -20306 3659 -20240 3693
rect -20306 3625 -20290 3659
rect -20256 3625 -20240 3659
rect -20306 3591 -20240 3625
rect -20306 3557 -20290 3591
rect -20256 3557 -20240 3591
rect -20306 3523 -20240 3557
rect -20306 3489 -20290 3523
rect -20256 3489 -20240 3523
rect -20306 3448 -20240 3489
rect -20210 4407 -20144 4448
rect -20210 4373 -20194 4407
rect -20160 4373 -20144 4407
rect -20210 4339 -20144 4373
rect -20210 4305 -20194 4339
rect -20160 4305 -20144 4339
rect -20210 4271 -20144 4305
rect -20210 4237 -20194 4271
rect -20160 4237 -20144 4271
rect -20210 4203 -20144 4237
rect -20210 4169 -20194 4203
rect -20160 4169 -20144 4203
rect -20210 4135 -20144 4169
rect -20210 4101 -20194 4135
rect -20160 4101 -20144 4135
rect -20210 4067 -20144 4101
rect -20210 4033 -20194 4067
rect -20160 4033 -20144 4067
rect -20210 3999 -20144 4033
rect -20210 3965 -20194 3999
rect -20160 3965 -20144 3999
rect -20210 3931 -20144 3965
rect -20210 3897 -20194 3931
rect -20160 3897 -20144 3931
rect -20210 3863 -20144 3897
rect -20210 3829 -20194 3863
rect -20160 3829 -20144 3863
rect -20210 3795 -20144 3829
rect -20210 3761 -20194 3795
rect -20160 3761 -20144 3795
rect -20210 3727 -20144 3761
rect -20210 3693 -20194 3727
rect -20160 3693 -20144 3727
rect -20210 3659 -20144 3693
rect -20210 3625 -20194 3659
rect -20160 3625 -20144 3659
rect -20210 3591 -20144 3625
rect -20210 3557 -20194 3591
rect -20160 3557 -20144 3591
rect -20210 3523 -20144 3557
rect -20210 3489 -20194 3523
rect -20160 3489 -20144 3523
rect -20210 3448 -20144 3489
rect -20114 4407 -20048 4448
rect -20114 4373 -20098 4407
rect -20064 4373 -20048 4407
rect -20114 4339 -20048 4373
rect -20114 4305 -20098 4339
rect -20064 4305 -20048 4339
rect -20114 4271 -20048 4305
rect -20114 4237 -20098 4271
rect -20064 4237 -20048 4271
rect -20114 4203 -20048 4237
rect -20114 4169 -20098 4203
rect -20064 4169 -20048 4203
rect -20114 4135 -20048 4169
rect -20114 4101 -20098 4135
rect -20064 4101 -20048 4135
rect -20114 4067 -20048 4101
rect -20114 4033 -20098 4067
rect -20064 4033 -20048 4067
rect -20114 3999 -20048 4033
rect -20114 3965 -20098 3999
rect -20064 3965 -20048 3999
rect -20114 3931 -20048 3965
rect -20114 3897 -20098 3931
rect -20064 3897 -20048 3931
rect -20114 3863 -20048 3897
rect -20114 3829 -20098 3863
rect -20064 3829 -20048 3863
rect -20114 3795 -20048 3829
rect -20114 3761 -20098 3795
rect -20064 3761 -20048 3795
rect -20114 3727 -20048 3761
rect -20114 3693 -20098 3727
rect -20064 3693 -20048 3727
rect -20114 3659 -20048 3693
rect -20114 3625 -20098 3659
rect -20064 3625 -20048 3659
rect -20114 3591 -20048 3625
rect -20114 3557 -20098 3591
rect -20064 3557 -20048 3591
rect -20114 3523 -20048 3557
rect -20114 3489 -20098 3523
rect -20064 3489 -20048 3523
rect -20114 3448 -20048 3489
rect -20018 4407 -19956 4448
rect -20018 4373 -20002 4407
rect -19968 4373 -19956 4407
rect -20018 4339 -19956 4373
rect -20018 4305 -20002 4339
rect -19968 4305 -19956 4339
rect -20018 4271 -19956 4305
rect -20018 4237 -20002 4271
rect -19968 4237 -19956 4271
rect -20018 4203 -19956 4237
rect -20018 4169 -20002 4203
rect -19968 4169 -19956 4203
rect -20018 4135 -19956 4169
rect -20018 4101 -20002 4135
rect -19968 4101 -19956 4135
rect -20018 4067 -19956 4101
rect -20018 4033 -20002 4067
rect -19968 4033 -19956 4067
rect -20018 3999 -19956 4033
rect -20018 3965 -20002 3999
rect -19968 3965 -19956 3999
rect -20018 3931 -19956 3965
rect -20018 3897 -20002 3931
rect -19968 3897 -19956 3931
rect -20018 3863 -19956 3897
rect -20018 3829 -20002 3863
rect -19968 3829 -19956 3863
rect -20018 3795 -19956 3829
rect -20018 3761 -20002 3795
rect -19968 3761 -19956 3795
rect -20018 3727 -19956 3761
rect -20018 3693 -20002 3727
rect -19968 3693 -19956 3727
rect -20018 3659 -19956 3693
rect -20018 3625 -20002 3659
rect -19968 3625 -19956 3659
rect -20018 3591 -19956 3625
rect -20018 3557 -20002 3591
rect -19968 3557 -19956 3591
rect -20018 3523 -19956 3557
rect -20018 3489 -20002 3523
rect -19968 3489 -19956 3523
rect -20018 3448 -19956 3489
rect -19770 4413 -19708 4454
rect -19770 4379 -19758 4413
rect -19724 4379 -19708 4413
rect -19770 4345 -19708 4379
rect -19770 4311 -19758 4345
rect -19724 4311 -19708 4345
rect -19770 4277 -19708 4311
rect -19770 4243 -19758 4277
rect -19724 4243 -19708 4277
rect -19770 4209 -19708 4243
rect -19770 4175 -19758 4209
rect -19724 4175 -19708 4209
rect -19770 4141 -19708 4175
rect -19770 4107 -19758 4141
rect -19724 4107 -19708 4141
rect -19770 4073 -19708 4107
rect -19770 4039 -19758 4073
rect -19724 4039 -19708 4073
rect -19770 4005 -19708 4039
rect -19770 3971 -19758 4005
rect -19724 3971 -19708 4005
rect -19770 3937 -19708 3971
rect -19770 3903 -19758 3937
rect -19724 3903 -19708 3937
rect -19770 3869 -19708 3903
rect -19770 3835 -19758 3869
rect -19724 3835 -19708 3869
rect -19770 3801 -19708 3835
rect -19770 3767 -19758 3801
rect -19724 3767 -19708 3801
rect -19770 3733 -19708 3767
rect -19770 3699 -19758 3733
rect -19724 3699 -19708 3733
rect -19770 3665 -19708 3699
rect -19770 3631 -19758 3665
rect -19724 3631 -19708 3665
rect -19770 3597 -19708 3631
rect -19770 3563 -19758 3597
rect -19724 3563 -19708 3597
rect -19770 3529 -19708 3563
rect -19770 3495 -19758 3529
rect -19724 3495 -19708 3529
rect -19770 3454 -19708 3495
rect -19678 4413 -19612 4454
rect -19678 4379 -19662 4413
rect -19628 4379 -19612 4413
rect -19678 4345 -19612 4379
rect -19678 4311 -19662 4345
rect -19628 4311 -19612 4345
rect -19678 4277 -19612 4311
rect -19678 4243 -19662 4277
rect -19628 4243 -19612 4277
rect -19678 4209 -19612 4243
rect -19678 4175 -19662 4209
rect -19628 4175 -19612 4209
rect -19678 4141 -19612 4175
rect -19678 4107 -19662 4141
rect -19628 4107 -19612 4141
rect -19678 4073 -19612 4107
rect -19678 4039 -19662 4073
rect -19628 4039 -19612 4073
rect -19678 4005 -19612 4039
rect -19678 3971 -19662 4005
rect -19628 3971 -19612 4005
rect -19678 3937 -19612 3971
rect -19678 3903 -19662 3937
rect -19628 3903 -19612 3937
rect -19678 3869 -19612 3903
rect -19678 3835 -19662 3869
rect -19628 3835 -19612 3869
rect -19678 3801 -19612 3835
rect -19678 3767 -19662 3801
rect -19628 3767 -19612 3801
rect -19678 3733 -19612 3767
rect -19678 3699 -19662 3733
rect -19628 3699 -19612 3733
rect -19678 3665 -19612 3699
rect -19678 3631 -19662 3665
rect -19628 3631 -19612 3665
rect -19678 3597 -19612 3631
rect -19678 3563 -19662 3597
rect -19628 3563 -19612 3597
rect -19678 3529 -19612 3563
rect -19678 3495 -19662 3529
rect -19628 3495 -19612 3529
rect -19678 3454 -19612 3495
rect -19582 4413 -19516 4454
rect -19582 4379 -19566 4413
rect -19532 4379 -19516 4413
rect -19582 4345 -19516 4379
rect -19582 4311 -19566 4345
rect -19532 4311 -19516 4345
rect -19582 4277 -19516 4311
rect -19582 4243 -19566 4277
rect -19532 4243 -19516 4277
rect -19582 4209 -19516 4243
rect -19582 4175 -19566 4209
rect -19532 4175 -19516 4209
rect -19582 4141 -19516 4175
rect -19582 4107 -19566 4141
rect -19532 4107 -19516 4141
rect -19582 4073 -19516 4107
rect -19582 4039 -19566 4073
rect -19532 4039 -19516 4073
rect -19582 4005 -19516 4039
rect -19582 3971 -19566 4005
rect -19532 3971 -19516 4005
rect -19582 3937 -19516 3971
rect -19582 3903 -19566 3937
rect -19532 3903 -19516 3937
rect -19582 3869 -19516 3903
rect -19582 3835 -19566 3869
rect -19532 3835 -19516 3869
rect -19582 3801 -19516 3835
rect -19582 3767 -19566 3801
rect -19532 3767 -19516 3801
rect -19582 3733 -19516 3767
rect -19582 3699 -19566 3733
rect -19532 3699 -19516 3733
rect -19582 3665 -19516 3699
rect -19582 3631 -19566 3665
rect -19532 3631 -19516 3665
rect -19582 3597 -19516 3631
rect -19582 3563 -19566 3597
rect -19532 3563 -19516 3597
rect -19582 3529 -19516 3563
rect -19582 3495 -19566 3529
rect -19532 3495 -19516 3529
rect -19582 3454 -19516 3495
rect -19486 4413 -19420 4454
rect -19486 4379 -19470 4413
rect -19436 4379 -19420 4413
rect -19486 4345 -19420 4379
rect -19486 4311 -19470 4345
rect -19436 4311 -19420 4345
rect -19486 4277 -19420 4311
rect -19486 4243 -19470 4277
rect -19436 4243 -19420 4277
rect -19486 4209 -19420 4243
rect -19486 4175 -19470 4209
rect -19436 4175 -19420 4209
rect -19486 4141 -19420 4175
rect -19486 4107 -19470 4141
rect -19436 4107 -19420 4141
rect -19486 4073 -19420 4107
rect -19486 4039 -19470 4073
rect -19436 4039 -19420 4073
rect -19486 4005 -19420 4039
rect -19486 3971 -19470 4005
rect -19436 3971 -19420 4005
rect -19486 3937 -19420 3971
rect -19486 3903 -19470 3937
rect -19436 3903 -19420 3937
rect -19486 3869 -19420 3903
rect -19486 3835 -19470 3869
rect -19436 3835 -19420 3869
rect -19486 3801 -19420 3835
rect -19486 3767 -19470 3801
rect -19436 3767 -19420 3801
rect -19486 3733 -19420 3767
rect -19486 3699 -19470 3733
rect -19436 3699 -19420 3733
rect -19486 3665 -19420 3699
rect -19486 3631 -19470 3665
rect -19436 3631 -19420 3665
rect -19486 3597 -19420 3631
rect -19486 3563 -19470 3597
rect -19436 3563 -19420 3597
rect -19486 3529 -19420 3563
rect -19486 3495 -19470 3529
rect -19436 3495 -19420 3529
rect -19486 3454 -19420 3495
rect -19390 4413 -19324 4454
rect -19390 4379 -19374 4413
rect -19340 4379 -19324 4413
rect -19390 4345 -19324 4379
rect -19390 4311 -19374 4345
rect -19340 4311 -19324 4345
rect -19390 4277 -19324 4311
rect -19390 4243 -19374 4277
rect -19340 4243 -19324 4277
rect -19390 4209 -19324 4243
rect -19390 4175 -19374 4209
rect -19340 4175 -19324 4209
rect -19390 4141 -19324 4175
rect -19390 4107 -19374 4141
rect -19340 4107 -19324 4141
rect -19390 4073 -19324 4107
rect -19390 4039 -19374 4073
rect -19340 4039 -19324 4073
rect -19390 4005 -19324 4039
rect -19390 3971 -19374 4005
rect -19340 3971 -19324 4005
rect -19390 3937 -19324 3971
rect -19390 3903 -19374 3937
rect -19340 3903 -19324 3937
rect -19390 3869 -19324 3903
rect -19390 3835 -19374 3869
rect -19340 3835 -19324 3869
rect -19390 3801 -19324 3835
rect -19390 3767 -19374 3801
rect -19340 3767 -19324 3801
rect -19390 3733 -19324 3767
rect -19390 3699 -19374 3733
rect -19340 3699 -19324 3733
rect -19390 3665 -19324 3699
rect -19390 3631 -19374 3665
rect -19340 3631 -19324 3665
rect -19390 3597 -19324 3631
rect -19390 3563 -19374 3597
rect -19340 3563 -19324 3597
rect -19390 3529 -19324 3563
rect -19390 3495 -19374 3529
rect -19340 3495 -19324 3529
rect -19390 3454 -19324 3495
rect -19294 4413 -19228 4454
rect -19294 4379 -19278 4413
rect -19244 4379 -19228 4413
rect -19294 4345 -19228 4379
rect -19294 4311 -19278 4345
rect -19244 4311 -19228 4345
rect -19294 4277 -19228 4311
rect -19294 4243 -19278 4277
rect -19244 4243 -19228 4277
rect -19294 4209 -19228 4243
rect -19294 4175 -19278 4209
rect -19244 4175 -19228 4209
rect -19294 4141 -19228 4175
rect -19294 4107 -19278 4141
rect -19244 4107 -19228 4141
rect -19294 4073 -19228 4107
rect -19294 4039 -19278 4073
rect -19244 4039 -19228 4073
rect -19294 4005 -19228 4039
rect -19294 3971 -19278 4005
rect -19244 3971 -19228 4005
rect -19294 3937 -19228 3971
rect -19294 3903 -19278 3937
rect -19244 3903 -19228 3937
rect -19294 3869 -19228 3903
rect -19294 3835 -19278 3869
rect -19244 3835 -19228 3869
rect -19294 3801 -19228 3835
rect -19294 3767 -19278 3801
rect -19244 3767 -19228 3801
rect -19294 3733 -19228 3767
rect -19294 3699 -19278 3733
rect -19244 3699 -19228 3733
rect -19294 3665 -19228 3699
rect -19294 3631 -19278 3665
rect -19244 3631 -19228 3665
rect -19294 3597 -19228 3631
rect -19294 3563 -19278 3597
rect -19244 3563 -19228 3597
rect -19294 3529 -19228 3563
rect -19294 3495 -19278 3529
rect -19244 3495 -19228 3529
rect -19294 3454 -19228 3495
rect -19198 4413 -19132 4454
rect -19198 4379 -19182 4413
rect -19148 4379 -19132 4413
rect -19198 4345 -19132 4379
rect -19198 4311 -19182 4345
rect -19148 4311 -19132 4345
rect -19198 4277 -19132 4311
rect -19198 4243 -19182 4277
rect -19148 4243 -19132 4277
rect -19198 4209 -19132 4243
rect -19198 4175 -19182 4209
rect -19148 4175 -19132 4209
rect -19198 4141 -19132 4175
rect -19198 4107 -19182 4141
rect -19148 4107 -19132 4141
rect -19198 4073 -19132 4107
rect -19198 4039 -19182 4073
rect -19148 4039 -19132 4073
rect -19198 4005 -19132 4039
rect -19198 3971 -19182 4005
rect -19148 3971 -19132 4005
rect -19198 3937 -19132 3971
rect -19198 3903 -19182 3937
rect -19148 3903 -19132 3937
rect -19198 3869 -19132 3903
rect -19198 3835 -19182 3869
rect -19148 3835 -19132 3869
rect -19198 3801 -19132 3835
rect -19198 3767 -19182 3801
rect -19148 3767 -19132 3801
rect -19198 3733 -19132 3767
rect -19198 3699 -19182 3733
rect -19148 3699 -19132 3733
rect -19198 3665 -19132 3699
rect -19198 3631 -19182 3665
rect -19148 3631 -19132 3665
rect -19198 3597 -19132 3631
rect -19198 3563 -19182 3597
rect -19148 3563 -19132 3597
rect -19198 3529 -19132 3563
rect -19198 3495 -19182 3529
rect -19148 3495 -19132 3529
rect -19198 3454 -19132 3495
rect -19102 4413 -19036 4454
rect -19102 4379 -19086 4413
rect -19052 4379 -19036 4413
rect -19102 4345 -19036 4379
rect -19102 4311 -19086 4345
rect -19052 4311 -19036 4345
rect -19102 4277 -19036 4311
rect -19102 4243 -19086 4277
rect -19052 4243 -19036 4277
rect -19102 4209 -19036 4243
rect -19102 4175 -19086 4209
rect -19052 4175 -19036 4209
rect -19102 4141 -19036 4175
rect -19102 4107 -19086 4141
rect -19052 4107 -19036 4141
rect -19102 4073 -19036 4107
rect -19102 4039 -19086 4073
rect -19052 4039 -19036 4073
rect -19102 4005 -19036 4039
rect -19102 3971 -19086 4005
rect -19052 3971 -19036 4005
rect -19102 3937 -19036 3971
rect -19102 3903 -19086 3937
rect -19052 3903 -19036 3937
rect -19102 3869 -19036 3903
rect -19102 3835 -19086 3869
rect -19052 3835 -19036 3869
rect -19102 3801 -19036 3835
rect -19102 3767 -19086 3801
rect -19052 3767 -19036 3801
rect -19102 3733 -19036 3767
rect -19102 3699 -19086 3733
rect -19052 3699 -19036 3733
rect -19102 3665 -19036 3699
rect -19102 3631 -19086 3665
rect -19052 3631 -19036 3665
rect -19102 3597 -19036 3631
rect -19102 3563 -19086 3597
rect -19052 3563 -19036 3597
rect -19102 3529 -19036 3563
rect -19102 3495 -19086 3529
rect -19052 3495 -19036 3529
rect -19102 3454 -19036 3495
rect -19006 4413 -18940 4454
rect -19006 4379 -18990 4413
rect -18956 4379 -18940 4413
rect -19006 4345 -18940 4379
rect -19006 4311 -18990 4345
rect -18956 4311 -18940 4345
rect -19006 4277 -18940 4311
rect -19006 4243 -18990 4277
rect -18956 4243 -18940 4277
rect -19006 4209 -18940 4243
rect -19006 4175 -18990 4209
rect -18956 4175 -18940 4209
rect -19006 4141 -18940 4175
rect -19006 4107 -18990 4141
rect -18956 4107 -18940 4141
rect -19006 4073 -18940 4107
rect -19006 4039 -18990 4073
rect -18956 4039 -18940 4073
rect -19006 4005 -18940 4039
rect -19006 3971 -18990 4005
rect -18956 3971 -18940 4005
rect -19006 3937 -18940 3971
rect -19006 3903 -18990 3937
rect -18956 3903 -18940 3937
rect -19006 3869 -18940 3903
rect -19006 3835 -18990 3869
rect -18956 3835 -18940 3869
rect -19006 3801 -18940 3835
rect -19006 3767 -18990 3801
rect -18956 3767 -18940 3801
rect -19006 3733 -18940 3767
rect -19006 3699 -18990 3733
rect -18956 3699 -18940 3733
rect -19006 3665 -18940 3699
rect -19006 3631 -18990 3665
rect -18956 3631 -18940 3665
rect -19006 3597 -18940 3631
rect -19006 3563 -18990 3597
rect -18956 3563 -18940 3597
rect -19006 3529 -18940 3563
rect -19006 3495 -18990 3529
rect -18956 3495 -18940 3529
rect -19006 3454 -18940 3495
rect -18910 4413 -18844 4454
rect -18910 4379 -18894 4413
rect -18860 4379 -18844 4413
rect -18910 4345 -18844 4379
rect -18910 4311 -18894 4345
rect -18860 4311 -18844 4345
rect -18910 4277 -18844 4311
rect -18910 4243 -18894 4277
rect -18860 4243 -18844 4277
rect -18910 4209 -18844 4243
rect -18910 4175 -18894 4209
rect -18860 4175 -18844 4209
rect -18910 4141 -18844 4175
rect -18910 4107 -18894 4141
rect -18860 4107 -18844 4141
rect -18910 4073 -18844 4107
rect -18910 4039 -18894 4073
rect -18860 4039 -18844 4073
rect -18910 4005 -18844 4039
rect -18910 3971 -18894 4005
rect -18860 3971 -18844 4005
rect -18910 3937 -18844 3971
rect -18910 3903 -18894 3937
rect -18860 3903 -18844 3937
rect -18910 3869 -18844 3903
rect -18910 3835 -18894 3869
rect -18860 3835 -18844 3869
rect -18910 3801 -18844 3835
rect -18910 3767 -18894 3801
rect -18860 3767 -18844 3801
rect -18910 3733 -18844 3767
rect -18910 3699 -18894 3733
rect -18860 3699 -18844 3733
rect -18910 3665 -18844 3699
rect -18910 3631 -18894 3665
rect -18860 3631 -18844 3665
rect -18910 3597 -18844 3631
rect -18910 3563 -18894 3597
rect -18860 3563 -18844 3597
rect -18910 3529 -18844 3563
rect -18910 3495 -18894 3529
rect -18860 3495 -18844 3529
rect -18910 3454 -18844 3495
rect -18814 4413 -18752 4454
rect -18814 4379 -18798 4413
rect -18764 4379 -18752 4413
rect -18814 4345 -18752 4379
rect -18814 4311 -18798 4345
rect -18764 4311 -18752 4345
rect -18814 4277 -18752 4311
rect -18814 4243 -18798 4277
rect -18764 4243 -18752 4277
rect -18814 4209 -18752 4243
rect -18814 4175 -18798 4209
rect -18764 4175 -18752 4209
rect -18814 4141 -18752 4175
rect -18814 4107 -18798 4141
rect -18764 4107 -18752 4141
rect -18814 4073 -18752 4107
rect -18814 4039 -18798 4073
rect -18764 4039 -18752 4073
rect -18814 4005 -18752 4039
rect -18814 3971 -18798 4005
rect -18764 3971 -18752 4005
rect -18814 3937 -18752 3971
rect -18814 3903 -18798 3937
rect -18764 3903 -18752 3937
rect -18814 3869 -18752 3903
rect -18814 3835 -18798 3869
rect -18764 3835 -18752 3869
rect -18814 3801 -18752 3835
rect -18814 3767 -18798 3801
rect -18764 3767 -18752 3801
rect -18814 3733 -18752 3767
rect -18814 3699 -18798 3733
rect -18764 3699 -18752 3733
rect -18814 3665 -18752 3699
rect -18814 3631 -18798 3665
rect -18764 3631 -18752 3665
rect -18814 3597 -18752 3631
rect -18814 3563 -18798 3597
rect -18764 3563 -18752 3597
rect -18814 3529 -18752 3563
rect -18814 3495 -18798 3529
rect -18764 3495 -18752 3529
rect -18814 3454 -18752 3495
rect -18602 4415 -18540 4456
rect -18602 4381 -18590 4415
rect -18556 4381 -18540 4415
rect -18602 4347 -18540 4381
rect -18602 4313 -18590 4347
rect -18556 4313 -18540 4347
rect -18602 4279 -18540 4313
rect -18602 4245 -18590 4279
rect -18556 4245 -18540 4279
rect -18602 4211 -18540 4245
rect -18602 4177 -18590 4211
rect -18556 4177 -18540 4211
rect -18602 4143 -18540 4177
rect -18602 4109 -18590 4143
rect -18556 4109 -18540 4143
rect -18602 4075 -18540 4109
rect -18602 4041 -18590 4075
rect -18556 4041 -18540 4075
rect -18602 4007 -18540 4041
rect -18602 3973 -18590 4007
rect -18556 3973 -18540 4007
rect -18602 3939 -18540 3973
rect -18602 3905 -18590 3939
rect -18556 3905 -18540 3939
rect -18602 3871 -18540 3905
rect -18602 3837 -18590 3871
rect -18556 3837 -18540 3871
rect -18602 3803 -18540 3837
rect -18602 3769 -18590 3803
rect -18556 3769 -18540 3803
rect -18602 3735 -18540 3769
rect -18602 3701 -18590 3735
rect -18556 3701 -18540 3735
rect -18602 3667 -18540 3701
rect -18602 3633 -18590 3667
rect -18556 3633 -18540 3667
rect -18602 3599 -18540 3633
rect -18602 3565 -18590 3599
rect -18556 3565 -18540 3599
rect -18602 3531 -18540 3565
rect -18602 3497 -18590 3531
rect -18556 3497 -18540 3531
rect -18602 3456 -18540 3497
rect -18510 4415 -18444 4456
rect -18510 4381 -18494 4415
rect -18460 4381 -18444 4415
rect -18510 4347 -18444 4381
rect -18510 4313 -18494 4347
rect -18460 4313 -18444 4347
rect -18510 4279 -18444 4313
rect -18510 4245 -18494 4279
rect -18460 4245 -18444 4279
rect -18510 4211 -18444 4245
rect -18510 4177 -18494 4211
rect -18460 4177 -18444 4211
rect -18510 4143 -18444 4177
rect -18510 4109 -18494 4143
rect -18460 4109 -18444 4143
rect -18510 4075 -18444 4109
rect -18510 4041 -18494 4075
rect -18460 4041 -18444 4075
rect -18510 4007 -18444 4041
rect -18510 3973 -18494 4007
rect -18460 3973 -18444 4007
rect -18510 3939 -18444 3973
rect -18510 3905 -18494 3939
rect -18460 3905 -18444 3939
rect -18510 3871 -18444 3905
rect -18510 3837 -18494 3871
rect -18460 3837 -18444 3871
rect -18510 3803 -18444 3837
rect -18510 3769 -18494 3803
rect -18460 3769 -18444 3803
rect -18510 3735 -18444 3769
rect -18510 3701 -18494 3735
rect -18460 3701 -18444 3735
rect -18510 3667 -18444 3701
rect -18510 3633 -18494 3667
rect -18460 3633 -18444 3667
rect -18510 3599 -18444 3633
rect -18510 3565 -18494 3599
rect -18460 3565 -18444 3599
rect -18510 3531 -18444 3565
rect -18510 3497 -18494 3531
rect -18460 3497 -18444 3531
rect -18510 3456 -18444 3497
rect -18414 4415 -18348 4456
rect -18414 4381 -18398 4415
rect -18364 4381 -18348 4415
rect -18414 4347 -18348 4381
rect -18414 4313 -18398 4347
rect -18364 4313 -18348 4347
rect -18414 4279 -18348 4313
rect -18414 4245 -18398 4279
rect -18364 4245 -18348 4279
rect -18414 4211 -18348 4245
rect -18414 4177 -18398 4211
rect -18364 4177 -18348 4211
rect -18414 4143 -18348 4177
rect -18414 4109 -18398 4143
rect -18364 4109 -18348 4143
rect -18414 4075 -18348 4109
rect -18414 4041 -18398 4075
rect -18364 4041 -18348 4075
rect -18414 4007 -18348 4041
rect -18414 3973 -18398 4007
rect -18364 3973 -18348 4007
rect -18414 3939 -18348 3973
rect -18414 3905 -18398 3939
rect -18364 3905 -18348 3939
rect -18414 3871 -18348 3905
rect -18414 3837 -18398 3871
rect -18364 3837 -18348 3871
rect -18414 3803 -18348 3837
rect -18414 3769 -18398 3803
rect -18364 3769 -18348 3803
rect -18414 3735 -18348 3769
rect -18414 3701 -18398 3735
rect -18364 3701 -18348 3735
rect -18414 3667 -18348 3701
rect -18414 3633 -18398 3667
rect -18364 3633 -18348 3667
rect -18414 3599 -18348 3633
rect -18414 3565 -18398 3599
rect -18364 3565 -18348 3599
rect -18414 3531 -18348 3565
rect -18414 3497 -18398 3531
rect -18364 3497 -18348 3531
rect -18414 3456 -18348 3497
rect -18318 4415 -18252 4456
rect -18318 4381 -18302 4415
rect -18268 4381 -18252 4415
rect -18318 4347 -18252 4381
rect -18318 4313 -18302 4347
rect -18268 4313 -18252 4347
rect -18318 4279 -18252 4313
rect -18318 4245 -18302 4279
rect -18268 4245 -18252 4279
rect -18318 4211 -18252 4245
rect -18318 4177 -18302 4211
rect -18268 4177 -18252 4211
rect -18318 4143 -18252 4177
rect -18318 4109 -18302 4143
rect -18268 4109 -18252 4143
rect -18318 4075 -18252 4109
rect -18318 4041 -18302 4075
rect -18268 4041 -18252 4075
rect -18318 4007 -18252 4041
rect -18318 3973 -18302 4007
rect -18268 3973 -18252 4007
rect -18318 3939 -18252 3973
rect -18318 3905 -18302 3939
rect -18268 3905 -18252 3939
rect -18318 3871 -18252 3905
rect -18318 3837 -18302 3871
rect -18268 3837 -18252 3871
rect -18318 3803 -18252 3837
rect -18318 3769 -18302 3803
rect -18268 3769 -18252 3803
rect -18318 3735 -18252 3769
rect -18318 3701 -18302 3735
rect -18268 3701 -18252 3735
rect -18318 3667 -18252 3701
rect -18318 3633 -18302 3667
rect -18268 3633 -18252 3667
rect -18318 3599 -18252 3633
rect -18318 3565 -18302 3599
rect -18268 3565 -18252 3599
rect -18318 3531 -18252 3565
rect -18318 3497 -18302 3531
rect -18268 3497 -18252 3531
rect -18318 3456 -18252 3497
rect -18222 4415 -18156 4456
rect -18222 4381 -18206 4415
rect -18172 4381 -18156 4415
rect -18222 4347 -18156 4381
rect -18222 4313 -18206 4347
rect -18172 4313 -18156 4347
rect -18222 4279 -18156 4313
rect -18222 4245 -18206 4279
rect -18172 4245 -18156 4279
rect -18222 4211 -18156 4245
rect -18222 4177 -18206 4211
rect -18172 4177 -18156 4211
rect -18222 4143 -18156 4177
rect -18222 4109 -18206 4143
rect -18172 4109 -18156 4143
rect -18222 4075 -18156 4109
rect -18222 4041 -18206 4075
rect -18172 4041 -18156 4075
rect -18222 4007 -18156 4041
rect -18222 3973 -18206 4007
rect -18172 3973 -18156 4007
rect -18222 3939 -18156 3973
rect -18222 3905 -18206 3939
rect -18172 3905 -18156 3939
rect -18222 3871 -18156 3905
rect -18222 3837 -18206 3871
rect -18172 3837 -18156 3871
rect -18222 3803 -18156 3837
rect -18222 3769 -18206 3803
rect -18172 3769 -18156 3803
rect -18222 3735 -18156 3769
rect -18222 3701 -18206 3735
rect -18172 3701 -18156 3735
rect -18222 3667 -18156 3701
rect -18222 3633 -18206 3667
rect -18172 3633 -18156 3667
rect -18222 3599 -18156 3633
rect -18222 3565 -18206 3599
rect -18172 3565 -18156 3599
rect -18222 3531 -18156 3565
rect -18222 3497 -18206 3531
rect -18172 3497 -18156 3531
rect -18222 3456 -18156 3497
rect -18126 4415 -18064 4456
rect 1472 4495 1534 4529
rect -18126 4381 -18110 4415
rect -18076 4381 -18064 4415
rect -18126 4347 -18064 4381
rect -18126 4313 -18110 4347
rect -18076 4313 -18064 4347
rect -18126 4279 -18064 4313
rect -18126 4245 -18110 4279
rect -18076 4245 -18064 4279
rect -18126 4211 -18064 4245
rect -18126 4177 -18110 4211
rect -18076 4177 -18064 4211
rect -18126 4143 -18064 4177
rect -18126 4109 -18110 4143
rect -18076 4109 -18064 4143
rect -18126 4075 -18064 4109
rect -18126 4041 -18110 4075
rect -18076 4041 -18064 4075
rect -18126 4007 -18064 4041
rect -18126 3973 -18110 4007
rect -18076 3973 -18064 4007
rect -18126 3939 -18064 3973
rect -18126 3905 -18110 3939
rect -18076 3905 -18064 3939
rect -18126 3871 -18064 3905
rect -18126 3837 -18110 3871
rect -18076 3837 -18064 3871
rect -18126 3803 -18064 3837
rect -18126 3769 -18110 3803
rect -18076 3769 -18064 3803
rect -18126 3735 -18064 3769
rect -18126 3701 -18110 3735
rect -18076 3701 -18064 3735
rect -18126 3667 -18064 3701
rect -18126 3633 -18110 3667
rect -18076 3633 -18064 3667
rect -18126 3599 -18064 3633
rect -18126 3565 -18110 3599
rect -18076 3565 -18064 3599
rect -18126 3531 -18064 3565
rect -18126 3497 -18110 3531
rect -18076 3497 -18064 3531
rect -18126 3456 -18064 3497
rect -16768 4413 -16706 4454
rect -16768 4379 -16756 4413
rect -16722 4379 -16706 4413
rect -16768 4345 -16706 4379
rect -16768 4311 -16756 4345
rect -16722 4311 -16706 4345
rect -16768 4277 -16706 4311
rect -16768 4243 -16756 4277
rect -16722 4243 -16706 4277
rect -16768 4209 -16706 4243
rect -16768 4175 -16756 4209
rect -16722 4175 -16706 4209
rect -16768 4141 -16706 4175
rect -16768 4107 -16756 4141
rect -16722 4107 -16706 4141
rect -16768 4073 -16706 4107
rect -16768 4039 -16756 4073
rect -16722 4039 -16706 4073
rect -16768 4005 -16706 4039
rect -16768 3971 -16756 4005
rect -16722 3971 -16706 4005
rect -16768 3937 -16706 3971
rect -16768 3903 -16756 3937
rect -16722 3903 -16706 3937
rect -16768 3869 -16706 3903
rect -16768 3835 -16756 3869
rect -16722 3835 -16706 3869
rect -16768 3801 -16706 3835
rect -16768 3767 -16756 3801
rect -16722 3767 -16706 3801
rect -16768 3733 -16706 3767
rect -16768 3699 -16756 3733
rect -16722 3699 -16706 3733
rect -16768 3665 -16706 3699
rect -16768 3631 -16756 3665
rect -16722 3631 -16706 3665
rect -16768 3597 -16706 3631
rect -16768 3563 -16756 3597
rect -16722 3563 -16706 3597
rect -16768 3529 -16706 3563
rect -16768 3495 -16756 3529
rect -16722 3495 -16706 3529
rect -16768 3454 -16706 3495
rect -16676 4413 -16610 4454
rect -16676 4379 -16660 4413
rect -16626 4379 -16610 4413
rect -16676 4345 -16610 4379
rect -16676 4311 -16660 4345
rect -16626 4311 -16610 4345
rect -16676 4277 -16610 4311
rect -16676 4243 -16660 4277
rect -16626 4243 -16610 4277
rect -16676 4209 -16610 4243
rect -16676 4175 -16660 4209
rect -16626 4175 -16610 4209
rect -16676 4141 -16610 4175
rect -16676 4107 -16660 4141
rect -16626 4107 -16610 4141
rect -16676 4073 -16610 4107
rect -16676 4039 -16660 4073
rect -16626 4039 -16610 4073
rect -16676 4005 -16610 4039
rect -16676 3971 -16660 4005
rect -16626 3971 -16610 4005
rect -16676 3937 -16610 3971
rect -16676 3903 -16660 3937
rect -16626 3903 -16610 3937
rect -16676 3869 -16610 3903
rect -16676 3835 -16660 3869
rect -16626 3835 -16610 3869
rect -16676 3801 -16610 3835
rect -16676 3767 -16660 3801
rect -16626 3767 -16610 3801
rect -16676 3733 -16610 3767
rect -16676 3699 -16660 3733
rect -16626 3699 -16610 3733
rect -16676 3665 -16610 3699
rect -16676 3631 -16660 3665
rect -16626 3631 -16610 3665
rect -16676 3597 -16610 3631
rect -16676 3563 -16660 3597
rect -16626 3563 -16610 3597
rect -16676 3529 -16610 3563
rect -16676 3495 -16660 3529
rect -16626 3495 -16610 3529
rect -16676 3454 -16610 3495
rect -16580 4413 -16514 4454
rect -16580 4379 -16564 4413
rect -16530 4379 -16514 4413
rect -16580 4345 -16514 4379
rect -16580 4311 -16564 4345
rect -16530 4311 -16514 4345
rect -16580 4277 -16514 4311
rect -16580 4243 -16564 4277
rect -16530 4243 -16514 4277
rect -16580 4209 -16514 4243
rect -16580 4175 -16564 4209
rect -16530 4175 -16514 4209
rect -16580 4141 -16514 4175
rect -16580 4107 -16564 4141
rect -16530 4107 -16514 4141
rect -16580 4073 -16514 4107
rect -16580 4039 -16564 4073
rect -16530 4039 -16514 4073
rect -16580 4005 -16514 4039
rect -16580 3971 -16564 4005
rect -16530 3971 -16514 4005
rect -16580 3937 -16514 3971
rect -16580 3903 -16564 3937
rect -16530 3903 -16514 3937
rect -16580 3869 -16514 3903
rect -16580 3835 -16564 3869
rect -16530 3835 -16514 3869
rect -16580 3801 -16514 3835
rect -16580 3767 -16564 3801
rect -16530 3767 -16514 3801
rect -16580 3733 -16514 3767
rect -16580 3699 -16564 3733
rect -16530 3699 -16514 3733
rect -16580 3665 -16514 3699
rect -16580 3631 -16564 3665
rect -16530 3631 -16514 3665
rect -16580 3597 -16514 3631
rect -16580 3563 -16564 3597
rect -16530 3563 -16514 3597
rect -16580 3529 -16514 3563
rect -16580 3495 -16564 3529
rect -16530 3495 -16514 3529
rect -16580 3454 -16514 3495
rect -16484 4413 -16418 4454
rect -16484 4379 -16468 4413
rect -16434 4379 -16418 4413
rect -16484 4345 -16418 4379
rect -16484 4311 -16468 4345
rect -16434 4311 -16418 4345
rect -16484 4277 -16418 4311
rect -16484 4243 -16468 4277
rect -16434 4243 -16418 4277
rect -16484 4209 -16418 4243
rect -16484 4175 -16468 4209
rect -16434 4175 -16418 4209
rect -16484 4141 -16418 4175
rect -16484 4107 -16468 4141
rect -16434 4107 -16418 4141
rect -16484 4073 -16418 4107
rect -16484 4039 -16468 4073
rect -16434 4039 -16418 4073
rect -16484 4005 -16418 4039
rect -16484 3971 -16468 4005
rect -16434 3971 -16418 4005
rect -16484 3937 -16418 3971
rect -16484 3903 -16468 3937
rect -16434 3903 -16418 3937
rect -16484 3869 -16418 3903
rect -16484 3835 -16468 3869
rect -16434 3835 -16418 3869
rect -16484 3801 -16418 3835
rect -16484 3767 -16468 3801
rect -16434 3767 -16418 3801
rect -16484 3733 -16418 3767
rect -16484 3699 -16468 3733
rect -16434 3699 -16418 3733
rect -16484 3665 -16418 3699
rect -16484 3631 -16468 3665
rect -16434 3631 -16418 3665
rect -16484 3597 -16418 3631
rect -16484 3563 -16468 3597
rect -16434 3563 -16418 3597
rect -16484 3529 -16418 3563
rect -16484 3495 -16468 3529
rect -16434 3495 -16418 3529
rect -16484 3454 -16418 3495
rect -16388 4413 -16322 4454
rect -16388 4379 -16372 4413
rect -16338 4379 -16322 4413
rect -16388 4345 -16322 4379
rect -16388 4311 -16372 4345
rect -16338 4311 -16322 4345
rect -16388 4277 -16322 4311
rect -16388 4243 -16372 4277
rect -16338 4243 -16322 4277
rect -16388 4209 -16322 4243
rect -16388 4175 -16372 4209
rect -16338 4175 -16322 4209
rect -16388 4141 -16322 4175
rect -16388 4107 -16372 4141
rect -16338 4107 -16322 4141
rect -16388 4073 -16322 4107
rect -16388 4039 -16372 4073
rect -16338 4039 -16322 4073
rect -16388 4005 -16322 4039
rect -16388 3971 -16372 4005
rect -16338 3971 -16322 4005
rect -16388 3937 -16322 3971
rect -16388 3903 -16372 3937
rect -16338 3903 -16322 3937
rect -16388 3869 -16322 3903
rect -16388 3835 -16372 3869
rect -16338 3835 -16322 3869
rect -16388 3801 -16322 3835
rect -16388 3767 -16372 3801
rect -16338 3767 -16322 3801
rect -16388 3733 -16322 3767
rect -16388 3699 -16372 3733
rect -16338 3699 -16322 3733
rect -16388 3665 -16322 3699
rect -16388 3631 -16372 3665
rect -16338 3631 -16322 3665
rect -16388 3597 -16322 3631
rect -16388 3563 -16372 3597
rect -16338 3563 -16322 3597
rect -16388 3529 -16322 3563
rect -16388 3495 -16372 3529
rect -16338 3495 -16322 3529
rect -16388 3454 -16322 3495
rect -16292 4413 -16226 4454
rect -16292 4379 -16276 4413
rect -16242 4379 -16226 4413
rect -16292 4345 -16226 4379
rect -16292 4311 -16276 4345
rect -16242 4311 -16226 4345
rect -16292 4277 -16226 4311
rect -16292 4243 -16276 4277
rect -16242 4243 -16226 4277
rect -16292 4209 -16226 4243
rect -16292 4175 -16276 4209
rect -16242 4175 -16226 4209
rect -16292 4141 -16226 4175
rect -16292 4107 -16276 4141
rect -16242 4107 -16226 4141
rect -16292 4073 -16226 4107
rect -16292 4039 -16276 4073
rect -16242 4039 -16226 4073
rect -16292 4005 -16226 4039
rect -16292 3971 -16276 4005
rect -16242 3971 -16226 4005
rect -16292 3937 -16226 3971
rect -16292 3903 -16276 3937
rect -16242 3903 -16226 3937
rect -16292 3869 -16226 3903
rect -16292 3835 -16276 3869
rect -16242 3835 -16226 3869
rect -16292 3801 -16226 3835
rect -16292 3767 -16276 3801
rect -16242 3767 -16226 3801
rect -16292 3733 -16226 3767
rect -16292 3699 -16276 3733
rect -16242 3699 -16226 3733
rect -16292 3665 -16226 3699
rect -16292 3631 -16276 3665
rect -16242 3631 -16226 3665
rect -16292 3597 -16226 3631
rect -16292 3563 -16276 3597
rect -16242 3563 -16226 3597
rect -16292 3529 -16226 3563
rect -16292 3495 -16276 3529
rect -16242 3495 -16226 3529
rect -16292 3454 -16226 3495
rect -16196 4413 -16130 4454
rect -16196 4379 -16180 4413
rect -16146 4379 -16130 4413
rect -16196 4345 -16130 4379
rect -16196 4311 -16180 4345
rect -16146 4311 -16130 4345
rect -16196 4277 -16130 4311
rect -16196 4243 -16180 4277
rect -16146 4243 -16130 4277
rect -16196 4209 -16130 4243
rect -16196 4175 -16180 4209
rect -16146 4175 -16130 4209
rect -16196 4141 -16130 4175
rect -16196 4107 -16180 4141
rect -16146 4107 -16130 4141
rect -16196 4073 -16130 4107
rect -16196 4039 -16180 4073
rect -16146 4039 -16130 4073
rect -16196 4005 -16130 4039
rect -16196 3971 -16180 4005
rect -16146 3971 -16130 4005
rect -16196 3937 -16130 3971
rect -16196 3903 -16180 3937
rect -16146 3903 -16130 3937
rect -16196 3869 -16130 3903
rect -16196 3835 -16180 3869
rect -16146 3835 -16130 3869
rect -16196 3801 -16130 3835
rect -16196 3767 -16180 3801
rect -16146 3767 -16130 3801
rect -16196 3733 -16130 3767
rect -16196 3699 -16180 3733
rect -16146 3699 -16130 3733
rect -16196 3665 -16130 3699
rect -16196 3631 -16180 3665
rect -16146 3631 -16130 3665
rect -16196 3597 -16130 3631
rect -16196 3563 -16180 3597
rect -16146 3563 -16130 3597
rect -16196 3529 -16130 3563
rect -16196 3495 -16180 3529
rect -16146 3495 -16130 3529
rect -16196 3454 -16130 3495
rect -16100 4413 -16034 4454
rect -16100 4379 -16084 4413
rect -16050 4379 -16034 4413
rect -16100 4345 -16034 4379
rect -16100 4311 -16084 4345
rect -16050 4311 -16034 4345
rect -16100 4277 -16034 4311
rect -16100 4243 -16084 4277
rect -16050 4243 -16034 4277
rect -16100 4209 -16034 4243
rect -16100 4175 -16084 4209
rect -16050 4175 -16034 4209
rect -16100 4141 -16034 4175
rect -16100 4107 -16084 4141
rect -16050 4107 -16034 4141
rect -16100 4073 -16034 4107
rect -16100 4039 -16084 4073
rect -16050 4039 -16034 4073
rect -16100 4005 -16034 4039
rect -16100 3971 -16084 4005
rect -16050 3971 -16034 4005
rect -16100 3937 -16034 3971
rect -16100 3903 -16084 3937
rect -16050 3903 -16034 3937
rect -16100 3869 -16034 3903
rect -16100 3835 -16084 3869
rect -16050 3835 -16034 3869
rect -16100 3801 -16034 3835
rect -16100 3767 -16084 3801
rect -16050 3767 -16034 3801
rect -16100 3733 -16034 3767
rect -16100 3699 -16084 3733
rect -16050 3699 -16034 3733
rect -16100 3665 -16034 3699
rect -16100 3631 -16084 3665
rect -16050 3631 -16034 3665
rect -16100 3597 -16034 3631
rect -16100 3563 -16084 3597
rect -16050 3563 -16034 3597
rect -16100 3529 -16034 3563
rect -16100 3495 -16084 3529
rect -16050 3495 -16034 3529
rect -16100 3454 -16034 3495
rect -16004 4413 -15938 4454
rect -16004 4379 -15988 4413
rect -15954 4379 -15938 4413
rect -16004 4345 -15938 4379
rect -16004 4311 -15988 4345
rect -15954 4311 -15938 4345
rect -16004 4277 -15938 4311
rect -16004 4243 -15988 4277
rect -15954 4243 -15938 4277
rect -16004 4209 -15938 4243
rect -16004 4175 -15988 4209
rect -15954 4175 -15938 4209
rect -16004 4141 -15938 4175
rect -16004 4107 -15988 4141
rect -15954 4107 -15938 4141
rect -16004 4073 -15938 4107
rect -16004 4039 -15988 4073
rect -15954 4039 -15938 4073
rect -16004 4005 -15938 4039
rect -16004 3971 -15988 4005
rect -15954 3971 -15938 4005
rect -16004 3937 -15938 3971
rect -16004 3903 -15988 3937
rect -15954 3903 -15938 3937
rect -16004 3869 -15938 3903
rect -16004 3835 -15988 3869
rect -15954 3835 -15938 3869
rect -16004 3801 -15938 3835
rect -16004 3767 -15988 3801
rect -15954 3767 -15938 3801
rect -16004 3733 -15938 3767
rect -16004 3699 -15988 3733
rect -15954 3699 -15938 3733
rect -16004 3665 -15938 3699
rect -16004 3631 -15988 3665
rect -15954 3631 -15938 3665
rect -16004 3597 -15938 3631
rect -16004 3563 -15988 3597
rect -15954 3563 -15938 3597
rect -16004 3529 -15938 3563
rect -16004 3495 -15988 3529
rect -15954 3495 -15938 3529
rect -16004 3454 -15938 3495
rect -15908 4413 -15842 4454
rect -15908 4379 -15892 4413
rect -15858 4379 -15842 4413
rect -15908 4345 -15842 4379
rect -15908 4311 -15892 4345
rect -15858 4311 -15842 4345
rect -15908 4277 -15842 4311
rect -15908 4243 -15892 4277
rect -15858 4243 -15842 4277
rect -15908 4209 -15842 4243
rect -15908 4175 -15892 4209
rect -15858 4175 -15842 4209
rect -15908 4141 -15842 4175
rect -15908 4107 -15892 4141
rect -15858 4107 -15842 4141
rect -15908 4073 -15842 4107
rect -15908 4039 -15892 4073
rect -15858 4039 -15842 4073
rect -15908 4005 -15842 4039
rect -15908 3971 -15892 4005
rect -15858 3971 -15842 4005
rect -15908 3937 -15842 3971
rect -15908 3903 -15892 3937
rect -15858 3903 -15842 3937
rect -15908 3869 -15842 3903
rect -15908 3835 -15892 3869
rect -15858 3835 -15842 3869
rect -15908 3801 -15842 3835
rect -15908 3767 -15892 3801
rect -15858 3767 -15842 3801
rect -15908 3733 -15842 3767
rect -15908 3699 -15892 3733
rect -15858 3699 -15842 3733
rect -15908 3665 -15842 3699
rect -15908 3631 -15892 3665
rect -15858 3631 -15842 3665
rect -15908 3597 -15842 3631
rect -15908 3563 -15892 3597
rect -15858 3563 -15842 3597
rect -15908 3529 -15842 3563
rect -15908 3495 -15892 3529
rect -15858 3495 -15842 3529
rect -15908 3454 -15842 3495
rect -15812 4413 -15746 4454
rect -15812 4379 -15796 4413
rect -15762 4379 -15746 4413
rect -15812 4345 -15746 4379
rect -15812 4311 -15796 4345
rect -15762 4311 -15746 4345
rect -15812 4277 -15746 4311
rect -15812 4243 -15796 4277
rect -15762 4243 -15746 4277
rect -15812 4209 -15746 4243
rect -15812 4175 -15796 4209
rect -15762 4175 -15746 4209
rect -15812 4141 -15746 4175
rect -15812 4107 -15796 4141
rect -15762 4107 -15746 4141
rect -15812 4073 -15746 4107
rect -15812 4039 -15796 4073
rect -15762 4039 -15746 4073
rect -15812 4005 -15746 4039
rect -15812 3971 -15796 4005
rect -15762 3971 -15746 4005
rect -15812 3937 -15746 3971
rect -15812 3903 -15796 3937
rect -15762 3903 -15746 3937
rect -15812 3869 -15746 3903
rect -15812 3835 -15796 3869
rect -15762 3835 -15746 3869
rect -15812 3801 -15746 3835
rect -15812 3767 -15796 3801
rect -15762 3767 -15746 3801
rect -15812 3733 -15746 3767
rect -15812 3699 -15796 3733
rect -15762 3699 -15746 3733
rect -15812 3665 -15746 3699
rect -15812 3631 -15796 3665
rect -15762 3631 -15746 3665
rect -15812 3597 -15746 3631
rect -15812 3563 -15796 3597
rect -15762 3563 -15746 3597
rect -15812 3529 -15746 3563
rect -15812 3495 -15796 3529
rect -15762 3495 -15746 3529
rect -15812 3454 -15746 3495
rect -15716 4413 -15650 4454
rect -15716 4379 -15700 4413
rect -15666 4379 -15650 4413
rect -15716 4345 -15650 4379
rect -15716 4311 -15700 4345
rect -15666 4311 -15650 4345
rect -15716 4277 -15650 4311
rect -15716 4243 -15700 4277
rect -15666 4243 -15650 4277
rect -15716 4209 -15650 4243
rect -15716 4175 -15700 4209
rect -15666 4175 -15650 4209
rect -15716 4141 -15650 4175
rect -15716 4107 -15700 4141
rect -15666 4107 -15650 4141
rect -15716 4073 -15650 4107
rect -15716 4039 -15700 4073
rect -15666 4039 -15650 4073
rect -15716 4005 -15650 4039
rect -15716 3971 -15700 4005
rect -15666 3971 -15650 4005
rect -15716 3937 -15650 3971
rect -15716 3903 -15700 3937
rect -15666 3903 -15650 3937
rect -15716 3869 -15650 3903
rect -15716 3835 -15700 3869
rect -15666 3835 -15650 3869
rect -15716 3801 -15650 3835
rect -15716 3767 -15700 3801
rect -15666 3767 -15650 3801
rect -15716 3733 -15650 3767
rect -15716 3699 -15700 3733
rect -15666 3699 -15650 3733
rect -15716 3665 -15650 3699
rect -15716 3631 -15700 3665
rect -15666 3631 -15650 3665
rect -15716 3597 -15650 3631
rect -15716 3563 -15700 3597
rect -15666 3563 -15650 3597
rect -15716 3529 -15650 3563
rect -15716 3495 -15700 3529
rect -15666 3495 -15650 3529
rect -15716 3454 -15650 3495
rect -15620 4413 -15554 4454
rect -15620 4379 -15604 4413
rect -15570 4379 -15554 4413
rect -15620 4345 -15554 4379
rect -15620 4311 -15604 4345
rect -15570 4311 -15554 4345
rect -15620 4277 -15554 4311
rect -15620 4243 -15604 4277
rect -15570 4243 -15554 4277
rect -15620 4209 -15554 4243
rect -15620 4175 -15604 4209
rect -15570 4175 -15554 4209
rect -15620 4141 -15554 4175
rect -15620 4107 -15604 4141
rect -15570 4107 -15554 4141
rect -15620 4073 -15554 4107
rect -15620 4039 -15604 4073
rect -15570 4039 -15554 4073
rect -15620 4005 -15554 4039
rect -15620 3971 -15604 4005
rect -15570 3971 -15554 4005
rect -15620 3937 -15554 3971
rect -15620 3903 -15604 3937
rect -15570 3903 -15554 3937
rect -15620 3869 -15554 3903
rect -15620 3835 -15604 3869
rect -15570 3835 -15554 3869
rect -15620 3801 -15554 3835
rect -15620 3767 -15604 3801
rect -15570 3767 -15554 3801
rect -15620 3733 -15554 3767
rect -15620 3699 -15604 3733
rect -15570 3699 -15554 3733
rect -15620 3665 -15554 3699
rect -15620 3631 -15604 3665
rect -15570 3631 -15554 3665
rect -15620 3597 -15554 3631
rect -15620 3563 -15604 3597
rect -15570 3563 -15554 3597
rect -15620 3529 -15554 3563
rect -15620 3495 -15604 3529
rect -15570 3495 -15554 3529
rect -15620 3454 -15554 3495
rect -15524 4413 -15458 4454
rect -15524 4379 -15508 4413
rect -15474 4379 -15458 4413
rect -15524 4345 -15458 4379
rect -15524 4311 -15508 4345
rect -15474 4311 -15458 4345
rect -15524 4277 -15458 4311
rect -15524 4243 -15508 4277
rect -15474 4243 -15458 4277
rect -15524 4209 -15458 4243
rect -15524 4175 -15508 4209
rect -15474 4175 -15458 4209
rect -15524 4141 -15458 4175
rect -15524 4107 -15508 4141
rect -15474 4107 -15458 4141
rect -15524 4073 -15458 4107
rect -15524 4039 -15508 4073
rect -15474 4039 -15458 4073
rect -15524 4005 -15458 4039
rect -15524 3971 -15508 4005
rect -15474 3971 -15458 4005
rect -15524 3937 -15458 3971
rect -15524 3903 -15508 3937
rect -15474 3903 -15458 3937
rect -15524 3869 -15458 3903
rect -15524 3835 -15508 3869
rect -15474 3835 -15458 3869
rect -15524 3801 -15458 3835
rect -15524 3767 -15508 3801
rect -15474 3767 -15458 3801
rect -15524 3733 -15458 3767
rect -15524 3699 -15508 3733
rect -15474 3699 -15458 3733
rect -15524 3665 -15458 3699
rect -15524 3631 -15508 3665
rect -15474 3631 -15458 3665
rect -15524 3597 -15458 3631
rect -15524 3563 -15508 3597
rect -15474 3563 -15458 3597
rect -15524 3529 -15458 3563
rect -15524 3495 -15508 3529
rect -15474 3495 -15458 3529
rect -15524 3454 -15458 3495
rect -15428 4413 -15362 4454
rect -15428 4379 -15412 4413
rect -15378 4379 -15362 4413
rect -15428 4345 -15362 4379
rect -15428 4311 -15412 4345
rect -15378 4311 -15362 4345
rect -15428 4277 -15362 4311
rect -15428 4243 -15412 4277
rect -15378 4243 -15362 4277
rect -15428 4209 -15362 4243
rect -15428 4175 -15412 4209
rect -15378 4175 -15362 4209
rect -15428 4141 -15362 4175
rect -15428 4107 -15412 4141
rect -15378 4107 -15362 4141
rect -15428 4073 -15362 4107
rect -15428 4039 -15412 4073
rect -15378 4039 -15362 4073
rect -15428 4005 -15362 4039
rect -15428 3971 -15412 4005
rect -15378 3971 -15362 4005
rect -15428 3937 -15362 3971
rect -15428 3903 -15412 3937
rect -15378 3903 -15362 3937
rect -15428 3869 -15362 3903
rect -15428 3835 -15412 3869
rect -15378 3835 -15362 3869
rect -15428 3801 -15362 3835
rect -15428 3767 -15412 3801
rect -15378 3767 -15362 3801
rect -15428 3733 -15362 3767
rect -15428 3699 -15412 3733
rect -15378 3699 -15362 3733
rect -15428 3665 -15362 3699
rect -15428 3631 -15412 3665
rect -15378 3631 -15362 3665
rect -15428 3597 -15362 3631
rect -15428 3563 -15412 3597
rect -15378 3563 -15362 3597
rect -15428 3529 -15362 3563
rect -15428 3495 -15412 3529
rect -15378 3495 -15362 3529
rect -15428 3454 -15362 3495
rect -15332 4413 -15266 4454
rect -15332 4379 -15316 4413
rect -15282 4379 -15266 4413
rect -15332 4345 -15266 4379
rect -15332 4311 -15316 4345
rect -15282 4311 -15266 4345
rect -15332 4277 -15266 4311
rect -15332 4243 -15316 4277
rect -15282 4243 -15266 4277
rect -15332 4209 -15266 4243
rect -15332 4175 -15316 4209
rect -15282 4175 -15266 4209
rect -15332 4141 -15266 4175
rect -15332 4107 -15316 4141
rect -15282 4107 -15266 4141
rect -15332 4073 -15266 4107
rect -15332 4039 -15316 4073
rect -15282 4039 -15266 4073
rect -15332 4005 -15266 4039
rect -15332 3971 -15316 4005
rect -15282 3971 -15266 4005
rect -15332 3937 -15266 3971
rect -15332 3903 -15316 3937
rect -15282 3903 -15266 3937
rect -15332 3869 -15266 3903
rect -15332 3835 -15316 3869
rect -15282 3835 -15266 3869
rect -15332 3801 -15266 3835
rect -15332 3767 -15316 3801
rect -15282 3767 -15266 3801
rect -15332 3733 -15266 3767
rect -15332 3699 -15316 3733
rect -15282 3699 -15266 3733
rect -15332 3665 -15266 3699
rect -15332 3631 -15316 3665
rect -15282 3631 -15266 3665
rect -15332 3597 -15266 3631
rect -15332 3563 -15316 3597
rect -15282 3563 -15266 3597
rect -15332 3529 -15266 3563
rect -15332 3495 -15316 3529
rect -15282 3495 -15266 3529
rect -15332 3454 -15266 3495
rect -15236 4413 -15170 4454
rect -15236 4379 -15220 4413
rect -15186 4379 -15170 4413
rect -15236 4345 -15170 4379
rect -15236 4311 -15220 4345
rect -15186 4311 -15170 4345
rect -15236 4277 -15170 4311
rect -15236 4243 -15220 4277
rect -15186 4243 -15170 4277
rect -15236 4209 -15170 4243
rect -15236 4175 -15220 4209
rect -15186 4175 -15170 4209
rect -15236 4141 -15170 4175
rect -15236 4107 -15220 4141
rect -15186 4107 -15170 4141
rect -15236 4073 -15170 4107
rect -15236 4039 -15220 4073
rect -15186 4039 -15170 4073
rect -15236 4005 -15170 4039
rect -15236 3971 -15220 4005
rect -15186 3971 -15170 4005
rect -15236 3937 -15170 3971
rect -15236 3903 -15220 3937
rect -15186 3903 -15170 3937
rect -15236 3869 -15170 3903
rect -15236 3835 -15220 3869
rect -15186 3835 -15170 3869
rect -15236 3801 -15170 3835
rect -15236 3767 -15220 3801
rect -15186 3767 -15170 3801
rect -15236 3733 -15170 3767
rect -15236 3699 -15220 3733
rect -15186 3699 -15170 3733
rect -15236 3665 -15170 3699
rect -15236 3631 -15220 3665
rect -15186 3631 -15170 3665
rect -15236 3597 -15170 3631
rect -15236 3563 -15220 3597
rect -15186 3563 -15170 3597
rect -15236 3529 -15170 3563
rect -15236 3495 -15220 3529
rect -15186 3495 -15170 3529
rect -15236 3454 -15170 3495
rect -15140 4413 -15074 4454
rect -15140 4379 -15124 4413
rect -15090 4379 -15074 4413
rect -15140 4345 -15074 4379
rect -15140 4311 -15124 4345
rect -15090 4311 -15074 4345
rect -15140 4277 -15074 4311
rect -15140 4243 -15124 4277
rect -15090 4243 -15074 4277
rect -15140 4209 -15074 4243
rect -15140 4175 -15124 4209
rect -15090 4175 -15074 4209
rect -15140 4141 -15074 4175
rect -15140 4107 -15124 4141
rect -15090 4107 -15074 4141
rect -15140 4073 -15074 4107
rect -15140 4039 -15124 4073
rect -15090 4039 -15074 4073
rect -15140 4005 -15074 4039
rect -15140 3971 -15124 4005
rect -15090 3971 -15074 4005
rect -15140 3937 -15074 3971
rect -15140 3903 -15124 3937
rect -15090 3903 -15074 3937
rect -15140 3869 -15074 3903
rect -15140 3835 -15124 3869
rect -15090 3835 -15074 3869
rect -15140 3801 -15074 3835
rect -15140 3767 -15124 3801
rect -15090 3767 -15074 3801
rect -15140 3733 -15074 3767
rect -15140 3699 -15124 3733
rect -15090 3699 -15074 3733
rect -15140 3665 -15074 3699
rect -15140 3631 -15124 3665
rect -15090 3631 -15074 3665
rect -15140 3597 -15074 3631
rect -15140 3563 -15124 3597
rect -15090 3563 -15074 3597
rect -15140 3529 -15074 3563
rect -15140 3495 -15124 3529
rect -15090 3495 -15074 3529
rect -15140 3454 -15074 3495
rect -15044 4413 -14978 4454
rect -15044 4379 -15028 4413
rect -14994 4379 -14978 4413
rect -15044 4345 -14978 4379
rect -15044 4311 -15028 4345
rect -14994 4311 -14978 4345
rect -15044 4277 -14978 4311
rect -15044 4243 -15028 4277
rect -14994 4243 -14978 4277
rect -15044 4209 -14978 4243
rect -15044 4175 -15028 4209
rect -14994 4175 -14978 4209
rect -15044 4141 -14978 4175
rect -15044 4107 -15028 4141
rect -14994 4107 -14978 4141
rect -15044 4073 -14978 4107
rect -15044 4039 -15028 4073
rect -14994 4039 -14978 4073
rect -15044 4005 -14978 4039
rect -15044 3971 -15028 4005
rect -14994 3971 -14978 4005
rect -15044 3937 -14978 3971
rect -15044 3903 -15028 3937
rect -14994 3903 -14978 3937
rect -15044 3869 -14978 3903
rect -15044 3835 -15028 3869
rect -14994 3835 -14978 3869
rect -15044 3801 -14978 3835
rect -15044 3767 -15028 3801
rect -14994 3767 -14978 3801
rect -15044 3733 -14978 3767
rect -15044 3699 -15028 3733
rect -14994 3699 -14978 3733
rect -15044 3665 -14978 3699
rect -15044 3631 -15028 3665
rect -14994 3631 -14978 3665
rect -15044 3597 -14978 3631
rect -15044 3563 -15028 3597
rect -14994 3563 -14978 3597
rect -15044 3529 -14978 3563
rect -15044 3495 -15028 3529
rect -14994 3495 -14978 3529
rect -15044 3454 -14978 3495
rect -14948 4413 -14882 4454
rect -14948 4379 -14932 4413
rect -14898 4379 -14882 4413
rect -14948 4345 -14882 4379
rect -14948 4311 -14932 4345
rect -14898 4311 -14882 4345
rect -14948 4277 -14882 4311
rect -14948 4243 -14932 4277
rect -14898 4243 -14882 4277
rect -14948 4209 -14882 4243
rect -14948 4175 -14932 4209
rect -14898 4175 -14882 4209
rect -14948 4141 -14882 4175
rect -14948 4107 -14932 4141
rect -14898 4107 -14882 4141
rect -14948 4073 -14882 4107
rect -14948 4039 -14932 4073
rect -14898 4039 -14882 4073
rect -14948 4005 -14882 4039
rect -14948 3971 -14932 4005
rect -14898 3971 -14882 4005
rect -14948 3937 -14882 3971
rect -14948 3903 -14932 3937
rect -14898 3903 -14882 3937
rect -14948 3869 -14882 3903
rect -14948 3835 -14932 3869
rect -14898 3835 -14882 3869
rect -14948 3801 -14882 3835
rect -14948 3767 -14932 3801
rect -14898 3767 -14882 3801
rect -14948 3733 -14882 3767
rect -14948 3699 -14932 3733
rect -14898 3699 -14882 3733
rect -14948 3665 -14882 3699
rect -14948 3631 -14932 3665
rect -14898 3631 -14882 3665
rect -14948 3597 -14882 3631
rect -14948 3563 -14932 3597
rect -14898 3563 -14882 3597
rect -14948 3529 -14882 3563
rect -14948 3495 -14932 3529
rect -14898 3495 -14882 3529
rect -14948 3454 -14882 3495
rect -14852 4413 -14790 4454
rect -14852 4379 -14836 4413
rect -14802 4379 -14790 4413
rect -14852 4345 -14790 4379
rect -14852 4311 -14836 4345
rect -14802 4311 -14790 4345
rect -14852 4277 -14790 4311
rect -14852 4243 -14836 4277
rect -14802 4243 -14790 4277
rect -14852 4209 -14790 4243
rect -14852 4175 -14836 4209
rect -14802 4175 -14790 4209
rect -14852 4141 -14790 4175
rect -14852 4107 -14836 4141
rect -14802 4107 -14790 4141
rect -14852 4073 -14790 4107
rect -14852 4039 -14836 4073
rect -14802 4039 -14790 4073
rect -14852 4005 -14790 4039
rect -14852 3971 -14836 4005
rect -14802 3971 -14790 4005
rect -14852 3937 -14790 3971
rect -14852 3903 -14836 3937
rect -14802 3903 -14790 3937
rect -14852 3869 -14790 3903
rect -14852 3835 -14836 3869
rect -14802 3835 -14790 3869
rect -14852 3801 -14790 3835
rect -14852 3767 -14836 3801
rect -14802 3767 -14790 3801
rect -14852 3733 -14790 3767
rect -14852 3699 -14836 3733
rect -14802 3699 -14790 3733
rect -14852 3665 -14790 3699
rect -14852 3631 -14836 3665
rect -14802 3631 -14790 3665
rect -14852 3597 -14790 3631
rect -14852 3563 -14836 3597
rect -14802 3563 -14790 3597
rect -14852 3529 -14790 3563
rect -14852 3495 -14836 3529
rect -14802 3495 -14790 3529
rect -14852 3454 -14790 3495
rect -14624 4419 -14562 4460
rect -14624 4385 -14612 4419
rect -14578 4385 -14562 4419
rect -14624 4351 -14562 4385
rect -14624 4317 -14612 4351
rect -14578 4317 -14562 4351
rect -14624 4283 -14562 4317
rect -14624 4249 -14612 4283
rect -14578 4249 -14562 4283
rect -14624 4215 -14562 4249
rect -14624 4181 -14612 4215
rect -14578 4181 -14562 4215
rect -14624 4147 -14562 4181
rect -14624 4113 -14612 4147
rect -14578 4113 -14562 4147
rect -14624 4079 -14562 4113
rect -14624 4045 -14612 4079
rect -14578 4045 -14562 4079
rect -14624 4011 -14562 4045
rect -14624 3977 -14612 4011
rect -14578 3977 -14562 4011
rect -14624 3943 -14562 3977
rect -14624 3909 -14612 3943
rect -14578 3909 -14562 3943
rect -14624 3875 -14562 3909
rect -14624 3841 -14612 3875
rect -14578 3841 -14562 3875
rect -14624 3807 -14562 3841
rect -14624 3773 -14612 3807
rect -14578 3773 -14562 3807
rect -14624 3739 -14562 3773
rect -14624 3705 -14612 3739
rect -14578 3705 -14562 3739
rect -14624 3671 -14562 3705
rect -14624 3637 -14612 3671
rect -14578 3637 -14562 3671
rect -14624 3603 -14562 3637
rect -14624 3569 -14612 3603
rect -14578 3569 -14562 3603
rect -14624 3535 -14562 3569
rect -14624 3501 -14612 3535
rect -14578 3501 -14562 3535
rect -14624 3460 -14562 3501
rect -14532 4419 -14466 4460
rect -14532 4385 -14516 4419
rect -14482 4385 -14466 4419
rect -14532 4351 -14466 4385
rect -14532 4317 -14516 4351
rect -14482 4317 -14466 4351
rect -14532 4283 -14466 4317
rect -14532 4249 -14516 4283
rect -14482 4249 -14466 4283
rect -14532 4215 -14466 4249
rect -14532 4181 -14516 4215
rect -14482 4181 -14466 4215
rect -14532 4147 -14466 4181
rect -14532 4113 -14516 4147
rect -14482 4113 -14466 4147
rect -14532 4079 -14466 4113
rect -14532 4045 -14516 4079
rect -14482 4045 -14466 4079
rect -14532 4011 -14466 4045
rect -14532 3977 -14516 4011
rect -14482 3977 -14466 4011
rect -14532 3943 -14466 3977
rect -14532 3909 -14516 3943
rect -14482 3909 -14466 3943
rect -14532 3875 -14466 3909
rect -14532 3841 -14516 3875
rect -14482 3841 -14466 3875
rect -14532 3807 -14466 3841
rect -14532 3773 -14516 3807
rect -14482 3773 -14466 3807
rect -14532 3739 -14466 3773
rect -14532 3705 -14516 3739
rect -14482 3705 -14466 3739
rect -14532 3671 -14466 3705
rect -14532 3637 -14516 3671
rect -14482 3637 -14466 3671
rect -14532 3603 -14466 3637
rect -14532 3569 -14516 3603
rect -14482 3569 -14466 3603
rect -14532 3535 -14466 3569
rect -14532 3501 -14516 3535
rect -14482 3501 -14466 3535
rect -14532 3460 -14466 3501
rect -14436 4419 -14370 4460
rect -14436 4385 -14420 4419
rect -14386 4385 -14370 4419
rect -14436 4351 -14370 4385
rect -14436 4317 -14420 4351
rect -14386 4317 -14370 4351
rect -14436 4283 -14370 4317
rect -14436 4249 -14420 4283
rect -14386 4249 -14370 4283
rect -14436 4215 -14370 4249
rect -14436 4181 -14420 4215
rect -14386 4181 -14370 4215
rect -14436 4147 -14370 4181
rect -14436 4113 -14420 4147
rect -14386 4113 -14370 4147
rect -14436 4079 -14370 4113
rect -14436 4045 -14420 4079
rect -14386 4045 -14370 4079
rect -14436 4011 -14370 4045
rect -14436 3977 -14420 4011
rect -14386 3977 -14370 4011
rect -14436 3943 -14370 3977
rect -14436 3909 -14420 3943
rect -14386 3909 -14370 3943
rect -14436 3875 -14370 3909
rect -14436 3841 -14420 3875
rect -14386 3841 -14370 3875
rect -14436 3807 -14370 3841
rect -14436 3773 -14420 3807
rect -14386 3773 -14370 3807
rect -14436 3739 -14370 3773
rect -14436 3705 -14420 3739
rect -14386 3705 -14370 3739
rect -14436 3671 -14370 3705
rect -14436 3637 -14420 3671
rect -14386 3637 -14370 3671
rect -14436 3603 -14370 3637
rect -14436 3569 -14420 3603
rect -14386 3569 -14370 3603
rect -14436 3535 -14370 3569
rect -14436 3501 -14420 3535
rect -14386 3501 -14370 3535
rect -14436 3460 -14370 3501
rect -14340 4419 -14274 4460
rect -14340 4385 -14324 4419
rect -14290 4385 -14274 4419
rect -14340 4351 -14274 4385
rect -14340 4317 -14324 4351
rect -14290 4317 -14274 4351
rect -14340 4283 -14274 4317
rect -14340 4249 -14324 4283
rect -14290 4249 -14274 4283
rect -14340 4215 -14274 4249
rect -14340 4181 -14324 4215
rect -14290 4181 -14274 4215
rect -14340 4147 -14274 4181
rect -14340 4113 -14324 4147
rect -14290 4113 -14274 4147
rect -14340 4079 -14274 4113
rect -14340 4045 -14324 4079
rect -14290 4045 -14274 4079
rect -14340 4011 -14274 4045
rect -14340 3977 -14324 4011
rect -14290 3977 -14274 4011
rect -14340 3943 -14274 3977
rect -14340 3909 -14324 3943
rect -14290 3909 -14274 3943
rect -14340 3875 -14274 3909
rect -14340 3841 -14324 3875
rect -14290 3841 -14274 3875
rect -14340 3807 -14274 3841
rect -14340 3773 -14324 3807
rect -14290 3773 -14274 3807
rect -14340 3739 -14274 3773
rect -14340 3705 -14324 3739
rect -14290 3705 -14274 3739
rect -14340 3671 -14274 3705
rect -14340 3637 -14324 3671
rect -14290 3637 -14274 3671
rect -14340 3603 -14274 3637
rect -14340 3569 -14324 3603
rect -14290 3569 -14274 3603
rect -14340 3535 -14274 3569
rect -14340 3501 -14324 3535
rect -14290 3501 -14274 3535
rect -14340 3460 -14274 3501
rect -14244 4419 -14178 4460
rect -14244 4385 -14228 4419
rect -14194 4385 -14178 4419
rect -14244 4351 -14178 4385
rect -14244 4317 -14228 4351
rect -14194 4317 -14178 4351
rect -14244 4283 -14178 4317
rect -14244 4249 -14228 4283
rect -14194 4249 -14178 4283
rect -14244 4215 -14178 4249
rect -14244 4181 -14228 4215
rect -14194 4181 -14178 4215
rect -14244 4147 -14178 4181
rect -14244 4113 -14228 4147
rect -14194 4113 -14178 4147
rect -14244 4079 -14178 4113
rect -14244 4045 -14228 4079
rect -14194 4045 -14178 4079
rect -14244 4011 -14178 4045
rect -14244 3977 -14228 4011
rect -14194 3977 -14178 4011
rect -14244 3943 -14178 3977
rect -14244 3909 -14228 3943
rect -14194 3909 -14178 3943
rect -14244 3875 -14178 3909
rect -14244 3841 -14228 3875
rect -14194 3841 -14178 3875
rect -14244 3807 -14178 3841
rect -14244 3773 -14228 3807
rect -14194 3773 -14178 3807
rect -14244 3739 -14178 3773
rect -14244 3705 -14228 3739
rect -14194 3705 -14178 3739
rect -14244 3671 -14178 3705
rect -14244 3637 -14228 3671
rect -14194 3637 -14178 3671
rect -14244 3603 -14178 3637
rect -14244 3569 -14228 3603
rect -14194 3569 -14178 3603
rect -14244 3535 -14178 3569
rect -14244 3501 -14228 3535
rect -14194 3501 -14178 3535
rect -14244 3460 -14178 3501
rect -14148 4419 -14082 4460
rect -14148 4385 -14132 4419
rect -14098 4385 -14082 4419
rect -14148 4351 -14082 4385
rect -14148 4317 -14132 4351
rect -14098 4317 -14082 4351
rect -14148 4283 -14082 4317
rect -14148 4249 -14132 4283
rect -14098 4249 -14082 4283
rect -14148 4215 -14082 4249
rect -14148 4181 -14132 4215
rect -14098 4181 -14082 4215
rect -14148 4147 -14082 4181
rect -14148 4113 -14132 4147
rect -14098 4113 -14082 4147
rect -14148 4079 -14082 4113
rect -14148 4045 -14132 4079
rect -14098 4045 -14082 4079
rect -14148 4011 -14082 4045
rect -14148 3977 -14132 4011
rect -14098 3977 -14082 4011
rect -14148 3943 -14082 3977
rect -14148 3909 -14132 3943
rect -14098 3909 -14082 3943
rect -14148 3875 -14082 3909
rect -14148 3841 -14132 3875
rect -14098 3841 -14082 3875
rect -14148 3807 -14082 3841
rect -14148 3773 -14132 3807
rect -14098 3773 -14082 3807
rect -14148 3739 -14082 3773
rect -14148 3705 -14132 3739
rect -14098 3705 -14082 3739
rect -14148 3671 -14082 3705
rect -14148 3637 -14132 3671
rect -14098 3637 -14082 3671
rect -14148 3603 -14082 3637
rect -14148 3569 -14132 3603
rect -14098 3569 -14082 3603
rect -14148 3535 -14082 3569
rect -14148 3501 -14132 3535
rect -14098 3501 -14082 3535
rect -14148 3460 -14082 3501
rect -14052 4419 -13986 4460
rect -14052 4385 -14036 4419
rect -14002 4385 -13986 4419
rect -14052 4351 -13986 4385
rect -14052 4317 -14036 4351
rect -14002 4317 -13986 4351
rect -14052 4283 -13986 4317
rect -14052 4249 -14036 4283
rect -14002 4249 -13986 4283
rect -14052 4215 -13986 4249
rect -14052 4181 -14036 4215
rect -14002 4181 -13986 4215
rect -14052 4147 -13986 4181
rect -14052 4113 -14036 4147
rect -14002 4113 -13986 4147
rect -14052 4079 -13986 4113
rect -14052 4045 -14036 4079
rect -14002 4045 -13986 4079
rect -14052 4011 -13986 4045
rect -14052 3977 -14036 4011
rect -14002 3977 -13986 4011
rect -14052 3943 -13986 3977
rect -14052 3909 -14036 3943
rect -14002 3909 -13986 3943
rect -14052 3875 -13986 3909
rect -14052 3841 -14036 3875
rect -14002 3841 -13986 3875
rect -14052 3807 -13986 3841
rect -14052 3773 -14036 3807
rect -14002 3773 -13986 3807
rect -14052 3739 -13986 3773
rect -14052 3705 -14036 3739
rect -14002 3705 -13986 3739
rect -14052 3671 -13986 3705
rect -14052 3637 -14036 3671
rect -14002 3637 -13986 3671
rect -14052 3603 -13986 3637
rect -14052 3569 -14036 3603
rect -14002 3569 -13986 3603
rect -14052 3535 -13986 3569
rect -14052 3501 -14036 3535
rect -14002 3501 -13986 3535
rect -14052 3460 -13986 3501
rect -13956 4419 -13890 4460
rect -13956 4385 -13940 4419
rect -13906 4385 -13890 4419
rect -13956 4351 -13890 4385
rect -13956 4317 -13940 4351
rect -13906 4317 -13890 4351
rect -13956 4283 -13890 4317
rect -13956 4249 -13940 4283
rect -13906 4249 -13890 4283
rect -13956 4215 -13890 4249
rect -13956 4181 -13940 4215
rect -13906 4181 -13890 4215
rect -13956 4147 -13890 4181
rect -13956 4113 -13940 4147
rect -13906 4113 -13890 4147
rect -13956 4079 -13890 4113
rect -13956 4045 -13940 4079
rect -13906 4045 -13890 4079
rect -13956 4011 -13890 4045
rect -13956 3977 -13940 4011
rect -13906 3977 -13890 4011
rect -13956 3943 -13890 3977
rect -13956 3909 -13940 3943
rect -13906 3909 -13890 3943
rect -13956 3875 -13890 3909
rect -13956 3841 -13940 3875
rect -13906 3841 -13890 3875
rect -13956 3807 -13890 3841
rect -13956 3773 -13940 3807
rect -13906 3773 -13890 3807
rect -13956 3739 -13890 3773
rect -13956 3705 -13940 3739
rect -13906 3705 -13890 3739
rect -13956 3671 -13890 3705
rect -13956 3637 -13940 3671
rect -13906 3637 -13890 3671
rect -13956 3603 -13890 3637
rect -13956 3569 -13940 3603
rect -13906 3569 -13890 3603
rect -13956 3535 -13890 3569
rect -13956 3501 -13940 3535
rect -13906 3501 -13890 3535
rect -13956 3460 -13890 3501
rect -13860 4419 -13794 4460
rect -13860 4385 -13844 4419
rect -13810 4385 -13794 4419
rect -13860 4351 -13794 4385
rect -13860 4317 -13844 4351
rect -13810 4317 -13794 4351
rect -13860 4283 -13794 4317
rect -13860 4249 -13844 4283
rect -13810 4249 -13794 4283
rect -13860 4215 -13794 4249
rect -13860 4181 -13844 4215
rect -13810 4181 -13794 4215
rect -13860 4147 -13794 4181
rect -13860 4113 -13844 4147
rect -13810 4113 -13794 4147
rect -13860 4079 -13794 4113
rect -13860 4045 -13844 4079
rect -13810 4045 -13794 4079
rect -13860 4011 -13794 4045
rect -13860 3977 -13844 4011
rect -13810 3977 -13794 4011
rect -13860 3943 -13794 3977
rect -13860 3909 -13844 3943
rect -13810 3909 -13794 3943
rect -13860 3875 -13794 3909
rect -13860 3841 -13844 3875
rect -13810 3841 -13794 3875
rect -13860 3807 -13794 3841
rect -13860 3773 -13844 3807
rect -13810 3773 -13794 3807
rect -13860 3739 -13794 3773
rect -13860 3705 -13844 3739
rect -13810 3705 -13794 3739
rect -13860 3671 -13794 3705
rect -13860 3637 -13844 3671
rect -13810 3637 -13794 3671
rect -13860 3603 -13794 3637
rect -13860 3569 -13844 3603
rect -13810 3569 -13794 3603
rect -13860 3535 -13794 3569
rect -13860 3501 -13844 3535
rect -13810 3501 -13794 3535
rect -13860 3460 -13794 3501
rect -13764 4419 -13698 4460
rect -13764 4385 -13748 4419
rect -13714 4385 -13698 4419
rect -13764 4351 -13698 4385
rect -13764 4317 -13748 4351
rect -13714 4317 -13698 4351
rect -13764 4283 -13698 4317
rect -13764 4249 -13748 4283
rect -13714 4249 -13698 4283
rect -13764 4215 -13698 4249
rect -13764 4181 -13748 4215
rect -13714 4181 -13698 4215
rect -13764 4147 -13698 4181
rect -13764 4113 -13748 4147
rect -13714 4113 -13698 4147
rect -13764 4079 -13698 4113
rect -13764 4045 -13748 4079
rect -13714 4045 -13698 4079
rect -13764 4011 -13698 4045
rect -13764 3977 -13748 4011
rect -13714 3977 -13698 4011
rect -13764 3943 -13698 3977
rect -13764 3909 -13748 3943
rect -13714 3909 -13698 3943
rect -13764 3875 -13698 3909
rect -13764 3841 -13748 3875
rect -13714 3841 -13698 3875
rect -13764 3807 -13698 3841
rect -13764 3773 -13748 3807
rect -13714 3773 -13698 3807
rect -13764 3739 -13698 3773
rect -13764 3705 -13748 3739
rect -13714 3705 -13698 3739
rect -13764 3671 -13698 3705
rect -13764 3637 -13748 3671
rect -13714 3637 -13698 3671
rect -13764 3603 -13698 3637
rect -13764 3569 -13748 3603
rect -13714 3569 -13698 3603
rect -13764 3535 -13698 3569
rect -13764 3501 -13748 3535
rect -13714 3501 -13698 3535
rect -13764 3460 -13698 3501
rect -13668 4419 -13602 4460
rect -13668 4385 -13652 4419
rect -13618 4385 -13602 4419
rect -13668 4351 -13602 4385
rect -13668 4317 -13652 4351
rect -13618 4317 -13602 4351
rect -13668 4283 -13602 4317
rect -13668 4249 -13652 4283
rect -13618 4249 -13602 4283
rect -13668 4215 -13602 4249
rect -13668 4181 -13652 4215
rect -13618 4181 -13602 4215
rect -13668 4147 -13602 4181
rect -13668 4113 -13652 4147
rect -13618 4113 -13602 4147
rect -13668 4079 -13602 4113
rect -13668 4045 -13652 4079
rect -13618 4045 -13602 4079
rect -13668 4011 -13602 4045
rect -13668 3977 -13652 4011
rect -13618 3977 -13602 4011
rect -13668 3943 -13602 3977
rect -13668 3909 -13652 3943
rect -13618 3909 -13602 3943
rect -13668 3875 -13602 3909
rect -13668 3841 -13652 3875
rect -13618 3841 -13602 3875
rect -13668 3807 -13602 3841
rect -13668 3773 -13652 3807
rect -13618 3773 -13602 3807
rect -13668 3739 -13602 3773
rect -13668 3705 -13652 3739
rect -13618 3705 -13602 3739
rect -13668 3671 -13602 3705
rect -13668 3637 -13652 3671
rect -13618 3637 -13602 3671
rect -13668 3603 -13602 3637
rect -13668 3569 -13652 3603
rect -13618 3569 -13602 3603
rect -13668 3535 -13602 3569
rect -13668 3501 -13652 3535
rect -13618 3501 -13602 3535
rect -13668 3460 -13602 3501
rect -13572 4419 -13506 4460
rect -13572 4385 -13556 4419
rect -13522 4385 -13506 4419
rect -13572 4351 -13506 4385
rect -13572 4317 -13556 4351
rect -13522 4317 -13506 4351
rect -13572 4283 -13506 4317
rect -13572 4249 -13556 4283
rect -13522 4249 -13506 4283
rect -13572 4215 -13506 4249
rect -13572 4181 -13556 4215
rect -13522 4181 -13506 4215
rect -13572 4147 -13506 4181
rect -13572 4113 -13556 4147
rect -13522 4113 -13506 4147
rect -13572 4079 -13506 4113
rect -13572 4045 -13556 4079
rect -13522 4045 -13506 4079
rect -13572 4011 -13506 4045
rect -13572 3977 -13556 4011
rect -13522 3977 -13506 4011
rect -13572 3943 -13506 3977
rect -13572 3909 -13556 3943
rect -13522 3909 -13506 3943
rect -13572 3875 -13506 3909
rect -13572 3841 -13556 3875
rect -13522 3841 -13506 3875
rect -13572 3807 -13506 3841
rect -13572 3773 -13556 3807
rect -13522 3773 -13506 3807
rect -13572 3739 -13506 3773
rect -13572 3705 -13556 3739
rect -13522 3705 -13506 3739
rect -13572 3671 -13506 3705
rect -13572 3637 -13556 3671
rect -13522 3637 -13506 3671
rect -13572 3603 -13506 3637
rect -13572 3569 -13556 3603
rect -13522 3569 -13506 3603
rect -13572 3535 -13506 3569
rect -13572 3501 -13556 3535
rect -13522 3501 -13506 3535
rect -13572 3460 -13506 3501
rect -13476 4419 -13410 4460
rect -13476 4385 -13460 4419
rect -13426 4385 -13410 4419
rect -13476 4351 -13410 4385
rect -13476 4317 -13460 4351
rect -13426 4317 -13410 4351
rect -13476 4283 -13410 4317
rect -13476 4249 -13460 4283
rect -13426 4249 -13410 4283
rect -13476 4215 -13410 4249
rect -13476 4181 -13460 4215
rect -13426 4181 -13410 4215
rect -13476 4147 -13410 4181
rect -13476 4113 -13460 4147
rect -13426 4113 -13410 4147
rect -13476 4079 -13410 4113
rect -13476 4045 -13460 4079
rect -13426 4045 -13410 4079
rect -13476 4011 -13410 4045
rect -13476 3977 -13460 4011
rect -13426 3977 -13410 4011
rect -13476 3943 -13410 3977
rect -13476 3909 -13460 3943
rect -13426 3909 -13410 3943
rect -13476 3875 -13410 3909
rect -13476 3841 -13460 3875
rect -13426 3841 -13410 3875
rect -13476 3807 -13410 3841
rect -13476 3773 -13460 3807
rect -13426 3773 -13410 3807
rect -13476 3739 -13410 3773
rect -13476 3705 -13460 3739
rect -13426 3705 -13410 3739
rect -13476 3671 -13410 3705
rect -13476 3637 -13460 3671
rect -13426 3637 -13410 3671
rect -13476 3603 -13410 3637
rect -13476 3569 -13460 3603
rect -13426 3569 -13410 3603
rect -13476 3535 -13410 3569
rect -13476 3501 -13460 3535
rect -13426 3501 -13410 3535
rect -13476 3460 -13410 3501
rect -13380 4419 -13314 4460
rect -13380 4385 -13364 4419
rect -13330 4385 -13314 4419
rect -13380 4351 -13314 4385
rect -13380 4317 -13364 4351
rect -13330 4317 -13314 4351
rect -13380 4283 -13314 4317
rect -13380 4249 -13364 4283
rect -13330 4249 -13314 4283
rect -13380 4215 -13314 4249
rect -13380 4181 -13364 4215
rect -13330 4181 -13314 4215
rect -13380 4147 -13314 4181
rect -13380 4113 -13364 4147
rect -13330 4113 -13314 4147
rect -13380 4079 -13314 4113
rect -13380 4045 -13364 4079
rect -13330 4045 -13314 4079
rect -13380 4011 -13314 4045
rect -13380 3977 -13364 4011
rect -13330 3977 -13314 4011
rect -13380 3943 -13314 3977
rect -13380 3909 -13364 3943
rect -13330 3909 -13314 3943
rect -13380 3875 -13314 3909
rect -13380 3841 -13364 3875
rect -13330 3841 -13314 3875
rect -13380 3807 -13314 3841
rect -13380 3773 -13364 3807
rect -13330 3773 -13314 3807
rect -13380 3739 -13314 3773
rect -13380 3705 -13364 3739
rect -13330 3705 -13314 3739
rect -13380 3671 -13314 3705
rect -13380 3637 -13364 3671
rect -13330 3637 -13314 3671
rect -13380 3603 -13314 3637
rect -13380 3569 -13364 3603
rect -13330 3569 -13314 3603
rect -13380 3535 -13314 3569
rect -13380 3501 -13364 3535
rect -13330 3501 -13314 3535
rect -13380 3460 -13314 3501
rect -13284 4419 -13218 4460
rect -13284 4385 -13268 4419
rect -13234 4385 -13218 4419
rect -13284 4351 -13218 4385
rect -13284 4317 -13268 4351
rect -13234 4317 -13218 4351
rect -13284 4283 -13218 4317
rect -13284 4249 -13268 4283
rect -13234 4249 -13218 4283
rect -13284 4215 -13218 4249
rect -13284 4181 -13268 4215
rect -13234 4181 -13218 4215
rect -13284 4147 -13218 4181
rect -13284 4113 -13268 4147
rect -13234 4113 -13218 4147
rect -13284 4079 -13218 4113
rect -13284 4045 -13268 4079
rect -13234 4045 -13218 4079
rect -13284 4011 -13218 4045
rect -13284 3977 -13268 4011
rect -13234 3977 -13218 4011
rect -13284 3943 -13218 3977
rect -13284 3909 -13268 3943
rect -13234 3909 -13218 3943
rect -13284 3875 -13218 3909
rect -13284 3841 -13268 3875
rect -13234 3841 -13218 3875
rect -13284 3807 -13218 3841
rect -13284 3773 -13268 3807
rect -13234 3773 -13218 3807
rect -13284 3739 -13218 3773
rect -13284 3705 -13268 3739
rect -13234 3705 -13218 3739
rect -13284 3671 -13218 3705
rect -13284 3637 -13268 3671
rect -13234 3637 -13218 3671
rect -13284 3603 -13218 3637
rect -13284 3569 -13268 3603
rect -13234 3569 -13218 3603
rect -13284 3535 -13218 3569
rect -13284 3501 -13268 3535
rect -13234 3501 -13218 3535
rect -13284 3460 -13218 3501
rect -13188 4419 -13126 4460
rect -13188 4385 -13172 4419
rect -13138 4385 -13126 4419
rect -13188 4351 -13126 4385
rect -13188 4317 -13172 4351
rect -13138 4317 -13126 4351
rect -13188 4283 -13126 4317
rect -13188 4249 -13172 4283
rect -13138 4249 -13126 4283
rect -13188 4215 -13126 4249
rect -13188 4181 -13172 4215
rect -13138 4181 -13126 4215
rect -13188 4147 -13126 4181
rect -13188 4113 -13172 4147
rect -13138 4113 -13126 4147
rect -13188 4079 -13126 4113
rect -13188 4045 -13172 4079
rect -13138 4045 -13126 4079
rect -13188 4011 -13126 4045
rect -13188 3977 -13172 4011
rect -13138 3977 -13126 4011
rect -13188 3943 -13126 3977
rect -13188 3909 -13172 3943
rect -13138 3909 -13126 3943
rect -13188 3875 -13126 3909
rect -13188 3841 -13172 3875
rect -13138 3841 -13126 3875
rect -13188 3807 -13126 3841
rect -13188 3773 -13172 3807
rect -13138 3773 -13126 3807
rect -13188 3739 -13126 3773
rect -13188 3705 -13172 3739
rect -13138 3705 -13126 3739
rect -13188 3671 -13126 3705
rect -13188 3637 -13172 3671
rect -13138 3637 -13126 3671
rect -13188 3603 -13126 3637
rect -13188 3569 -13172 3603
rect -13138 3569 -13126 3603
rect -13188 3535 -13126 3569
rect -13188 3501 -13172 3535
rect -13138 3501 -13126 3535
rect -13188 3460 -13126 3501
rect -12940 4425 -12878 4466
rect -12940 4391 -12928 4425
rect -12894 4391 -12878 4425
rect -12940 4357 -12878 4391
rect -12940 4323 -12928 4357
rect -12894 4323 -12878 4357
rect -12940 4289 -12878 4323
rect -12940 4255 -12928 4289
rect -12894 4255 -12878 4289
rect -12940 4221 -12878 4255
rect -12940 4187 -12928 4221
rect -12894 4187 -12878 4221
rect -12940 4153 -12878 4187
rect -12940 4119 -12928 4153
rect -12894 4119 -12878 4153
rect -12940 4085 -12878 4119
rect -12940 4051 -12928 4085
rect -12894 4051 -12878 4085
rect -12940 4017 -12878 4051
rect -12940 3983 -12928 4017
rect -12894 3983 -12878 4017
rect -12940 3949 -12878 3983
rect -12940 3915 -12928 3949
rect -12894 3915 -12878 3949
rect -12940 3881 -12878 3915
rect -12940 3847 -12928 3881
rect -12894 3847 -12878 3881
rect -12940 3813 -12878 3847
rect -12940 3779 -12928 3813
rect -12894 3779 -12878 3813
rect -12940 3745 -12878 3779
rect -12940 3711 -12928 3745
rect -12894 3711 -12878 3745
rect -12940 3677 -12878 3711
rect -12940 3643 -12928 3677
rect -12894 3643 -12878 3677
rect -12940 3609 -12878 3643
rect -12940 3575 -12928 3609
rect -12894 3575 -12878 3609
rect -12940 3541 -12878 3575
rect -12940 3507 -12928 3541
rect -12894 3507 -12878 3541
rect -12940 3466 -12878 3507
rect -12848 4425 -12782 4466
rect -12848 4391 -12832 4425
rect -12798 4391 -12782 4425
rect -12848 4357 -12782 4391
rect -12848 4323 -12832 4357
rect -12798 4323 -12782 4357
rect -12848 4289 -12782 4323
rect -12848 4255 -12832 4289
rect -12798 4255 -12782 4289
rect -12848 4221 -12782 4255
rect -12848 4187 -12832 4221
rect -12798 4187 -12782 4221
rect -12848 4153 -12782 4187
rect -12848 4119 -12832 4153
rect -12798 4119 -12782 4153
rect -12848 4085 -12782 4119
rect -12848 4051 -12832 4085
rect -12798 4051 -12782 4085
rect -12848 4017 -12782 4051
rect -12848 3983 -12832 4017
rect -12798 3983 -12782 4017
rect -12848 3949 -12782 3983
rect -12848 3915 -12832 3949
rect -12798 3915 -12782 3949
rect -12848 3881 -12782 3915
rect -12848 3847 -12832 3881
rect -12798 3847 -12782 3881
rect -12848 3813 -12782 3847
rect -12848 3779 -12832 3813
rect -12798 3779 -12782 3813
rect -12848 3745 -12782 3779
rect -12848 3711 -12832 3745
rect -12798 3711 -12782 3745
rect -12848 3677 -12782 3711
rect -12848 3643 -12832 3677
rect -12798 3643 -12782 3677
rect -12848 3609 -12782 3643
rect -12848 3575 -12832 3609
rect -12798 3575 -12782 3609
rect -12848 3541 -12782 3575
rect -12848 3507 -12832 3541
rect -12798 3507 -12782 3541
rect -12848 3466 -12782 3507
rect -12752 4425 -12686 4466
rect -12752 4391 -12736 4425
rect -12702 4391 -12686 4425
rect -12752 4357 -12686 4391
rect -12752 4323 -12736 4357
rect -12702 4323 -12686 4357
rect -12752 4289 -12686 4323
rect -12752 4255 -12736 4289
rect -12702 4255 -12686 4289
rect -12752 4221 -12686 4255
rect -12752 4187 -12736 4221
rect -12702 4187 -12686 4221
rect -12752 4153 -12686 4187
rect -12752 4119 -12736 4153
rect -12702 4119 -12686 4153
rect -12752 4085 -12686 4119
rect -12752 4051 -12736 4085
rect -12702 4051 -12686 4085
rect -12752 4017 -12686 4051
rect -12752 3983 -12736 4017
rect -12702 3983 -12686 4017
rect -12752 3949 -12686 3983
rect -12752 3915 -12736 3949
rect -12702 3915 -12686 3949
rect -12752 3881 -12686 3915
rect -12752 3847 -12736 3881
rect -12702 3847 -12686 3881
rect -12752 3813 -12686 3847
rect -12752 3779 -12736 3813
rect -12702 3779 -12686 3813
rect -12752 3745 -12686 3779
rect -12752 3711 -12736 3745
rect -12702 3711 -12686 3745
rect -12752 3677 -12686 3711
rect -12752 3643 -12736 3677
rect -12702 3643 -12686 3677
rect -12752 3609 -12686 3643
rect -12752 3575 -12736 3609
rect -12702 3575 -12686 3609
rect -12752 3541 -12686 3575
rect -12752 3507 -12736 3541
rect -12702 3507 -12686 3541
rect -12752 3466 -12686 3507
rect -12656 4425 -12590 4466
rect -12656 4391 -12640 4425
rect -12606 4391 -12590 4425
rect -12656 4357 -12590 4391
rect -12656 4323 -12640 4357
rect -12606 4323 -12590 4357
rect -12656 4289 -12590 4323
rect -12656 4255 -12640 4289
rect -12606 4255 -12590 4289
rect -12656 4221 -12590 4255
rect -12656 4187 -12640 4221
rect -12606 4187 -12590 4221
rect -12656 4153 -12590 4187
rect -12656 4119 -12640 4153
rect -12606 4119 -12590 4153
rect -12656 4085 -12590 4119
rect -12656 4051 -12640 4085
rect -12606 4051 -12590 4085
rect -12656 4017 -12590 4051
rect -12656 3983 -12640 4017
rect -12606 3983 -12590 4017
rect -12656 3949 -12590 3983
rect -12656 3915 -12640 3949
rect -12606 3915 -12590 3949
rect -12656 3881 -12590 3915
rect -12656 3847 -12640 3881
rect -12606 3847 -12590 3881
rect -12656 3813 -12590 3847
rect -12656 3779 -12640 3813
rect -12606 3779 -12590 3813
rect -12656 3745 -12590 3779
rect -12656 3711 -12640 3745
rect -12606 3711 -12590 3745
rect -12656 3677 -12590 3711
rect -12656 3643 -12640 3677
rect -12606 3643 -12590 3677
rect -12656 3609 -12590 3643
rect -12656 3575 -12640 3609
rect -12606 3575 -12590 3609
rect -12656 3541 -12590 3575
rect -12656 3507 -12640 3541
rect -12606 3507 -12590 3541
rect -12656 3466 -12590 3507
rect -12560 4425 -12494 4466
rect -12560 4391 -12544 4425
rect -12510 4391 -12494 4425
rect -12560 4357 -12494 4391
rect -12560 4323 -12544 4357
rect -12510 4323 -12494 4357
rect -12560 4289 -12494 4323
rect -12560 4255 -12544 4289
rect -12510 4255 -12494 4289
rect -12560 4221 -12494 4255
rect -12560 4187 -12544 4221
rect -12510 4187 -12494 4221
rect -12560 4153 -12494 4187
rect -12560 4119 -12544 4153
rect -12510 4119 -12494 4153
rect -12560 4085 -12494 4119
rect -12560 4051 -12544 4085
rect -12510 4051 -12494 4085
rect -12560 4017 -12494 4051
rect -12560 3983 -12544 4017
rect -12510 3983 -12494 4017
rect -12560 3949 -12494 3983
rect -12560 3915 -12544 3949
rect -12510 3915 -12494 3949
rect -12560 3881 -12494 3915
rect -12560 3847 -12544 3881
rect -12510 3847 -12494 3881
rect -12560 3813 -12494 3847
rect -12560 3779 -12544 3813
rect -12510 3779 -12494 3813
rect -12560 3745 -12494 3779
rect -12560 3711 -12544 3745
rect -12510 3711 -12494 3745
rect -12560 3677 -12494 3711
rect -12560 3643 -12544 3677
rect -12510 3643 -12494 3677
rect -12560 3609 -12494 3643
rect -12560 3575 -12544 3609
rect -12510 3575 -12494 3609
rect -12560 3541 -12494 3575
rect -12560 3507 -12544 3541
rect -12510 3507 -12494 3541
rect -12560 3466 -12494 3507
rect -12464 4425 -12398 4466
rect -12464 4391 -12448 4425
rect -12414 4391 -12398 4425
rect -12464 4357 -12398 4391
rect -12464 4323 -12448 4357
rect -12414 4323 -12398 4357
rect -12464 4289 -12398 4323
rect -12464 4255 -12448 4289
rect -12414 4255 -12398 4289
rect -12464 4221 -12398 4255
rect -12464 4187 -12448 4221
rect -12414 4187 -12398 4221
rect -12464 4153 -12398 4187
rect -12464 4119 -12448 4153
rect -12414 4119 -12398 4153
rect -12464 4085 -12398 4119
rect -12464 4051 -12448 4085
rect -12414 4051 -12398 4085
rect -12464 4017 -12398 4051
rect -12464 3983 -12448 4017
rect -12414 3983 -12398 4017
rect -12464 3949 -12398 3983
rect -12464 3915 -12448 3949
rect -12414 3915 -12398 3949
rect -12464 3881 -12398 3915
rect -12464 3847 -12448 3881
rect -12414 3847 -12398 3881
rect -12464 3813 -12398 3847
rect -12464 3779 -12448 3813
rect -12414 3779 -12398 3813
rect -12464 3745 -12398 3779
rect -12464 3711 -12448 3745
rect -12414 3711 -12398 3745
rect -12464 3677 -12398 3711
rect -12464 3643 -12448 3677
rect -12414 3643 -12398 3677
rect -12464 3609 -12398 3643
rect -12464 3575 -12448 3609
rect -12414 3575 -12398 3609
rect -12464 3541 -12398 3575
rect -12464 3507 -12448 3541
rect -12414 3507 -12398 3541
rect -12464 3466 -12398 3507
rect -12368 4425 -12302 4466
rect -12368 4391 -12352 4425
rect -12318 4391 -12302 4425
rect -12368 4357 -12302 4391
rect -12368 4323 -12352 4357
rect -12318 4323 -12302 4357
rect -12368 4289 -12302 4323
rect -12368 4255 -12352 4289
rect -12318 4255 -12302 4289
rect -12368 4221 -12302 4255
rect -12368 4187 -12352 4221
rect -12318 4187 -12302 4221
rect -12368 4153 -12302 4187
rect -12368 4119 -12352 4153
rect -12318 4119 -12302 4153
rect -12368 4085 -12302 4119
rect -12368 4051 -12352 4085
rect -12318 4051 -12302 4085
rect -12368 4017 -12302 4051
rect -12368 3983 -12352 4017
rect -12318 3983 -12302 4017
rect -12368 3949 -12302 3983
rect -12368 3915 -12352 3949
rect -12318 3915 -12302 3949
rect -12368 3881 -12302 3915
rect -12368 3847 -12352 3881
rect -12318 3847 -12302 3881
rect -12368 3813 -12302 3847
rect -12368 3779 -12352 3813
rect -12318 3779 -12302 3813
rect -12368 3745 -12302 3779
rect -12368 3711 -12352 3745
rect -12318 3711 -12302 3745
rect -12368 3677 -12302 3711
rect -12368 3643 -12352 3677
rect -12318 3643 -12302 3677
rect -12368 3609 -12302 3643
rect -12368 3575 -12352 3609
rect -12318 3575 -12302 3609
rect -12368 3541 -12302 3575
rect -12368 3507 -12352 3541
rect -12318 3507 -12302 3541
rect -12368 3466 -12302 3507
rect -12272 4425 -12206 4466
rect -12272 4391 -12256 4425
rect -12222 4391 -12206 4425
rect -12272 4357 -12206 4391
rect -12272 4323 -12256 4357
rect -12222 4323 -12206 4357
rect -12272 4289 -12206 4323
rect -12272 4255 -12256 4289
rect -12222 4255 -12206 4289
rect -12272 4221 -12206 4255
rect -12272 4187 -12256 4221
rect -12222 4187 -12206 4221
rect -12272 4153 -12206 4187
rect -12272 4119 -12256 4153
rect -12222 4119 -12206 4153
rect -12272 4085 -12206 4119
rect -12272 4051 -12256 4085
rect -12222 4051 -12206 4085
rect -12272 4017 -12206 4051
rect -12272 3983 -12256 4017
rect -12222 3983 -12206 4017
rect -12272 3949 -12206 3983
rect -12272 3915 -12256 3949
rect -12222 3915 -12206 3949
rect -12272 3881 -12206 3915
rect -12272 3847 -12256 3881
rect -12222 3847 -12206 3881
rect -12272 3813 -12206 3847
rect -12272 3779 -12256 3813
rect -12222 3779 -12206 3813
rect -12272 3745 -12206 3779
rect -12272 3711 -12256 3745
rect -12222 3711 -12206 3745
rect -12272 3677 -12206 3711
rect -12272 3643 -12256 3677
rect -12222 3643 -12206 3677
rect -12272 3609 -12206 3643
rect -12272 3575 -12256 3609
rect -12222 3575 -12206 3609
rect -12272 3541 -12206 3575
rect -12272 3507 -12256 3541
rect -12222 3507 -12206 3541
rect -12272 3466 -12206 3507
rect -12176 4425 -12110 4466
rect -12176 4391 -12160 4425
rect -12126 4391 -12110 4425
rect -12176 4357 -12110 4391
rect -12176 4323 -12160 4357
rect -12126 4323 -12110 4357
rect -12176 4289 -12110 4323
rect -12176 4255 -12160 4289
rect -12126 4255 -12110 4289
rect -12176 4221 -12110 4255
rect -12176 4187 -12160 4221
rect -12126 4187 -12110 4221
rect -12176 4153 -12110 4187
rect -12176 4119 -12160 4153
rect -12126 4119 -12110 4153
rect -12176 4085 -12110 4119
rect -12176 4051 -12160 4085
rect -12126 4051 -12110 4085
rect -12176 4017 -12110 4051
rect -12176 3983 -12160 4017
rect -12126 3983 -12110 4017
rect -12176 3949 -12110 3983
rect -12176 3915 -12160 3949
rect -12126 3915 -12110 3949
rect -12176 3881 -12110 3915
rect -12176 3847 -12160 3881
rect -12126 3847 -12110 3881
rect -12176 3813 -12110 3847
rect -12176 3779 -12160 3813
rect -12126 3779 -12110 3813
rect -12176 3745 -12110 3779
rect -12176 3711 -12160 3745
rect -12126 3711 -12110 3745
rect -12176 3677 -12110 3711
rect -12176 3643 -12160 3677
rect -12126 3643 -12110 3677
rect -12176 3609 -12110 3643
rect -12176 3575 -12160 3609
rect -12126 3575 -12110 3609
rect -12176 3541 -12110 3575
rect -12176 3507 -12160 3541
rect -12126 3507 -12110 3541
rect -12176 3466 -12110 3507
rect -12080 4425 -12014 4466
rect -12080 4391 -12064 4425
rect -12030 4391 -12014 4425
rect -12080 4357 -12014 4391
rect -12080 4323 -12064 4357
rect -12030 4323 -12014 4357
rect -12080 4289 -12014 4323
rect -12080 4255 -12064 4289
rect -12030 4255 -12014 4289
rect -12080 4221 -12014 4255
rect -12080 4187 -12064 4221
rect -12030 4187 -12014 4221
rect -12080 4153 -12014 4187
rect -12080 4119 -12064 4153
rect -12030 4119 -12014 4153
rect -12080 4085 -12014 4119
rect -12080 4051 -12064 4085
rect -12030 4051 -12014 4085
rect -12080 4017 -12014 4051
rect -12080 3983 -12064 4017
rect -12030 3983 -12014 4017
rect -12080 3949 -12014 3983
rect -12080 3915 -12064 3949
rect -12030 3915 -12014 3949
rect -12080 3881 -12014 3915
rect -12080 3847 -12064 3881
rect -12030 3847 -12014 3881
rect -12080 3813 -12014 3847
rect -12080 3779 -12064 3813
rect -12030 3779 -12014 3813
rect -12080 3745 -12014 3779
rect -12080 3711 -12064 3745
rect -12030 3711 -12014 3745
rect -12080 3677 -12014 3711
rect -12080 3643 -12064 3677
rect -12030 3643 -12014 3677
rect -12080 3609 -12014 3643
rect -12080 3575 -12064 3609
rect -12030 3575 -12014 3609
rect -12080 3541 -12014 3575
rect -12080 3507 -12064 3541
rect -12030 3507 -12014 3541
rect -12080 3466 -12014 3507
rect -11984 4425 -11922 4466
rect -11984 4391 -11968 4425
rect -11934 4391 -11922 4425
rect -11984 4357 -11922 4391
rect -11984 4323 -11968 4357
rect -11934 4323 -11922 4357
rect -11984 4289 -11922 4323
rect -11984 4255 -11968 4289
rect -11934 4255 -11922 4289
rect -11984 4221 -11922 4255
rect -11984 4187 -11968 4221
rect -11934 4187 -11922 4221
rect -11984 4153 -11922 4187
rect -11984 4119 -11968 4153
rect -11934 4119 -11922 4153
rect -11984 4085 -11922 4119
rect -11984 4051 -11968 4085
rect -11934 4051 -11922 4085
rect -11984 4017 -11922 4051
rect -11984 3983 -11968 4017
rect -11934 3983 -11922 4017
rect -11984 3949 -11922 3983
rect -11984 3915 -11968 3949
rect -11934 3915 -11922 3949
rect -11984 3881 -11922 3915
rect -11984 3847 -11968 3881
rect -11934 3847 -11922 3881
rect -11984 3813 -11922 3847
rect -11984 3779 -11968 3813
rect -11934 3779 -11922 3813
rect -11984 3745 -11922 3779
rect -11984 3711 -11968 3745
rect -11934 3711 -11922 3745
rect -11984 3677 -11922 3711
rect -11984 3643 -11968 3677
rect -11934 3643 -11922 3677
rect -11984 3609 -11922 3643
rect -11984 3575 -11968 3609
rect -11934 3575 -11922 3609
rect -11984 3541 -11922 3575
rect -11984 3507 -11968 3541
rect -11934 3507 -11922 3541
rect -11984 3466 -11922 3507
rect -11772 4427 -11710 4468
rect -11772 4393 -11760 4427
rect -11726 4393 -11710 4427
rect -11772 4359 -11710 4393
rect -11772 4325 -11760 4359
rect -11726 4325 -11710 4359
rect -11772 4291 -11710 4325
rect -11772 4257 -11760 4291
rect -11726 4257 -11710 4291
rect -11772 4223 -11710 4257
rect -11772 4189 -11760 4223
rect -11726 4189 -11710 4223
rect -11772 4155 -11710 4189
rect -11772 4121 -11760 4155
rect -11726 4121 -11710 4155
rect -11772 4087 -11710 4121
rect -11772 4053 -11760 4087
rect -11726 4053 -11710 4087
rect -11772 4019 -11710 4053
rect -11772 3985 -11760 4019
rect -11726 3985 -11710 4019
rect -11772 3951 -11710 3985
rect -11772 3917 -11760 3951
rect -11726 3917 -11710 3951
rect -11772 3883 -11710 3917
rect -11772 3849 -11760 3883
rect -11726 3849 -11710 3883
rect -11772 3815 -11710 3849
rect -11772 3781 -11760 3815
rect -11726 3781 -11710 3815
rect -11772 3747 -11710 3781
rect -11772 3713 -11760 3747
rect -11726 3713 -11710 3747
rect -11772 3679 -11710 3713
rect -11772 3645 -11760 3679
rect -11726 3645 -11710 3679
rect -11772 3611 -11710 3645
rect -11772 3577 -11760 3611
rect -11726 3577 -11710 3611
rect -11772 3543 -11710 3577
rect -11772 3509 -11760 3543
rect -11726 3509 -11710 3543
rect -11772 3468 -11710 3509
rect -11680 4427 -11614 4468
rect -11680 4393 -11664 4427
rect -11630 4393 -11614 4427
rect -11680 4359 -11614 4393
rect -11680 4325 -11664 4359
rect -11630 4325 -11614 4359
rect -11680 4291 -11614 4325
rect -11680 4257 -11664 4291
rect -11630 4257 -11614 4291
rect -11680 4223 -11614 4257
rect -11680 4189 -11664 4223
rect -11630 4189 -11614 4223
rect -11680 4155 -11614 4189
rect -11680 4121 -11664 4155
rect -11630 4121 -11614 4155
rect -11680 4087 -11614 4121
rect -11680 4053 -11664 4087
rect -11630 4053 -11614 4087
rect -11680 4019 -11614 4053
rect -11680 3985 -11664 4019
rect -11630 3985 -11614 4019
rect -11680 3951 -11614 3985
rect -11680 3917 -11664 3951
rect -11630 3917 -11614 3951
rect -11680 3883 -11614 3917
rect -11680 3849 -11664 3883
rect -11630 3849 -11614 3883
rect -11680 3815 -11614 3849
rect -11680 3781 -11664 3815
rect -11630 3781 -11614 3815
rect -11680 3747 -11614 3781
rect -11680 3713 -11664 3747
rect -11630 3713 -11614 3747
rect -11680 3679 -11614 3713
rect -11680 3645 -11664 3679
rect -11630 3645 -11614 3679
rect -11680 3611 -11614 3645
rect -11680 3577 -11664 3611
rect -11630 3577 -11614 3611
rect -11680 3543 -11614 3577
rect -11680 3509 -11664 3543
rect -11630 3509 -11614 3543
rect -11680 3468 -11614 3509
rect -11584 4427 -11518 4468
rect -11584 4393 -11568 4427
rect -11534 4393 -11518 4427
rect -11584 4359 -11518 4393
rect -11584 4325 -11568 4359
rect -11534 4325 -11518 4359
rect -11584 4291 -11518 4325
rect -11584 4257 -11568 4291
rect -11534 4257 -11518 4291
rect -11584 4223 -11518 4257
rect -11584 4189 -11568 4223
rect -11534 4189 -11518 4223
rect -11584 4155 -11518 4189
rect -11584 4121 -11568 4155
rect -11534 4121 -11518 4155
rect -11584 4087 -11518 4121
rect -11584 4053 -11568 4087
rect -11534 4053 -11518 4087
rect -11584 4019 -11518 4053
rect -11584 3985 -11568 4019
rect -11534 3985 -11518 4019
rect -11584 3951 -11518 3985
rect -11584 3917 -11568 3951
rect -11534 3917 -11518 3951
rect -11584 3883 -11518 3917
rect -11584 3849 -11568 3883
rect -11534 3849 -11518 3883
rect -11584 3815 -11518 3849
rect -11584 3781 -11568 3815
rect -11534 3781 -11518 3815
rect -11584 3747 -11518 3781
rect -11584 3713 -11568 3747
rect -11534 3713 -11518 3747
rect -11584 3679 -11518 3713
rect -11584 3645 -11568 3679
rect -11534 3645 -11518 3679
rect -11584 3611 -11518 3645
rect -11584 3577 -11568 3611
rect -11534 3577 -11518 3611
rect -11584 3543 -11518 3577
rect -11584 3509 -11568 3543
rect -11534 3509 -11518 3543
rect -11584 3468 -11518 3509
rect -11488 4427 -11422 4468
rect -11488 4393 -11472 4427
rect -11438 4393 -11422 4427
rect -11488 4359 -11422 4393
rect -11488 4325 -11472 4359
rect -11438 4325 -11422 4359
rect -11488 4291 -11422 4325
rect -11488 4257 -11472 4291
rect -11438 4257 -11422 4291
rect -11488 4223 -11422 4257
rect -11488 4189 -11472 4223
rect -11438 4189 -11422 4223
rect -11488 4155 -11422 4189
rect -11488 4121 -11472 4155
rect -11438 4121 -11422 4155
rect -11488 4087 -11422 4121
rect -11488 4053 -11472 4087
rect -11438 4053 -11422 4087
rect -11488 4019 -11422 4053
rect -11488 3985 -11472 4019
rect -11438 3985 -11422 4019
rect -11488 3951 -11422 3985
rect -11488 3917 -11472 3951
rect -11438 3917 -11422 3951
rect -11488 3883 -11422 3917
rect -11488 3849 -11472 3883
rect -11438 3849 -11422 3883
rect -11488 3815 -11422 3849
rect -11488 3781 -11472 3815
rect -11438 3781 -11422 3815
rect -11488 3747 -11422 3781
rect -11488 3713 -11472 3747
rect -11438 3713 -11422 3747
rect -11488 3679 -11422 3713
rect -11488 3645 -11472 3679
rect -11438 3645 -11422 3679
rect -11488 3611 -11422 3645
rect -11488 3577 -11472 3611
rect -11438 3577 -11422 3611
rect -11488 3543 -11422 3577
rect -11488 3509 -11472 3543
rect -11438 3509 -11422 3543
rect -11488 3468 -11422 3509
rect -11392 4427 -11326 4468
rect -11392 4393 -11376 4427
rect -11342 4393 -11326 4427
rect -11392 4359 -11326 4393
rect -11392 4325 -11376 4359
rect -11342 4325 -11326 4359
rect -11392 4291 -11326 4325
rect -11392 4257 -11376 4291
rect -11342 4257 -11326 4291
rect -11392 4223 -11326 4257
rect -11392 4189 -11376 4223
rect -11342 4189 -11326 4223
rect -11392 4155 -11326 4189
rect -11392 4121 -11376 4155
rect -11342 4121 -11326 4155
rect -11392 4087 -11326 4121
rect -11392 4053 -11376 4087
rect -11342 4053 -11326 4087
rect -11392 4019 -11326 4053
rect -11392 3985 -11376 4019
rect -11342 3985 -11326 4019
rect -11392 3951 -11326 3985
rect -11392 3917 -11376 3951
rect -11342 3917 -11326 3951
rect -11392 3883 -11326 3917
rect -11392 3849 -11376 3883
rect -11342 3849 -11326 3883
rect -11392 3815 -11326 3849
rect -11392 3781 -11376 3815
rect -11342 3781 -11326 3815
rect -11392 3747 -11326 3781
rect -11392 3713 -11376 3747
rect -11342 3713 -11326 3747
rect -11392 3679 -11326 3713
rect -11392 3645 -11376 3679
rect -11342 3645 -11326 3679
rect -11392 3611 -11326 3645
rect -11392 3577 -11376 3611
rect -11342 3577 -11326 3611
rect -11392 3543 -11326 3577
rect -11392 3509 -11376 3543
rect -11342 3509 -11326 3543
rect -11392 3468 -11326 3509
rect -11296 4427 -11234 4468
rect -11296 4393 -11280 4427
rect -11246 4393 -11234 4427
rect -11296 4359 -11234 4393
rect -11296 4325 -11280 4359
rect -11246 4325 -11234 4359
rect -11296 4291 -11234 4325
rect -11296 4257 -11280 4291
rect -11246 4257 -11234 4291
rect -11296 4223 -11234 4257
rect -11296 4189 -11280 4223
rect -11246 4189 -11234 4223
rect -11296 4155 -11234 4189
rect -11296 4121 -11280 4155
rect -11246 4121 -11234 4155
rect -11296 4087 -11234 4121
rect -11296 4053 -11280 4087
rect -11246 4053 -11234 4087
rect -11296 4019 -11234 4053
rect -11296 3985 -11280 4019
rect -11246 3985 -11234 4019
rect -11296 3951 -11234 3985
rect -11296 3917 -11280 3951
rect -11246 3917 -11234 3951
rect -11296 3883 -11234 3917
rect -11296 3849 -11280 3883
rect -11246 3849 -11234 3883
rect -11296 3815 -11234 3849
rect -11296 3781 -11280 3815
rect -11246 3781 -11234 3815
rect -11296 3747 -11234 3781
rect -11296 3713 -11280 3747
rect -11246 3713 -11234 3747
rect -11296 3679 -11234 3713
rect -11296 3645 -11280 3679
rect -11246 3645 -11234 3679
rect -11296 3611 -11234 3645
rect -11296 3577 -11280 3611
rect -11246 3577 -11234 3611
rect -11296 3543 -11234 3577
rect -11296 3509 -11280 3543
rect -11246 3509 -11234 3543
rect -11296 3468 -11234 3509
rect -10302 4411 -10240 4452
rect -10302 4377 -10290 4411
rect -10256 4377 -10240 4411
rect -10302 4343 -10240 4377
rect -10302 4309 -10290 4343
rect -10256 4309 -10240 4343
rect -10302 4275 -10240 4309
rect -10302 4241 -10290 4275
rect -10256 4241 -10240 4275
rect -10302 4207 -10240 4241
rect -10302 4173 -10290 4207
rect -10256 4173 -10240 4207
rect -10302 4139 -10240 4173
rect -10302 4105 -10290 4139
rect -10256 4105 -10240 4139
rect -10302 4071 -10240 4105
rect -10302 4037 -10290 4071
rect -10256 4037 -10240 4071
rect -10302 4003 -10240 4037
rect -10302 3969 -10290 4003
rect -10256 3969 -10240 4003
rect -10302 3935 -10240 3969
rect -10302 3901 -10290 3935
rect -10256 3901 -10240 3935
rect -10302 3867 -10240 3901
rect -10302 3833 -10290 3867
rect -10256 3833 -10240 3867
rect -10302 3799 -10240 3833
rect -10302 3765 -10290 3799
rect -10256 3765 -10240 3799
rect -10302 3731 -10240 3765
rect -10302 3697 -10290 3731
rect -10256 3697 -10240 3731
rect -10302 3663 -10240 3697
rect -10302 3629 -10290 3663
rect -10256 3629 -10240 3663
rect -10302 3595 -10240 3629
rect -10302 3561 -10290 3595
rect -10256 3561 -10240 3595
rect -10302 3527 -10240 3561
rect -10302 3493 -10290 3527
rect -10256 3493 -10240 3527
rect -10302 3452 -10240 3493
rect -10210 4411 -10144 4452
rect -10210 4377 -10194 4411
rect -10160 4377 -10144 4411
rect -10210 4343 -10144 4377
rect -10210 4309 -10194 4343
rect -10160 4309 -10144 4343
rect -10210 4275 -10144 4309
rect -10210 4241 -10194 4275
rect -10160 4241 -10144 4275
rect -10210 4207 -10144 4241
rect -10210 4173 -10194 4207
rect -10160 4173 -10144 4207
rect -10210 4139 -10144 4173
rect -10210 4105 -10194 4139
rect -10160 4105 -10144 4139
rect -10210 4071 -10144 4105
rect -10210 4037 -10194 4071
rect -10160 4037 -10144 4071
rect -10210 4003 -10144 4037
rect -10210 3969 -10194 4003
rect -10160 3969 -10144 4003
rect -10210 3935 -10144 3969
rect -10210 3901 -10194 3935
rect -10160 3901 -10144 3935
rect -10210 3867 -10144 3901
rect -10210 3833 -10194 3867
rect -10160 3833 -10144 3867
rect -10210 3799 -10144 3833
rect -10210 3765 -10194 3799
rect -10160 3765 -10144 3799
rect -10210 3731 -10144 3765
rect -10210 3697 -10194 3731
rect -10160 3697 -10144 3731
rect -10210 3663 -10144 3697
rect -10210 3629 -10194 3663
rect -10160 3629 -10144 3663
rect -10210 3595 -10144 3629
rect -10210 3561 -10194 3595
rect -10160 3561 -10144 3595
rect -10210 3527 -10144 3561
rect -10210 3493 -10194 3527
rect -10160 3493 -10144 3527
rect -10210 3452 -10144 3493
rect -10114 4411 -10048 4452
rect -10114 4377 -10098 4411
rect -10064 4377 -10048 4411
rect -10114 4343 -10048 4377
rect -10114 4309 -10098 4343
rect -10064 4309 -10048 4343
rect -10114 4275 -10048 4309
rect -10114 4241 -10098 4275
rect -10064 4241 -10048 4275
rect -10114 4207 -10048 4241
rect -10114 4173 -10098 4207
rect -10064 4173 -10048 4207
rect -10114 4139 -10048 4173
rect -10114 4105 -10098 4139
rect -10064 4105 -10048 4139
rect -10114 4071 -10048 4105
rect -10114 4037 -10098 4071
rect -10064 4037 -10048 4071
rect -10114 4003 -10048 4037
rect -10114 3969 -10098 4003
rect -10064 3969 -10048 4003
rect -10114 3935 -10048 3969
rect -10114 3901 -10098 3935
rect -10064 3901 -10048 3935
rect -10114 3867 -10048 3901
rect -10114 3833 -10098 3867
rect -10064 3833 -10048 3867
rect -10114 3799 -10048 3833
rect -10114 3765 -10098 3799
rect -10064 3765 -10048 3799
rect -10114 3731 -10048 3765
rect -10114 3697 -10098 3731
rect -10064 3697 -10048 3731
rect -10114 3663 -10048 3697
rect -10114 3629 -10098 3663
rect -10064 3629 -10048 3663
rect -10114 3595 -10048 3629
rect -10114 3561 -10098 3595
rect -10064 3561 -10048 3595
rect -10114 3527 -10048 3561
rect -10114 3493 -10098 3527
rect -10064 3493 -10048 3527
rect -10114 3452 -10048 3493
rect -10018 4411 -9952 4452
rect -10018 4377 -10002 4411
rect -9968 4377 -9952 4411
rect -10018 4343 -9952 4377
rect -10018 4309 -10002 4343
rect -9968 4309 -9952 4343
rect -10018 4275 -9952 4309
rect -10018 4241 -10002 4275
rect -9968 4241 -9952 4275
rect -10018 4207 -9952 4241
rect -10018 4173 -10002 4207
rect -9968 4173 -9952 4207
rect -10018 4139 -9952 4173
rect -10018 4105 -10002 4139
rect -9968 4105 -9952 4139
rect -10018 4071 -9952 4105
rect -10018 4037 -10002 4071
rect -9968 4037 -9952 4071
rect -10018 4003 -9952 4037
rect -10018 3969 -10002 4003
rect -9968 3969 -9952 4003
rect -10018 3935 -9952 3969
rect -10018 3901 -10002 3935
rect -9968 3901 -9952 3935
rect -10018 3867 -9952 3901
rect -10018 3833 -10002 3867
rect -9968 3833 -9952 3867
rect -10018 3799 -9952 3833
rect -10018 3765 -10002 3799
rect -9968 3765 -9952 3799
rect -10018 3731 -9952 3765
rect -10018 3697 -10002 3731
rect -9968 3697 -9952 3731
rect -10018 3663 -9952 3697
rect -10018 3629 -10002 3663
rect -9968 3629 -9952 3663
rect -10018 3595 -9952 3629
rect -10018 3561 -10002 3595
rect -9968 3561 -9952 3595
rect -10018 3527 -9952 3561
rect -10018 3493 -10002 3527
rect -9968 3493 -9952 3527
rect -10018 3452 -9952 3493
rect -9922 4411 -9856 4452
rect -9922 4377 -9906 4411
rect -9872 4377 -9856 4411
rect -9922 4343 -9856 4377
rect -9922 4309 -9906 4343
rect -9872 4309 -9856 4343
rect -9922 4275 -9856 4309
rect -9922 4241 -9906 4275
rect -9872 4241 -9856 4275
rect -9922 4207 -9856 4241
rect -9922 4173 -9906 4207
rect -9872 4173 -9856 4207
rect -9922 4139 -9856 4173
rect -9922 4105 -9906 4139
rect -9872 4105 -9856 4139
rect -9922 4071 -9856 4105
rect -9922 4037 -9906 4071
rect -9872 4037 -9856 4071
rect -9922 4003 -9856 4037
rect -9922 3969 -9906 4003
rect -9872 3969 -9856 4003
rect -9922 3935 -9856 3969
rect -9922 3901 -9906 3935
rect -9872 3901 -9856 3935
rect -9922 3867 -9856 3901
rect -9922 3833 -9906 3867
rect -9872 3833 -9856 3867
rect -9922 3799 -9856 3833
rect -9922 3765 -9906 3799
rect -9872 3765 -9856 3799
rect -9922 3731 -9856 3765
rect -9922 3697 -9906 3731
rect -9872 3697 -9856 3731
rect -9922 3663 -9856 3697
rect -9922 3629 -9906 3663
rect -9872 3629 -9856 3663
rect -9922 3595 -9856 3629
rect -9922 3561 -9906 3595
rect -9872 3561 -9856 3595
rect -9922 3527 -9856 3561
rect -9922 3493 -9906 3527
rect -9872 3493 -9856 3527
rect -9922 3452 -9856 3493
rect -9826 4411 -9760 4452
rect -9826 4377 -9810 4411
rect -9776 4377 -9760 4411
rect -9826 4343 -9760 4377
rect -9826 4309 -9810 4343
rect -9776 4309 -9760 4343
rect -9826 4275 -9760 4309
rect -9826 4241 -9810 4275
rect -9776 4241 -9760 4275
rect -9826 4207 -9760 4241
rect -9826 4173 -9810 4207
rect -9776 4173 -9760 4207
rect -9826 4139 -9760 4173
rect -9826 4105 -9810 4139
rect -9776 4105 -9760 4139
rect -9826 4071 -9760 4105
rect -9826 4037 -9810 4071
rect -9776 4037 -9760 4071
rect -9826 4003 -9760 4037
rect -9826 3969 -9810 4003
rect -9776 3969 -9760 4003
rect -9826 3935 -9760 3969
rect -9826 3901 -9810 3935
rect -9776 3901 -9760 3935
rect -9826 3867 -9760 3901
rect -9826 3833 -9810 3867
rect -9776 3833 -9760 3867
rect -9826 3799 -9760 3833
rect -9826 3765 -9810 3799
rect -9776 3765 -9760 3799
rect -9826 3731 -9760 3765
rect -9826 3697 -9810 3731
rect -9776 3697 -9760 3731
rect -9826 3663 -9760 3697
rect -9826 3629 -9810 3663
rect -9776 3629 -9760 3663
rect -9826 3595 -9760 3629
rect -9826 3561 -9810 3595
rect -9776 3561 -9760 3595
rect -9826 3527 -9760 3561
rect -9826 3493 -9810 3527
rect -9776 3493 -9760 3527
rect -9826 3452 -9760 3493
rect -9730 4411 -9664 4452
rect -9730 4377 -9714 4411
rect -9680 4377 -9664 4411
rect -9730 4343 -9664 4377
rect -9730 4309 -9714 4343
rect -9680 4309 -9664 4343
rect -9730 4275 -9664 4309
rect -9730 4241 -9714 4275
rect -9680 4241 -9664 4275
rect -9730 4207 -9664 4241
rect -9730 4173 -9714 4207
rect -9680 4173 -9664 4207
rect -9730 4139 -9664 4173
rect -9730 4105 -9714 4139
rect -9680 4105 -9664 4139
rect -9730 4071 -9664 4105
rect -9730 4037 -9714 4071
rect -9680 4037 -9664 4071
rect -9730 4003 -9664 4037
rect -9730 3969 -9714 4003
rect -9680 3969 -9664 4003
rect -9730 3935 -9664 3969
rect -9730 3901 -9714 3935
rect -9680 3901 -9664 3935
rect -9730 3867 -9664 3901
rect -9730 3833 -9714 3867
rect -9680 3833 -9664 3867
rect -9730 3799 -9664 3833
rect -9730 3765 -9714 3799
rect -9680 3765 -9664 3799
rect -9730 3731 -9664 3765
rect -9730 3697 -9714 3731
rect -9680 3697 -9664 3731
rect -9730 3663 -9664 3697
rect -9730 3629 -9714 3663
rect -9680 3629 -9664 3663
rect -9730 3595 -9664 3629
rect -9730 3561 -9714 3595
rect -9680 3561 -9664 3595
rect -9730 3527 -9664 3561
rect -9730 3493 -9714 3527
rect -9680 3493 -9664 3527
rect -9730 3452 -9664 3493
rect -9634 4411 -9568 4452
rect -9634 4377 -9618 4411
rect -9584 4377 -9568 4411
rect -9634 4343 -9568 4377
rect -9634 4309 -9618 4343
rect -9584 4309 -9568 4343
rect -9634 4275 -9568 4309
rect -9634 4241 -9618 4275
rect -9584 4241 -9568 4275
rect -9634 4207 -9568 4241
rect -9634 4173 -9618 4207
rect -9584 4173 -9568 4207
rect -9634 4139 -9568 4173
rect -9634 4105 -9618 4139
rect -9584 4105 -9568 4139
rect -9634 4071 -9568 4105
rect -9634 4037 -9618 4071
rect -9584 4037 -9568 4071
rect -9634 4003 -9568 4037
rect -9634 3969 -9618 4003
rect -9584 3969 -9568 4003
rect -9634 3935 -9568 3969
rect -9634 3901 -9618 3935
rect -9584 3901 -9568 3935
rect -9634 3867 -9568 3901
rect -9634 3833 -9618 3867
rect -9584 3833 -9568 3867
rect -9634 3799 -9568 3833
rect -9634 3765 -9618 3799
rect -9584 3765 -9568 3799
rect -9634 3731 -9568 3765
rect -9634 3697 -9618 3731
rect -9584 3697 -9568 3731
rect -9634 3663 -9568 3697
rect -9634 3629 -9618 3663
rect -9584 3629 -9568 3663
rect -9634 3595 -9568 3629
rect -9634 3561 -9618 3595
rect -9584 3561 -9568 3595
rect -9634 3527 -9568 3561
rect -9634 3493 -9618 3527
rect -9584 3493 -9568 3527
rect -9634 3452 -9568 3493
rect -9538 4411 -9472 4452
rect -9538 4377 -9522 4411
rect -9488 4377 -9472 4411
rect -9538 4343 -9472 4377
rect -9538 4309 -9522 4343
rect -9488 4309 -9472 4343
rect -9538 4275 -9472 4309
rect -9538 4241 -9522 4275
rect -9488 4241 -9472 4275
rect -9538 4207 -9472 4241
rect -9538 4173 -9522 4207
rect -9488 4173 -9472 4207
rect -9538 4139 -9472 4173
rect -9538 4105 -9522 4139
rect -9488 4105 -9472 4139
rect -9538 4071 -9472 4105
rect -9538 4037 -9522 4071
rect -9488 4037 -9472 4071
rect -9538 4003 -9472 4037
rect -9538 3969 -9522 4003
rect -9488 3969 -9472 4003
rect -9538 3935 -9472 3969
rect -9538 3901 -9522 3935
rect -9488 3901 -9472 3935
rect -9538 3867 -9472 3901
rect -9538 3833 -9522 3867
rect -9488 3833 -9472 3867
rect -9538 3799 -9472 3833
rect -9538 3765 -9522 3799
rect -9488 3765 -9472 3799
rect -9538 3731 -9472 3765
rect -9538 3697 -9522 3731
rect -9488 3697 -9472 3731
rect -9538 3663 -9472 3697
rect -9538 3629 -9522 3663
rect -9488 3629 -9472 3663
rect -9538 3595 -9472 3629
rect -9538 3561 -9522 3595
rect -9488 3561 -9472 3595
rect -9538 3527 -9472 3561
rect -9538 3493 -9522 3527
rect -9488 3493 -9472 3527
rect -9538 3452 -9472 3493
rect -9442 4411 -9376 4452
rect -9442 4377 -9426 4411
rect -9392 4377 -9376 4411
rect -9442 4343 -9376 4377
rect -9442 4309 -9426 4343
rect -9392 4309 -9376 4343
rect -9442 4275 -9376 4309
rect -9442 4241 -9426 4275
rect -9392 4241 -9376 4275
rect -9442 4207 -9376 4241
rect -9442 4173 -9426 4207
rect -9392 4173 -9376 4207
rect -9442 4139 -9376 4173
rect -9442 4105 -9426 4139
rect -9392 4105 -9376 4139
rect -9442 4071 -9376 4105
rect -9442 4037 -9426 4071
rect -9392 4037 -9376 4071
rect -9442 4003 -9376 4037
rect -9442 3969 -9426 4003
rect -9392 3969 -9376 4003
rect -9442 3935 -9376 3969
rect -9442 3901 -9426 3935
rect -9392 3901 -9376 3935
rect -9442 3867 -9376 3901
rect -9442 3833 -9426 3867
rect -9392 3833 -9376 3867
rect -9442 3799 -9376 3833
rect -9442 3765 -9426 3799
rect -9392 3765 -9376 3799
rect -9442 3731 -9376 3765
rect -9442 3697 -9426 3731
rect -9392 3697 -9376 3731
rect -9442 3663 -9376 3697
rect -9442 3629 -9426 3663
rect -9392 3629 -9376 3663
rect -9442 3595 -9376 3629
rect -9442 3561 -9426 3595
rect -9392 3561 -9376 3595
rect -9442 3527 -9376 3561
rect -9442 3493 -9426 3527
rect -9392 3493 -9376 3527
rect -9442 3452 -9376 3493
rect -9346 4411 -9280 4452
rect -9346 4377 -9330 4411
rect -9296 4377 -9280 4411
rect -9346 4343 -9280 4377
rect -9346 4309 -9330 4343
rect -9296 4309 -9280 4343
rect -9346 4275 -9280 4309
rect -9346 4241 -9330 4275
rect -9296 4241 -9280 4275
rect -9346 4207 -9280 4241
rect -9346 4173 -9330 4207
rect -9296 4173 -9280 4207
rect -9346 4139 -9280 4173
rect -9346 4105 -9330 4139
rect -9296 4105 -9280 4139
rect -9346 4071 -9280 4105
rect -9346 4037 -9330 4071
rect -9296 4037 -9280 4071
rect -9346 4003 -9280 4037
rect -9346 3969 -9330 4003
rect -9296 3969 -9280 4003
rect -9346 3935 -9280 3969
rect -9346 3901 -9330 3935
rect -9296 3901 -9280 3935
rect -9346 3867 -9280 3901
rect -9346 3833 -9330 3867
rect -9296 3833 -9280 3867
rect -9346 3799 -9280 3833
rect -9346 3765 -9330 3799
rect -9296 3765 -9280 3799
rect -9346 3731 -9280 3765
rect -9346 3697 -9330 3731
rect -9296 3697 -9280 3731
rect -9346 3663 -9280 3697
rect -9346 3629 -9330 3663
rect -9296 3629 -9280 3663
rect -9346 3595 -9280 3629
rect -9346 3561 -9330 3595
rect -9296 3561 -9280 3595
rect -9346 3527 -9280 3561
rect -9346 3493 -9330 3527
rect -9296 3493 -9280 3527
rect -9346 3452 -9280 3493
rect -9250 4411 -9184 4452
rect -9250 4377 -9234 4411
rect -9200 4377 -9184 4411
rect -9250 4343 -9184 4377
rect -9250 4309 -9234 4343
rect -9200 4309 -9184 4343
rect -9250 4275 -9184 4309
rect -9250 4241 -9234 4275
rect -9200 4241 -9184 4275
rect -9250 4207 -9184 4241
rect -9250 4173 -9234 4207
rect -9200 4173 -9184 4207
rect -9250 4139 -9184 4173
rect -9250 4105 -9234 4139
rect -9200 4105 -9184 4139
rect -9250 4071 -9184 4105
rect -9250 4037 -9234 4071
rect -9200 4037 -9184 4071
rect -9250 4003 -9184 4037
rect -9250 3969 -9234 4003
rect -9200 3969 -9184 4003
rect -9250 3935 -9184 3969
rect -9250 3901 -9234 3935
rect -9200 3901 -9184 3935
rect -9250 3867 -9184 3901
rect -9250 3833 -9234 3867
rect -9200 3833 -9184 3867
rect -9250 3799 -9184 3833
rect -9250 3765 -9234 3799
rect -9200 3765 -9184 3799
rect -9250 3731 -9184 3765
rect -9250 3697 -9234 3731
rect -9200 3697 -9184 3731
rect -9250 3663 -9184 3697
rect -9250 3629 -9234 3663
rect -9200 3629 -9184 3663
rect -9250 3595 -9184 3629
rect -9250 3561 -9234 3595
rect -9200 3561 -9184 3595
rect -9250 3527 -9184 3561
rect -9250 3493 -9234 3527
rect -9200 3493 -9184 3527
rect -9250 3452 -9184 3493
rect -9154 4411 -9088 4452
rect -9154 4377 -9138 4411
rect -9104 4377 -9088 4411
rect -9154 4343 -9088 4377
rect -9154 4309 -9138 4343
rect -9104 4309 -9088 4343
rect -9154 4275 -9088 4309
rect -9154 4241 -9138 4275
rect -9104 4241 -9088 4275
rect -9154 4207 -9088 4241
rect -9154 4173 -9138 4207
rect -9104 4173 -9088 4207
rect -9154 4139 -9088 4173
rect -9154 4105 -9138 4139
rect -9104 4105 -9088 4139
rect -9154 4071 -9088 4105
rect -9154 4037 -9138 4071
rect -9104 4037 -9088 4071
rect -9154 4003 -9088 4037
rect -9154 3969 -9138 4003
rect -9104 3969 -9088 4003
rect -9154 3935 -9088 3969
rect -9154 3901 -9138 3935
rect -9104 3901 -9088 3935
rect -9154 3867 -9088 3901
rect -9154 3833 -9138 3867
rect -9104 3833 -9088 3867
rect -9154 3799 -9088 3833
rect -9154 3765 -9138 3799
rect -9104 3765 -9088 3799
rect -9154 3731 -9088 3765
rect -9154 3697 -9138 3731
rect -9104 3697 -9088 3731
rect -9154 3663 -9088 3697
rect -9154 3629 -9138 3663
rect -9104 3629 -9088 3663
rect -9154 3595 -9088 3629
rect -9154 3561 -9138 3595
rect -9104 3561 -9088 3595
rect -9154 3527 -9088 3561
rect -9154 3493 -9138 3527
rect -9104 3493 -9088 3527
rect -9154 3452 -9088 3493
rect -9058 4411 -8992 4452
rect -9058 4377 -9042 4411
rect -9008 4377 -8992 4411
rect -9058 4343 -8992 4377
rect -9058 4309 -9042 4343
rect -9008 4309 -8992 4343
rect -9058 4275 -8992 4309
rect -9058 4241 -9042 4275
rect -9008 4241 -8992 4275
rect -9058 4207 -8992 4241
rect -9058 4173 -9042 4207
rect -9008 4173 -8992 4207
rect -9058 4139 -8992 4173
rect -9058 4105 -9042 4139
rect -9008 4105 -8992 4139
rect -9058 4071 -8992 4105
rect -9058 4037 -9042 4071
rect -9008 4037 -8992 4071
rect -9058 4003 -8992 4037
rect -9058 3969 -9042 4003
rect -9008 3969 -8992 4003
rect -9058 3935 -8992 3969
rect -9058 3901 -9042 3935
rect -9008 3901 -8992 3935
rect -9058 3867 -8992 3901
rect -9058 3833 -9042 3867
rect -9008 3833 -8992 3867
rect -9058 3799 -8992 3833
rect -9058 3765 -9042 3799
rect -9008 3765 -8992 3799
rect -9058 3731 -8992 3765
rect -9058 3697 -9042 3731
rect -9008 3697 -8992 3731
rect -9058 3663 -8992 3697
rect -9058 3629 -9042 3663
rect -9008 3629 -8992 3663
rect -9058 3595 -8992 3629
rect -9058 3561 -9042 3595
rect -9008 3561 -8992 3595
rect -9058 3527 -8992 3561
rect -9058 3493 -9042 3527
rect -9008 3493 -8992 3527
rect -9058 3452 -8992 3493
rect -8962 4411 -8896 4452
rect -8962 4377 -8946 4411
rect -8912 4377 -8896 4411
rect -8962 4343 -8896 4377
rect -8962 4309 -8946 4343
rect -8912 4309 -8896 4343
rect -8962 4275 -8896 4309
rect -8962 4241 -8946 4275
rect -8912 4241 -8896 4275
rect -8962 4207 -8896 4241
rect -8962 4173 -8946 4207
rect -8912 4173 -8896 4207
rect -8962 4139 -8896 4173
rect -8962 4105 -8946 4139
rect -8912 4105 -8896 4139
rect -8962 4071 -8896 4105
rect -8962 4037 -8946 4071
rect -8912 4037 -8896 4071
rect -8962 4003 -8896 4037
rect -8962 3969 -8946 4003
rect -8912 3969 -8896 4003
rect -8962 3935 -8896 3969
rect -8962 3901 -8946 3935
rect -8912 3901 -8896 3935
rect -8962 3867 -8896 3901
rect -8962 3833 -8946 3867
rect -8912 3833 -8896 3867
rect -8962 3799 -8896 3833
rect -8962 3765 -8946 3799
rect -8912 3765 -8896 3799
rect -8962 3731 -8896 3765
rect -8962 3697 -8946 3731
rect -8912 3697 -8896 3731
rect -8962 3663 -8896 3697
rect -8962 3629 -8946 3663
rect -8912 3629 -8896 3663
rect -8962 3595 -8896 3629
rect -8962 3561 -8946 3595
rect -8912 3561 -8896 3595
rect -8962 3527 -8896 3561
rect -8962 3493 -8946 3527
rect -8912 3493 -8896 3527
rect -8962 3452 -8896 3493
rect -8866 4411 -8800 4452
rect -8866 4377 -8850 4411
rect -8816 4377 -8800 4411
rect -8866 4343 -8800 4377
rect -8866 4309 -8850 4343
rect -8816 4309 -8800 4343
rect -8866 4275 -8800 4309
rect -8866 4241 -8850 4275
rect -8816 4241 -8800 4275
rect -8866 4207 -8800 4241
rect -8866 4173 -8850 4207
rect -8816 4173 -8800 4207
rect -8866 4139 -8800 4173
rect -8866 4105 -8850 4139
rect -8816 4105 -8800 4139
rect -8866 4071 -8800 4105
rect -8866 4037 -8850 4071
rect -8816 4037 -8800 4071
rect -8866 4003 -8800 4037
rect -8866 3969 -8850 4003
rect -8816 3969 -8800 4003
rect -8866 3935 -8800 3969
rect -8866 3901 -8850 3935
rect -8816 3901 -8800 3935
rect -8866 3867 -8800 3901
rect -8866 3833 -8850 3867
rect -8816 3833 -8800 3867
rect -8866 3799 -8800 3833
rect -8866 3765 -8850 3799
rect -8816 3765 -8800 3799
rect -8866 3731 -8800 3765
rect -8866 3697 -8850 3731
rect -8816 3697 -8800 3731
rect -8866 3663 -8800 3697
rect -8866 3629 -8850 3663
rect -8816 3629 -8800 3663
rect -8866 3595 -8800 3629
rect -8866 3561 -8850 3595
rect -8816 3561 -8800 3595
rect -8866 3527 -8800 3561
rect -8866 3493 -8850 3527
rect -8816 3493 -8800 3527
rect -8866 3452 -8800 3493
rect -8770 4411 -8704 4452
rect -8770 4377 -8754 4411
rect -8720 4377 -8704 4411
rect -8770 4343 -8704 4377
rect -8770 4309 -8754 4343
rect -8720 4309 -8704 4343
rect -8770 4275 -8704 4309
rect -8770 4241 -8754 4275
rect -8720 4241 -8704 4275
rect -8770 4207 -8704 4241
rect -8770 4173 -8754 4207
rect -8720 4173 -8704 4207
rect -8770 4139 -8704 4173
rect -8770 4105 -8754 4139
rect -8720 4105 -8704 4139
rect -8770 4071 -8704 4105
rect -8770 4037 -8754 4071
rect -8720 4037 -8704 4071
rect -8770 4003 -8704 4037
rect -8770 3969 -8754 4003
rect -8720 3969 -8704 4003
rect -8770 3935 -8704 3969
rect -8770 3901 -8754 3935
rect -8720 3901 -8704 3935
rect -8770 3867 -8704 3901
rect -8770 3833 -8754 3867
rect -8720 3833 -8704 3867
rect -8770 3799 -8704 3833
rect -8770 3765 -8754 3799
rect -8720 3765 -8704 3799
rect -8770 3731 -8704 3765
rect -8770 3697 -8754 3731
rect -8720 3697 -8704 3731
rect -8770 3663 -8704 3697
rect -8770 3629 -8754 3663
rect -8720 3629 -8704 3663
rect -8770 3595 -8704 3629
rect -8770 3561 -8754 3595
rect -8720 3561 -8704 3595
rect -8770 3527 -8704 3561
rect -8770 3493 -8754 3527
rect -8720 3493 -8704 3527
rect -8770 3452 -8704 3493
rect -8674 4411 -8608 4452
rect -8674 4377 -8658 4411
rect -8624 4377 -8608 4411
rect -8674 4343 -8608 4377
rect -8674 4309 -8658 4343
rect -8624 4309 -8608 4343
rect -8674 4275 -8608 4309
rect -8674 4241 -8658 4275
rect -8624 4241 -8608 4275
rect -8674 4207 -8608 4241
rect -8674 4173 -8658 4207
rect -8624 4173 -8608 4207
rect -8674 4139 -8608 4173
rect -8674 4105 -8658 4139
rect -8624 4105 -8608 4139
rect -8674 4071 -8608 4105
rect -8674 4037 -8658 4071
rect -8624 4037 -8608 4071
rect -8674 4003 -8608 4037
rect -8674 3969 -8658 4003
rect -8624 3969 -8608 4003
rect -8674 3935 -8608 3969
rect -8674 3901 -8658 3935
rect -8624 3901 -8608 3935
rect -8674 3867 -8608 3901
rect -8674 3833 -8658 3867
rect -8624 3833 -8608 3867
rect -8674 3799 -8608 3833
rect -8674 3765 -8658 3799
rect -8624 3765 -8608 3799
rect -8674 3731 -8608 3765
rect -8674 3697 -8658 3731
rect -8624 3697 -8608 3731
rect -8674 3663 -8608 3697
rect -8674 3629 -8658 3663
rect -8624 3629 -8608 3663
rect -8674 3595 -8608 3629
rect -8674 3561 -8658 3595
rect -8624 3561 -8608 3595
rect -8674 3527 -8608 3561
rect -8674 3493 -8658 3527
rect -8624 3493 -8608 3527
rect -8674 3452 -8608 3493
rect -8578 4411 -8512 4452
rect -8578 4377 -8562 4411
rect -8528 4377 -8512 4411
rect -8578 4343 -8512 4377
rect -8578 4309 -8562 4343
rect -8528 4309 -8512 4343
rect -8578 4275 -8512 4309
rect -8578 4241 -8562 4275
rect -8528 4241 -8512 4275
rect -8578 4207 -8512 4241
rect -8578 4173 -8562 4207
rect -8528 4173 -8512 4207
rect -8578 4139 -8512 4173
rect -8578 4105 -8562 4139
rect -8528 4105 -8512 4139
rect -8578 4071 -8512 4105
rect -8578 4037 -8562 4071
rect -8528 4037 -8512 4071
rect -8578 4003 -8512 4037
rect -8578 3969 -8562 4003
rect -8528 3969 -8512 4003
rect -8578 3935 -8512 3969
rect -8578 3901 -8562 3935
rect -8528 3901 -8512 3935
rect -8578 3867 -8512 3901
rect -8578 3833 -8562 3867
rect -8528 3833 -8512 3867
rect -8578 3799 -8512 3833
rect -8578 3765 -8562 3799
rect -8528 3765 -8512 3799
rect -8578 3731 -8512 3765
rect -8578 3697 -8562 3731
rect -8528 3697 -8512 3731
rect -8578 3663 -8512 3697
rect -8578 3629 -8562 3663
rect -8528 3629 -8512 3663
rect -8578 3595 -8512 3629
rect -8578 3561 -8562 3595
rect -8528 3561 -8512 3595
rect -8578 3527 -8512 3561
rect -8578 3493 -8562 3527
rect -8528 3493 -8512 3527
rect -8578 3452 -8512 3493
rect -8482 4411 -8416 4452
rect -8482 4377 -8466 4411
rect -8432 4377 -8416 4411
rect -8482 4343 -8416 4377
rect -8482 4309 -8466 4343
rect -8432 4309 -8416 4343
rect -8482 4275 -8416 4309
rect -8482 4241 -8466 4275
rect -8432 4241 -8416 4275
rect -8482 4207 -8416 4241
rect -8482 4173 -8466 4207
rect -8432 4173 -8416 4207
rect -8482 4139 -8416 4173
rect -8482 4105 -8466 4139
rect -8432 4105 -8416 4139
rect -8482 4071 -8416 4105
rect -8482 4037 -8466 4071
rect -8432 4037 -8416 4071
rect -8482 4003 -8416 4037
rect -8482 3969 -8466 4003
rect -8432 3969 -8416 4003
rect -8482 3935 -8416 3969
rect -8482 3901 -8466 3935
rect -8432 3901 -8416 3935
rect -8482 3867 -8416 3901
rect -8482 3833 -8466 3867
rect -8432 3833 -8416 3867
rect -8482 3799 -8416 3833
rect -8482 3765 -8466 3799
rect -8432 3765 -8416 3799
rect -8482 3731 -8416 3765
rect -8482 3697 -8466 3731
rect -8432 3697 -8416 3731
rect -8482 3663 -8416 3697
rect -8482 3629 -8466 3663
rect -8432 3629 -8416 3663
rect -8482 3595 -8416 3629
rect -8482 3561 -8466 3595
rect -8432 3561 -8416 3595
rect -8482 3527 -8416 3561
rect -8482 3493 -8466 3527
rect -8432 3493 -8416 3527
rect -8482 3452 -8416 3493
rect -8386 4411 -8324 4452
rect -8386 4377 -8370 4411
rect -8336 4377 -8324 4411
rect -8386 4343 -8324 4377
rect -8386 4309 -8370 4343
rect -8336 4309 -8324 4343
rect -8386 4275 -8324 4309
rect -8386 4241 -8370 4275
rect -8336 4241 -8324 4275
rect -8386 4207 -8324 4241
rect -8386 4173 -8370 4207
rect -8336 4173 -8324 4207
rect -8386 4139 -8324 4173
rect -8386 4105 -8370 4139
rect -8336 4105 -8324 4139
rect -8386 4071 -8324 4105
rect -8386 4037 -8370 4071
rect -8336 4037 -8324 4071
rect -8386 4003 -8324 4037
rect -8386 3969 -8370 4003
rect -8336 3969 -8324 4003
rect -8386 3935 -8324 3969
rect -8386 3901 -8370 3935
rect -8336 3901 -8324 3935
rect -8386 3867 -8324 3901
rect -8386 3833 -8370 3867
rect -8336 3833 -8324 3867
rect -8386 3799 -8324 3833
rect -8386 3765 -8370 3799
rect -8336 3765 -8324 3799
rect -8386 3731 -8324 3765
rect -8386 3697 -8370 3731
rect -8336 3697 -8324 3731
rect -8386 3663 -8324 3697
rect -8386 3629 -8370 3663
rect -8336 3629 -8324 3663
rect -8386 3595 -8324 3629
rect -8386 3561 -8370 3595
rect -8336 3561 -8324 3595
rect -8386 3527 -8324 3561
rect -8386 3493 -8370 3527
rect -8336 3493 -8324 3527
rect -8386 3452 -8324 3493
rect -8158 4417 -8096 4458
rect -8158 4383 -8146 4417
rect -8112 4383 -8096 4417
rect -8158 4349 -8096 4383
rect -8158 4315 -8146 4349
rect -8112 4315 -8096 4349
rect -8158 4281 -8096 4315
rect -8158 4247 -8146 4281
rect -8112 4247 -8096 4281
rect -8158 4213 -8096 4247
rect -8158 4179 -8146 4213
rect -8112 4179 -8096 4213
rect -8158 4145 -8096 4179
rect -8158 4111 -8146 4145
rect -8112 4111 -8096 4145
rect -8158 4077 -8096 4111
rect -8158 4043 -8146 4077
rect -8112 4043 -8096 4077
rect -8158 4009 -8096 4043
rect -8158 3975 -8146 4009
rect -8112 3975 -8096 4009
rect -8158 3941 -8096 3975
rect -8158 3907 -8146 3941
rect -8112 3907 -8096 3941
rect -8158 3873 -8096 3907
rect -8158 3839 -8146 3873
rect -8112 3839 -8096 3873
rect -8158 3805 -8096 3839
rect -8158 3771 -8146 3805
rect -8112 3771 -8096 3805
rect -8158 3737 -8096 3771
rect -8158 3703 -8146 3737
rect -8112 3703 -8096 3737
rect -8158 3669 -8096 3703
rect -8158 3635 -8146 3669
rect -8112 3635 -8096 3669
rect -8158 3601 -8096 3635
rect -8158 3567 -8146 3601
rect -8112 3567 -8096 3601
rect -8158 3533 -8096 3567
rect -8158 3499 -8146 3533
rect -8112 3499 -8096 3533
rect -8158 3458 -8096 3499
rect -8066 4417 -8000 4458
rect -8066 4383 -8050 4417
rect -8016 4383 -8000 4417
rect -8066 4349 -8000 4383
rect -8066 4315 -8050 4349
rect -8016 4315 -8000 4349
rect -8066 4281 -8000 4315
rect -8066 4247 -8050 4281
rect -8016 4247 -8000 4281
rect -8066 4213 -8000 4247
rect -8066 4179 -8050 4213
rect -8016 4179 -8000 4213
rect -8066 4145 -8000 4179
rect -8066 4111 -8050 4145
rect -8016 4111 -8000 4145
rect -8066 4077 -8000 4111
rect -8066 4043 -8050 4077
rect -8016 4043 -8000 4077
rect -8066 4009 -8000 4043
rect -8066 3975 -8050 4009
rect -8016 3975 -8000 4009
rect -8066 3941 -8000 3975
rect -8066 3907 -8050 3941
rect -8016 3907 -8000 3941
rect -8066 3873 -8000 3907
rect -8066 3839 -8050 3873
rect -8016 3839 -8000 3873
rect -8066 3805 -8000 3839
rect -8066 3771 -8050 3805
rect -8016 3771 -8000 3805
rect -8066 3737 -8000 3771
rect -8066 3703 -8050 3737
rect -8016 3703 -8000 3737
rect -8066 3669 -8000 3703
rect -8066 3635 -8050 3669
rect -8016 3635 -8000 3669
rect -8066 3601 -8000 3635
rect -8066 3567 -8050 3601
rect -8016 3567 -8000 3601
rect -8066 3533 -8000 3567
rect -8066 3499 -8050 3533
rect -8016 3499 -8000 3533
rect -8066 3458 -8000 3499
rect -7970 4417 -7904 4458
rect -7970 4383 -7954 4417
rect -7920 4383 -7904 4417
rect -7970 4349 -7904 4383
rect -7970 4315 -7954 4349
rect -7920 4315 -7904 4349
rect -7970 4281 -7904 4315
rect -7970 4247 -7954 4281
rect -7920 4247 -7904 4281
rect -7970 4213 -7904 4247
rect -7970 4179 -7954 4213
rect -7920 4179 -7904 4213
rect -7970 4145 -7904 4179
rect -7970 4111 -7954 4145
rect -7920 4111 -7904 4145
rect -7970 4077 -7904 4111
rect -7970 4043 -7954 4077
rect -7920 4043 -7904 4077
rect -7970 4009 -7904 4043
rect -7970 3975 -7954 4009
rect -7920 3975 -7904 4009
rect -7970 3941 -7904 3975
rect -7970 3907 -7954 3941
rect -7920 3907 -7904 3941
rect -7970 3873 -7904 3907
rect -7970 3839 -7954 3873
rect -7920 3839 -7904 3873
rect -7970 3805 -7904 3839
rect -7970 3771 -7954 3805
rect -7920 3771 -7904 3805
rect -7970 3737 -7904 3771
rect -7970 3703 -7954 3737
rect -7920 3703 -7904 3737
rect -7970 3669 -7904 3703
rect -7970 3635 -7954 3669
rect -7920 3635 -7904 3669
rect -7970 3601 -7904 3635
rect -7970 3567 -7954 3601
rect -7920 3567 -7904 3601
rect -7970 3533 -7904 3567
rect -7970 3499 -7954 3533
rect -7920 3499 -7904 3533
rect -7970 3458 -7904 3499
rect -7874 4417 -7808 4458
rect -7874 4383 -7858 4417
rect -7824 4383 -7808 4417
rect -7874 4349 -7808 4383
rect -7874 4315 -7858 4349
rect -7824 4315 -7808 4349
rect -7874 4281 -7808 4315
rect -7874 4247 -7858 4281
rect -7824 4247 -7808 4281
rect -7874 4213 -7808 4247
rect -7874 4179 -7858 4213
rect -7824 4179 -7808 4213
rect -7874 4145 -7808 4179
rect -7874 4111 -7858 4145
rect -7824 4111 -7808 4145
rect -7874 4077 -7808 4111
rect -7874 4043 -7858 4077
rect -7824 4043 -7808 4077
rect -7874 4009 -7808 4043
rect -7874 3975 -7858 4009
rect -7824 3975 -7808 4009
rect -7874 3941 -7808 3975
rect -7874 3907 -7858 3941
rect -7824 3907 -7808 3941
rect -7874 3873 -7808 3907
rect -7874 3839 -7858 3873
rect -7824 3839 -7808 3873
rect -7874 3805 -7808 3839
rect -7874 3771 -7858 3805
rect -7824 3771 -7808 3805
rect -7874 3737 -7808 3771
rect -7874 3703 -7858 3737
rect -7824 3703 -7808 3737
rect -7874 3669 -7808 3703
rect -7874 3635 -7858 3669
rect -7824 3635 -7808 3669
rect -7874 3601 -7808 3635
rect -7874 3567 -7858 3601
rect -7824 3567 -7808 3601
rect -7874 3533 -7808 3567
rect -7874 3499 -7858 3533
rect -7824 3499 -7808 3533
rect -7874 3458 -7808 3499
rect -7778 4417 -7712 4458
rect -7778 4383 -7762 4417
rect -7728 4383 -7712 4417
rect -7778 4349 -7712 4383
rect -7778 4315 -7762 4349
rect -7728 4315 -7712 4349
rect -7778 4281 -7712 4315
rect -7778 4247 -7762 4281
rect -7728 4247 -7712 4281
rect -7778 4213 -7712 4247
rect -7778 4179 -7762 4213
rect -7728 4179 -7712 4213
rect -7778 4145 -7712 4179
rect -7778 4111 -7762 4145
rect -7728 4111 -7712 4145
rect -7778 4077 -7712 4111
rect -7778 4043 -7762 4077
rect -7728 4043 -7712 4077
rect -7778 4009 -7712 4043
rect -7778 3975 -7762 4009
rect -7728 3975 -7712 4009
rect -7778 3941 -7712 3975
rect -7778 3907 -7762 3941
rect -7728 3907 -7712 3941
rect -7778 3873 -7712 3907
rect -7778 3839 -7762 3873
rect -7728 3839 -7712 3873
rect -7778 3805 -7712 3839
rect -7778 3771 -7762 3805
rect -7728 3771 -7712 3805
rect -7778 3737 -7712 3771
rect -7778 3703 -7762 3737
rect -7728 3703 -7712 3737
rect -7778 3669 -7712 3703
rect -7778 3635 -7762 3669
rect -7728 3635 -7712 3669
rect -7778 3601 -7712 3635
rect -7778 3567 -7762 3601
rect -7728 3567 -7712 3601
rect -7778 3533 -7712 3567
rect -7778 3499 -7762 3533
rect -7728 3499 -7712 3533
rect -7778 3458 -7712 3499
rect -7682 4417 -7616 4458
rect -7682 4383 -7666 4417
rect -7632 4383 -7616 4417
rect -7682 4349 -7616 4383
rect -7682 4315 -7666 4349
rect -7632 4315 -7616 4349
rect -7682 4281 -7616 4315
rect -7682 4247 -7666 4281
rect -7632 4247 -7616 4281
rect -7682 4213 -7616 4247
rect -7682 4179 -7666 4213
rect -7632 4179 -7616 4213
rect -7682 4145 -7616 4179
rect -7682 4111 -7666 4145
rect -7632 4111 -7616 4145
rect -7682 4077 -7616 4111
rect -7682 4043 -7666 4077
rect -7632 4043 -7616 4077
rect -7682 4009 -7616 4043
rect -7682 3975 -7666 4009
rect -7632 3975 -7616 4009
rect -7682 3941 -7616 3975
rect -7682 3907 -7666 3941
rect -7632 3907 -7616 3941
rect -7682 3873 -7616 3907
rect -7682 3839 -7666 3873
rect -7632 3839 -7616 3873
rect -7682 3805 -7616 3839
rect -7682 3771 -7666 3805
rect -7632 3771 -7616 3805
rect -7682 3737 -7616 3771
rect -7682 3703 -7666 3737
rect -7632 3703 -7616 3737
rect -7682 3669 -7616 3703
rect -7682 3635 -7666 3669
rect -7632 3635 -7616 3669
rect -7682 3601 -7616 3635
rect -7682 3567 -7666 3601
rect -7632 3567 -7616 3601
rect -7682 3533 -7616 3567
rect -7682 3499 -7666 3533
rect -7632 3499 -7616 3533
rect -7682 3458 -7616 3499
rect -7586 4417 -7520 4458
rect -7586 4383 -7570 4417
rect -7536 4383 -7520 4417
rect -7586 4349 -7520 4383
rect -7586 4315 -7570 4349
rect -7536 4315 -7520 4349
rect -7586 4281 -7520 4315
rect -7586 4247 -7570 4281
rect -7536 4247 -7520 4281
rect -7586 4213 -7520 4247
rect -7586 4179 -7570 4213
rect -7536 4179 -7520 4213
rect -7586 4145 -7520 4179
rect -7586 4111 -7570 4145
rect -7536 4111 -7520 4145
rect -7586 4077 -7520 4111
rect -7586 4043 -7570 4077
rect -7536 4043 -7520 4077
rect -7586 4009 -7520 4043
rect -7586 3975 -7570 4009
rect -7536 3975 -7520 4009
rect -7586 3941 -7520 3975
rect -7586 3907 -7570 3941
rect -7536 3907 -7520 3941
rect -7586 3873 -7520 3907
rect -7586 3839 -7570 3873
rect -7536 3839 -7520 3873
rect -7586 3805 -7520 3839
rect -7586 3771 -7570 3805
rect -7536 3771 -7520 3805
rect -7586 3737 -7520 3771
rect -7586 3703 -7570 3737
rect -7536 3703 -7520 3737
rect -7586 3669 -7520 3703
rect -7586 3635 -7570 3669
rect -7536 3635 -7520 3669
rect -7586 3601 -7520 3635
rect -7586 3567 -7570 3601
rect -7536 3567 -7520 3601
rect -7586 3533 -7520 3567
rect -7586 3499 -7570 3533
rect -7536 3499 -7520 3533
rect -7586 3458 -7520 3499
rect -7490 4417 -7424 4458
rect -7490 4383 -7474 4417
rect -7440 4383 -7424 4417
rect -7490 4349 -7424 4383
rect -7490 4315 -7474 4349
rect -7440 4315 -7424 4349
rect -7490 4281 -7424 4315
rect -7490 4247 -7474 4281
rect -7440 4247 -7424 4281
rect -7490 4213 -7424 4247
rect -7490 4179 -7474 4213
rect -7440 4179 -7424 4213
rect -7490 4145 -7424 4179
rect -7490 4111 -7474 4145
rect -7440 4111 -7424 4145
rect -7490 4077 -7424 4111
rect -7490 4043 -7474 4077
rect -7440 4043 -7424 4077
rect -7490 4009 -7424 4043
rect -7490 3975 -7474 4009
rect -7440 3975 -7424 4009
rect -7490 3941 -7424 3975
rect -7490 3907 -7474 3941
rect -7440 3907 -7424 3941
rect -7490 3873 -7424 3907
rect -7490 3839 -7474 3873
rect -7440 3839 -7424 3873
rect -7490 3805 -7424 3839
rect -7490 3771 -7474 3805
rect -7440 3771 -7424 3805
rect -7490 3737 -7424 3771
rect -7490 3703 -7474 3737
rect -7440 3703 -7424 3737
rect -7490 3669 -7424 3703
rect -7490 3635 -7474 3669
rect -7440 3635 -7424 3669
rect -7490 3601 -7424 3635
rect -7490 3567 -7474 3601
rect -7440 3567 -7424 3601
rect -7490 3533 -7424 3567
rect -7490 3499 -7474 3533
rect -7440 3499 -7424 3533
rect -7490 3458 -7424 3499
rect -7394 4417 -7328 4458
rect -7394 4383 -7378 4417
rect -7344 4383 -7328 4417
rect -7394 4349 -7328 4383
rect -7394 4315 -7378 4349
rect -7344 4315 -7328 4349
rect -7394 4281 -7328 4315
rect -7394 4247 -7378 4281
rect -7344 4247 -7328 4281
rect -7394 4213 -7328 4247
rect -7394 4179 -7378 4213
rect -7344 4179 -7328 4213
rect -7394 4145 -7328 4179
rect -7394 4111 -7378 4145
rect -7344 4111 -7328 4145
rect -7394 4077 -7328 4111
rect -7394 4043 -7378 4077
rect -7344 4043 -7328 4077
rect -7394 4009 -7328 4043
rect -7394 3975 -7378 4009
rect -7344 3975 -7328 4009
rect -7394 3941 -7328 3975
rect -7394 3907 -7378 3941
rect -7344 3907 -7328 3941
rect -7394 3873 -7328 3907
rect -7394 3839 -7378 3873
rect -7344 3839 -7328 3873
rect -7394 3805 -7328 3839
rect -7394 3771 -7378 3805
rect -7344 3771 -7328 3805
rect -7394 3737 -7328 3771
rect -7394 3703 -7378 3737
rect -7344 3703 -7328 3737
rect -7394 3669 -7328 3703
rect -7394 3635 -7378 3669
rect -7344 3635 -7328 3669
rect -7394 3601 -7328 3635
rect -7394 3567 -7378 3601
rect -7344 3567 -7328 3601
rect -7394 3533 -7328 3567
rect -7394 3499 -7378 3533
rect -7344 3499 -7328 3533
rect -7394 3458 -7328 3499
rect -7298 4417 -7232 4458
rect -7298 4383 -7282 4417
rect -7248 4383 -7232 4417
rect -7298 4349 -7232 4383
rect -7298 4315 -7282 4349
rect -7248 4315 -7232 4349
rect -7298 4281 -7232 4315
rect -7298 4247 -7282 4281
rect -7248 4247 -7232 4281
rect -7298 4213 -7232 4247
rect -7298 4179 -7282 4213
rect -7248 4179 -7232 4213
rect -7298 4145 -7232 4179
rect -7298 4111 -7282 4145
rect -7248 4111 -7232 4145
rect -7298 4077 -7232 4111
rect -7298 4043 -7282 4077
rect -7248 4043 -7232 4077
rect -7298 4009 -7232 4043
rect -7298 3975 -7282 4009
rect -7248 3975 -7232 4009
rect -7298 3941 -7232 3975
rect -7298 3907 -7282 3941
rect -7248 3907 -7232 3941
rect -7298 3873 -7232 3907
rect -7298 3839 -7282 3873
rect -7248 3839 -7232 3873
rect -7298 3805 -7232 3839
rect -7298 3771 -7282 3805
rect -7248 3771 -7232 3805
rect -7298 3737 -7232 3771
rect -7298 3703 -7282 3737
rect -7248 3703 -7232 3737
rect -7298 3669 -7232 3703
rect -7298 3635 -7282 3669
rect -7248 3635 -7232 3669
rect -7298 3601 -7232 3635
rect -7298 3567 -7282 3601
rect -7248 3567 -7232 3601
rect -7298 3533 -7232 3567
rect -7298 3499 -7282 3533
rect -7248 3499 -7232 3533
rect -7298 3458 -7232 3499
rect -7202 4417 -7136 4458
rect -7202 4383 -7186 4417
rect -7152 4383 -7136 4417
rect -7202 4349 -7136 4383
rect -7202 4315 -7186 4349
rect -7152 4315 -7136 4349
rect -7202 4281 -7136 4315
rect -7202 4247 -7186 4281
rect -7152 4247 -7136 4281
rect -7202 4213 -7136 4247
rect -7202 4179 -7186 4213
rect -7152 4179 -7136 4213
rect -7202 4145 -7136 4179
rect -7202 4111 -7186 4145
rect -7152 4111 -7136 4145
rect -7202 4077 -7136 4111
rect -7202 4043 -7186 4077
rect -7152 4043 -7136 4077
rect -7202 4009 -7136 4043
rect -7202 3975 -7186 4009
rect -7152 3975 -7136 4009
rect -7202 3941 -7136 3975
rect -7202 3907 -7186 3941
rect -7152 3907 -7136 3941
rect -7202 3873 -7136 3907
rect -7202 3839 -7186 3873
rect -7152 3839 -7136 3873
rect -7202 3805 -7136 3839
rect -7202 3771 -7186 3805
rect -7152 3771 -7136 3805
rect -7202 3737 -7136 3771
rect -7202 3703 -7186 3737
rect -7152 3703 -7136 3737
rect -7202 3669 -7136 3703
rect -7202 3635 -7186 3669
rect -7152 3635 -7136 3669
rect -7202 3601 -7136 3635
rect -7202 3567 -7186 3601
rect -7152 3567 -7136 3601
rect -7202 3533 -7136 3567
rect -7202 3499 -7186 3533
rect -7152 3499 -7136 3533
rect -7202 3458 -7136 3499
rect -7106 4417 -7040 4458
rect -7106 4383 -7090 4417
rect -7056 4383 -7040 4417
rect -7106 4349 -7040 4383
rect -7106 4315 -7090 4349
rect -7056 4315 -7040 4349
rect -7106 4281 -7040 4315
rect -7106 4247 -7090 4281
rect -7056 4247 -7040 4281
rect -7106 4213 -7040 4247
rect -7106 4179 -7090 4213
rect -7056 4179 -7040 4213
rect -7106 4145 -7040 4179
rect -7106 4111 -7090 4145
rect -7056 4111 -7040 4145
rect -7106 4077 -7040 4111
rect -7106 4043 -7090 4077
rect -7056 4043 -7040 4077
rect -7106 4009 -7040 4043
rect -7106 3975 -7090 4009
rect -7056 3975 -7040 4009
rect -7106 3941 -7040 3975
rect -7106 3907 -7090 3941
rect -7056 3907 -7040 3941
rect -7106 3873 -7040 3907
rect -7106 3839 -7090 3873
rect -7056 3839 -7040 3873
rect -7106 3805 -7040 3839
rect -7106 3771 -7090 3805
rect -7056 3771 -7040 3805
rect -7106 3737 -7040 3771
rect -7106 3703 -7090 3737
rect -7056 3703 -7040 3737
rect -7106 3669 -7040 3703
rect -7106 3635 -7090 3669
rect -7056 3635 -7040 3669
rect -7106 3601 -7040 3635
rect -7106 3567 -7090 3601
rect -7056 3567 -7040 3601
rect -7106 3533 -7040 3567
rect -7106 3499 -7090 3533
rect -7056 3499 -7040 3533
rect -7106 3458 -7040 3499
rect -7010 4417 -6944 4458
rect -7010 4383 -6994 4417
rect -6960 4383 -6944 4417
rect -7010 4349 -6944 4383
rect -7010 4315 -6994 4349
rect -6960 4315 -6944 4349
rect -7010 4281 -6944 4315
rect -7010 4247 -6994 4281
rect -6960 4247 -6944 4281
rect -7010 4213 -6944 4247
rect -7010 4179 -6994 4213
rect -6960 4179 -6944 4213
rect -7010 4145 -6944 4179
rect -7010 4111 -6994 4145
rect -6960 4111 -6944 4145
rect -7010 4077 -6944 4111
rect -7010 4043 -6994 4077
rect -6960 4043 -6944 4077
rect -7010 4009 -6944 4043
rect -7010 3975 -6994 4009
rect -6960 3975 -6944 4009
rect -7010 3941 -6944 3975
rect -7010 3907 -6994 3941
rect -6960 3907 -6944 3941
rect -7010 3873 -6944 3907
rect -7010 3839 -6994 3873
rect -6960 3839 -6944 3873
rect -7010 3805 -6944 3839
rect -7010 3771 -6994 3805
rect -6960 3771 -6944 3805
rect -7010 3737 -6944 3771
rect -7010 3703 -6994 3737
rect -6960 3703 -6944 3737
rect -7010 3669 -6944 3703
rect -7010 3635 -6994 3669
rect -6960 3635 -6944 3669
rect -7010 3601 -6944 3635
rect -7010 3567 -6994 3601
rect -6960 3567 -6944 3601
rect -7010 3533 -6944 3567
rect -7010 3499 -6994 3533
rect -6960 3499 -6944 3533
rect -7010 3458 -6944 3499
rect -6914 4417 -6848 4458
rect -6914 4383 -6898 4417
rect -6864 4383 -6848 4417
rect -6914 4349 -6848 4383
rect -6914 4315 -6898 4349
rect -6864 4315 -6848 4349
rect -6914 4281 -6848 4315
rect -6914 4247 -6898 4281
rect -6864 4247 -6848 4281
rect -6914 4213 -6848 4247
rect -6914 4179 -6898 4213
rect -6864 4179 -6848 4213
rect -6914 4145 -6848 4179
rect -6914 4111 -6898 4145
rect -6864 4111 -6848 4145
rect -6914 4077 -6848 4111
rect -6914 4043 -6898 4077
rect -6864 4043 -6848 4077
rect -6914 4009 -6848 4043
rect -6914 3975 -6898 4009
rect -6864 3975 -6848 4009
rect -6914 3941 -6848 3975
rect -6914 3907 -6898 3941
rect -6864 3907 -6848 3941
rect -6914 3873 -6848 3907
rect -6914 3839 -6898 3873
rect -6864 3839 -6848 3873
rect -6914 3805 -6848 3839
rect -6914 3771 -6898 3805
rect -6864 3771 -6848 3805
rect -6914 3737 -6848 3771
rect -6914 3703 -6898 3737
rect -6864 3703 -6848 3737
rect -6914 3669 -6848 3703
rect -6914 3635 -6898 3669
rect -6864 3635 -6848 3669
rect -6914 3601 -6848 3635
rect -6914 3567 -6898 3601
rect -6864 3567 -6848 3601
rect -6914 3533 -6848 3567
rect -6914 3499 -6898 3533
rect -6864 3499 -6848 3533
rect -6914 3458 -6848 3499
rect -6818 4417 -6752 4458
rect -6818 4383 -6802 4417
rect -6768 4383 -6752 4417
rect -6818 4349 -6752 4383
rect -6818 4315 -6802 4349
rect -6768 4315 -6752 4349
rect -6818 4281 -6752 4315
rect -6818 4247 -6802 4281
rect -6768 4247 -6752 4281
rect -6818 4213 -6752 4247
rect -6818 4179 -6802 4213
rect -6768 4179 -6752 4213
rect -6818 4145 -6752 4179
rect -6818 4111 -6802 4145
rect -6768 4111 -6752 4145
rect -6818 4077 -6752 4111
rect -6818 4043 -6802 4077
rect -6768 4043 -6752 4077
rect -6818 4009 -6752 4043
rect -6818 3975 -6802 4009
rect -6768 3975 -6752 4009
rect -6818 3941 -6752 3975
rect -6818 3907 -6802 3941
rect -6768 3907 -6752 3941
rect -6818 3873 -6752 3907
rect -6818 3839 -6802 3873
rect -6768 3839 -6752 3873
rect -6818 3805 -6752 3839
rect -6818 3771 -6802 3805
rect -6768 3771 -6752 3805
rect -6818 3737 -6752 3771
rect -6818 3703 -6802 3737
rect -6768 3703 -6752 3737
rect -6818 3669 -6752 3703
rect -6818 3635 -6802 3669
rect -6768 3635 -6752 3669
rect -6818 3601 -6752 3635
rect -6818 3567 -6802 3601
rect -6768 3567 -6752 3601
rect -6818 3533 -6752 3567
rect -6818 3499 -6802 3533
rect -6768 3499 -6752 3533
rect -6818 3458 -6752 3499
rect -6722 4417 -6660 4458
rect -6722 4383 -6706 4417
rect -6672 4383 -6660 4417
rect -6722 4349 -6660 4383
rect -6722 4315 -6706 4349
rect -6672 4315 -6660 4349
rect -6722 4281 -6660 4315
rect -6722 4247 -6706 4281
rect -6672 4247 -6660 4281
rect -6722 4213 -6660 4247
rect -6722 4179 -6706 4213
rect -6672 4179 -6660 4213
rect -6722 4145 -6660 4179
rect -6722 4111 -6706 4145
rect -6672 4111 -6660 4145
rect -6722 4077 -6660 4111
rect -6722 4043 -6706 4077
rect -6672 4043 -6660 4077
rect -6722 4009 -6660 4043
rect -6722 3975 -6706 4009
rect -6672 3975 -6660 4009
rect -6722 3941 -6660 3975
rect -6722 3907 -6706 3941
rect -6672 3907 -6660 3941
rect -6722 3873 -6660 3907
rect -6722 3839 -6706 3873
rect -6672 3839 -6660 3873
rect -6722 3805 -6660 3839
rect -6722 3771 -6706 3805
rect -6672 3771 -6660 3805
rect -6722 3737 -6660 3771
rect -6722 3703 -6706 3737
rect -6672 3703 -6660 3737
rect -6722 3669 -6660 3703
rect -6722 3635 -6706 3669
rect -6672 3635 -6660 3669
rect -6722 3601 -6660 3635
rect -6722 3567 -6706 3601
rect -6672 3567 -6660 3601
rect -6722 3533 -6660 3567
rect -6722 3499 -6706 3533
rect -6672 3499 -6660 3533
rect -6722 3458 -6660 3499
rect -6474 4423 -6412 4464
rect -6474 4389 -6462 4423
rect -6428 4389 -6412 4423
rect -6474 4355 -6412 4389
rect -6474 4321 -6462 4355
rect -6428 4321 -6412 4355
rect -6474 4287 -6412 4321
rect -6474 4253 -6462 4287
rect -6428 4253 -6412 4287
rect -6474 4219 -6412 4253
rect -6474 4185 -6462 4219
rect -6428 4185 -6412 4219
rect -6474 4151 -6412 4185
rect -6474 4117 -6462 4151
rect -6428 4117 -6412 4151
rect -6474 4083 -6412 4117
rect -6474 4049 -6462 4083
rect -6428 4049 -6412 4083
rect -6474 4015 -6412 4049
rect -6474 3981 -6462 4015
rect -6428 3981 -6412 4015
rect -6474 3947 -6412 3981
rect -6474 3913 -6462 3947
rect -6428 3913 -6412 3947
rect -6474 3879 -6412 3913
rect -6474 3845 -6462 3879
rect -6428 3845 -6412 3879
rect -6474 3811 -6412 3845
rect -6474 3777 -6462 3811
rect -6428 3777 -6412 3811
rect -6474 3743 -6412 3777
rect -6474 3709 -6462 3743
rect -6428 3709 -6412 3743
rect -6474 3675 -6412 3709
rect -6474 3641 -6462 3675
rect -6428 3641 -6412 3675
rect -6474 3607 -6412 3641
rect -6474 3573 -6462 3607
rect -6428 3573 -6412 3607
rect -6474 3539 -6412 3573
rect -6474 3505 -6462 3539
rect -6428 3505 -6412 3539
rect -6474 3464 -6412 3505
rect -6382 4423 -6316 4464
rect -6382 4389 -6366 4423
rect -6332 4389 -6316 4423
rect -6382 4355 -6316 4389
rect -6382 4321 -6366 4355
rect -6332 4321 -6316 4355
rect -6382 4287 -6316 4321
rect -6382 4253 -6366 4287
rect -6332 4253 -6316 4287
rect -6382 4219 -6316 4253
rect -6382 4185 -6366 4219
rect -6332 4185 -6316 4219
rect -6382 4151 -6316 4185
rect -6382 4117 -6366 4151
rect -6332 4117 -6316 4151
rect -6382 4083 -6316 4117
rect -6382 4049 -6366 4083
rect -6332 4049 -6316 4083
rect -6382 4015 -6316 4049
rect -6382 3981 -6366 4015
rect -6332 3981 -6316 4015
rect -6382 3947 -6316 3981
rect -6382 3913 -6366 3947
rect -6332 3913 -6316 3947
rect -6382 3879 -6316 3913
rect -6382 3845 -6366 3879
rect -6332 3845 -6316 3879
rect -6382 3811 -6316 3845
rect -6382 3777 -6366 3811
rect -6332 3777 -6316 3811
rect -6382 3743 -6316 3777
rect -6382 3709 -6366 3743
rect -6332 3709 -6316 3743
rect -6382 3675 -6316 3709
rect -6382 3641 -6366 3675
rect -6332 3641 -6316 3675
rect -6382 3607 -6316 3641
rect -6382 3573 -6366 3607
rect -6332 3573 -6316 3607
rect -6382 3539 -6316 3573
rect -6382 3505 -6366 3539
rect -6332 3505 -6316 3539
rect -6382 3464 -6316 3505
rect -6286 4423 -6220 4464
rect -6286 4389 -6270 4423
rect -6236 4389 -6220 4423
rect -6286 4355 -6220 4389
rect -6286 4321 -6270 4355
rect -6236 4321 -6220 4355
rect -6286 4287 -6220 4321
rect -6286 4253 -6270 4287
rect -6236 4253 -6220 4287
rect -6286 4219 -6220 4253
rect -6286 4185 -6270 4219
rect -6236 4185 -6220 4219
rect -6286 4151 -6220 4185
rect -6286 4117 -6270 4151
rect -6236 4117 -6220 4151
rect -6286 4083 -6220 4117
rect -6286 4049 -6270 4083
rect -6236 4049 -6220 4083
rect -6286 4015 -6220 4049
rect -6286 3981 -6270 4015
rect -6236 3981 -6220 4015
rect -6286 3947 -6220 3981
rect -6286 3913 -6270 3947
rect -6236 3913 -6220 3947
rect -6286 3879 -6220 3913
rect -6286 3845 -6270 3879
rect -6236 3845 -6220 3879
rect -6286 3811 -6220 3845
rect -6286 3777 -6270 3811
rect -6236 3777 -6220 3811
rect -6286 3743 -6220 3777
rect -6286 3709 -6270 3743
rect -6236 3709 -6220 3743
rect -6286 3675 -6220 3709
rect -6286 3641 -6270 3675
rect -6236 3641 -6220 3675
rect -6286 3607 -6220 3641
rect -6286 3573 -6270 3607
rect -6236 3573 -6220 3607
rect -6286 3539 -6220 3573
rect -6286 3505 -6270 3539
rect -6236 3505 -6220 3539
rect -6286 3464 -6220 3505
rect -6190 4423 -6124 4464
rect -6190 4389 -6174 4423
rect -6140 4389 -6124 4423
rect -6190 4355 -6124 4389
rect -6190 4321 -6174 4355
rect -6140 4321 -6124 4355
rect -6190 4287 -6124 4321
rect -6190 4253 -6174 4287
rect -6140 4253 -6124 4287
rect -6190 4219 -6124 4253
rect -6190 4185 -6174 4219
rect -6140 4185 -6124 4219
rect -6190 4151 -6124 4185
rect -6190 4117 -6174 4151
rect -6140 4117 -6124 4151
rect -6190 4083 -6124 4117
rect -6190 4049 -6174 4083
rect -6140 4049 -6124 4083
rect -6190 4015 -6124 4049
rect -6190 3981 -6174 4015
rect -6140 3981 -6124 4015
rect -6190 3947 -6124 3981
rect -6190 3913 -6174 3947
rect -6140 3913 -6124 3947
rect -6190 3879 -6124 3913
rect -6190 3845 -6174 3879
rect -6140 3845 -6124 3879
rect -6190 3811 -6124 3845
rect -6190 3777 -6174 3811
rect -6140 3777 -6124 3811
rect -6190 3743 -6124 3777
rect -6190 3709 -6174 3743
rect -6140 3709 -6124 3743
rect -6190 3675 -6124 3709
rect -6190 3641 -6174 3675
rect -6140 3641 -6124 3675
rect -6190 3607 -6124 3641
rect -6190 3573 -6174 3607
rect -6140 3573 -6124 3607
rect -6190 3539 -6124 3573
rect -6190 3505 -6174 3539
rect -6140 3505 -6124 3539
rect -6190 3464 -6124 3505
rect -6094 4423 -6028 4464
rect -6094 4389 -6078 4423
rect -6044 4389 -6028 4423
rect -6094 4355 -6028 4389
rect -6094 4321 -6078 4355
rect -6044 4321 -6028 4355
rect -6094 4287 -6028 4321
rect -6094 4253 -6078 4287
rect -6044 4253 -6028 4287
rect -6094 4219 -6028 4253
rect -6094 4185 -6078 4219
rect -6044 4185 -6028 4219
rect -6094 4151 -6028 4185
rect -6094 4117 -6078 4151
rect -6044 4117 -6028 4151
rect -6094 4083 -6028 4117
rect -6094 4049 -6078 4083
rect -6044 4049 -6028 4083
rect -6094 4015 -6028 4049
rect -6094 3981 -6078 4015
rect -6044 3981 -6028 4015
rect -6094 3947 -6028 3981
rect -6094 3913 -6078 3947
rect -6044 3913 -6028 3947
rect -6094 3879 -6028 3913
rect -6094 3845 -6078 3879
rect -6044 3845 -6028 3879
rect -6094 3811 -6028 3845
rect -6094 3777 -6078 3811
rect -6044 3777 -6028 3811
rect -6094 3743 -6028 3777
rect -6094 3709 -6078 3743
rect -6044 3709 -6028 3743
rect -6094 3675 -6028 3709
rect -6094 3641 -6078 3675
rect -6044 3641 -6028 3675
rect -6094 3607 -6028 3641
rect -6094 3573 -6078 3607
rect -6044 3573 -6028 3607
rect -6094 3539 -6028 3573
rect -6094 3505 -6078 3539
rect -6044 3505 -6028 3539
rect -6094 3464 -6028 3505
rect -5998 4423 -5932 4464
rect -5998 4389 -5982 4423
rect -5948 4389 -5932 4423
rect -5998 4355 -5932 4389
rect -5998 4321 -5982 4355
rect -5948 4321 -5932 4355
rect -5998 4287 -5932 4321
rect -5998 4253 -5982 4287
rect -5948 4253 -5932 4287
rect -5998 4219 -5932 4253
rect -5998 4185 -5982 4219
rect -5948 4185 -5932 4219
rect -5998 4151 -5932 4185
rect -5998 4117 -5982 4151
rect -5948 4117 -5932 4151
rect -5998 4083 -5932 4117
rect -5998 4049 -5982 4083
rect -5948 4049 -5932 4083
rect -5998 4015 -5932 4049
rect -5998 3981 -5982 4015
rect -5948 3981 -5932 4015
rect -5998 3947 -5932 3981
rect -5998 3913 -5982 3947
rect -5948 3913 -5932 3947
rect -5998 3879 -5932 3913
rect -5998 3845 -5982 3879
rect -5948 3845 -5932 3879
rect -5998 3811 -5932 3845
rect -5998 3777 -5982 3811
rect -5948 3777 -5932 3811
rect -5998 3743 -5932 3777
rect -5998 3709 -5982 3743
rect -5948 3709 -5932 3743
rect -5998 3675 -5932 3709
rect -5998 3641 -5982 3675
rect -5948 3641 -5932 3675
rect -5998 3607 -5932 3641
rect -5998 3573 -5982 3607
rect -5948 3573 -5932 3607
rect -5998 3539 -5932 3573
rect -5998 3505 -5982 3539
rect -5948 3505 -5932 3539
rect -5998 3464 -5932 3505
rect -5902 4423 -5836 4464
rect -5902 4389 -5886 4423
rect -5852 4389 -5836 4423
rect -5902 4355 -5836 4389
rect -5902 4321 -5886 4355
rect -5852 4321 -5836 4355
rect -5902 4287 -5836 4321
rect -5902 4253 -5886 4287
rect -5852 4253 -5836 4287
rect -5902 4219 -5836 4253
rect -5902 4185 -5886 4219
rect -5852 4185 -5836 4219
rect -5902 4151 -5836 4185
rect -5902 4117 -5886 4151
rect -5852 4117 -5836 4151
rect -5902 4083 -5836 4117
rect -5902 4049 -5886 4083
rect -5852 4049 -5836 4083
rect -5902 4015 -5836 4049
rect -5902 3981 -5886 4015
rect -5852 3981 -5836 4015
rect -5902 3947 -5836 3981
rect -5902 3913 -5886 3947
rect -5852 3913 -5836 3947
rect -5902 3879 -5836 3913
rect -5902 3845 -5886 3879
rect -5852 3845 -5836 3879
rect -5902 3811 -5836 3845
rect -5902 3777 -5886 3811
rect -5852 3777 -5836 3811
rect -5902 3743 -5836 3777
rect -5902 3709 -5886 3743
rect -5852 3709 -5836 3743
rect -5902 3675 -5836 3709
rect -5902 3641 -5886 3675
rect -5852 3641 -5836 3675
rect -5902 3607 -5836 3641
rect -5902 3573 -5886 3607
rect -5852 3573 -5836 3607
rect -5902 3539 -5836 3573
rect -5902 3505 -5886 3539
rect -5852 3505 -5836 3539
rect -5902 3464 -5836 3505
rect -5806 4423 -5740 4464
rect -5806 4389 -5790 4423
rect -5756 4389 -5740 4423
rect -5806 4355 -5740 4389
rect -5806 4321 -5790 4355
rect -5756 4321 -5740 4355
rect -5806 4287 -5740 4321
rect -5806 4253 -5790 4287
rect -5756 4253 -5740 4287
rect -5806 4219 -5740 4253
rect -5806 4185 -5790 4219
rect -5756 4185 -5740 4219
rect -5806 4151 -5740 4185
rect -5806 4117 -5790 4151
rect -5756 4117 -5740 4151
rect -5806 4083 -5740 4117
rect -5806 4049 -5790 4083
rect -5756 4049 -5740 4083
rect -5806 4015 -5740 4049
rect -5806 3981 -5790 4015
rect -5756 3981 -5740 4015
rect -5806 3947 -5740 3981
rect -5806 3913 -5790 3947
rect -5756 3913 -5740 3947
rect -5806 3879 -5740 3913
rect -5806 3845 -5790 3879
rect -5756 3845 -5740 3879
rect -5806 3811 -5740 3845
rect -5806 3777 -5790 3811
rect -5756 3777 -5740 3811
rect -5806 3743 -5740 3777
rect -5806 3709 -5790 3743
rect -5756 3709 -5740 3743
rect -5806 3675 -5740 3709
rect -5806 3641 -5790 3675
rect -5756 3641 -5740 3675
rect -5806 3607 -5740 3641
rect -5806 3573 -5790 3607
rect -5756 3573 -5740 3607
rect -5806 3539 -5740 3573
rect -5806 3505 -5790 3539
rect -5756 3505 -5740 3539
rect -5806 3464 -5740 3505
rect -5710 4423 -5644 4464
rect -5710 4389 -5694 4423
rect -5660 4389 -5644 4423
rect -5710 4355 -5644 4389
rect -5710 4321 -5694 4355
rect -5660 4321 -5644 4355
rect -5710 4287 -5644 4321
rect -5710 4253 -5694 4287
rect -5660 4253 -5644 4287
rect -5710 4219 -5644 4253
rect -5710 4185 -5694 4219
rect -5660 4185 -5644 4219
rect -5710 4151 -5644 4185
rect -5710 4117 -5694 4151
rect -5660 4117 -5644 4151
rect -5710 4083 -5644 4117
rect -5710 4049 -5694 4083
rect -5660 4049 -5644 4083
rect -5710 4015 -5644 4049
rect -5710 3981 -5694 4015
rect -5660 3981 -5644 4015
rect -5710 3947 -5644 3981
rect -5710 3913 -5694 3947
rect -5660 3913 -5644 3947
rect -5710 3879 -5644 3913
rect -5710 3845 -5694 3879
rect -5660 3845 -5644 3879
rect -5710 3811 -5644 3845
rect -5710 3777 -5694 3811
rect -5660 3777 -5644 3811
rect -5710 3743 -5644 3777
rect -5710 3709 -5694 3743
rect -5660 3709 -5644 3743
rect -5710 3675 -5644 3709
rect -5710 3641 -5694 3675
rect -5660 3641 -5644 3675
rect -5710 3607 -5644 3641
rect -5710 3573 -5694 3607
rect -5660 3573 -5644 3607
rect -5710 3539 -5644 3573
rect -5710 3505 -5694 3539
rect -5660 3505 -5644 3539
rect -5710 3464 -5644 3505
rect -5614 4423 -5548 4464
rect -5614 4389 -5598 4423
rect -5564 4389 -5548 4423
rect -5614 4355 -5548 4389
rect -5614 4321 -5598 4355
rect -5564 4321 -5548 4355
rect -5614 4287 -5548 4321
rect -5614 4253 -5598 4287
rect -5564 4253 -5548 4287
rect -5614 4219 -5548 4253
rect -5614 4185 -5598 4219
rect -5564 4185 -5548 4219
rect -5614 4151 -5548 4185
rect -5614 4117 -5598 4151
rect -5564 4117 -5548 4151
rect -5614 4083 -5548 4117
rect -5614 4049 -5598 4083
rect -5564 4049 -5548 4083
rect -5614 4015 -5548 4049
rect -5614 3981 -5598 4015
rect -5564 3981 -5548 4015
rect -5614 3947 -5548 3981
rect -5614 3913 -5598 3947
rect -5564 3913 -5548 3947
rect -5614 3879 -5548 3913
rect -5614 3845 -5598 3879
rect -5564 3845 -5548 3879
rect -5614 3811 -5548 3845
rect -5614 3777 -5598 3811
rect -5564 3777 -5548 3811
rect -5614 3743 -5548 3777
rect -5614 3709 -5598 3743
rect -5564 3709 -5548 3743
rect -5614 3675 -5548 3709
rect -5614 3641 -5598 3675
rect -5564 3641 -5548 3675
rect -5614 3607 -5548 3641
rect -5614 3573 -5598 3607
rect -5564 3573 -5548 3607
rect -5614 3539 -5548 3573
rect -5614 3505 -5598 3539
rect -5564 3505 -5548 3539
rect -5614 3464 -5548 3505
rect -5518 4423 -5456 4464
rect -5518 4389 -5502 4423
rect -5468 4389 -5456 4423
rect -5518 4355 -5456 4389
rect -5518 4321 -5502 4355
rect -5468 4321 -5456 4355
rect -5518 4287 -5456 4321
rect -5518 4253 -5502 4287
rect -5468 4253 -5456 4287
rect -5518 4219 -5456 4253
rect -5518 4185 -5502 4219
rect -5468 4185 -5456 4219
rect -5518 4151 -5456 4185
rect -5518 4117 -5502 4151
rect -5468 4117 -5456 4151
rect -5518 4083 -5456 4117
rect -5518 4049 -5502 4083
rect -5468 4049 -5456 4083
rect -5518 4015 -5456 4049
rect -5518 3981 -5502 4015
rect -5468 3981 -5456 4015
rect -5518 3947 -5456 3981
rect -5518 3913 -5502 3947
rect -5468 3913 -5456 3947
rect -5518 3879 -5456 3913
rect -5518 3845 -5502 3879
rect -5468 3845 -5456 3879
rect -5518 3811 -5456 3845
rect -5518 3777 -5502 3811
rect -5468 3777 -5456 3811
rect -5518 3743 -5456 3777
rect -5518 3709 -5502 3743
rect -5468 3709 -5456 3743
rect -5518 3675 -5456 3709
rect -5518 3641 -5502 3675
rect -5468 3641 -5456 3675
rect -5518 3607 -5456 3641
rect -5518 3573 -5502 3607
rect -5468 3573 -5456 3607
rect -5518 3539 -5456 3573
rect -5518 3505 -5502 3539
rect -5468 3505 -5456 3539
rect -5518 3464 -5456 3505
rect -5306 4425 -5244 4466
rect -5306 4391 -5294 4425
rect -5260 4391 -5244 4425
rect -5306 4357 -5244 4391
rect -5306 4323 -5294 4357
rect -5260 4323 -5244 4357
rect -5306 4289 -5244 4323
rect -5306 4255 -5294 4289
rect -5260 4255 -5244 4289
rect -5306 4221 -5244 4255
rect -5306 4187 -5294 4221
rect -5260 4187 -5244 4221
rect -5306 4153 -5244 4187
rect -5306 4119 -5294 4153
rect -5260 4119 -5244 4153
rect -5306 4085 -5244 4119
rect -5306 4051 -5294 4085
rect -5260 4051 -5244 4085
rect -5306 4017 -5244 4051
rect -5306 3983 -5294 4017
rect -5260 3983 -5244 4017
rect -5306 3949 -5244 3983
rect -5306 3915 -5294 3949
rect -5260 3915 -5244 3949
rect -5306 3881 -5244 3915
rect -5306 3847 -5294 3881
rect -5260 3847 -5244 3881
rect -5306 3813 -5244 3847
rect -5306 3779 -5294 3813
rect -5260 3779 -5244 3813
rect -5306 3745 -5244 3779
rect -5306 3711 -5294 3745
rect -5260 3711 -5244 3745
rect -5306 3677 -5244 3711
rect -5306 3643 -5294 3677
rect -5260 3643 -5244 3677
rect -5306 3609 -5244 3643
rect -5306 3575 -5294 3609
rect -5260 3575 -5244 3609
rect -5306 3541 -5244 3575
rect -5306 3507 -5294 3541
rect -5260 3507 -5244 3541
rect -5306 3466 -5244 3507
rect -5214 4425 -5148 4466
rect -5214 4391 -5198 4425
rect -5164 4391 -5148 4425
rect -5214 4357 -5148 4391
rect -5214 4323 -5198 4357
rect -5164 4323 -5148 4357
rect -5214 4289 -5148 4323
rect -5214 4255 -5198 4289
rect -5164 4255 -5148 4289
rect -5214 4221 -5148 4255
rect -5214 4187 -5198 4221
rect -5164 4187 -5148 4221
rect -5214 4153 -5148 4187
rect -5214 4119 -5198 4153
rect -5164 4119 -5148 4153
rect -5214 4085 -5148 4119
rect -5214 4051 -5198 4085
rect -5164 4051 -5148 4085
rect -5214 4017 -5148 4051
rect -5214 3983 -5198 4017
rect -5164 3983 -5148 4017
rect -5214 3949 -5148 3983
rect -5214 3915 -5198 3949
rect -5164 3915 -5148 3949
rect -5214 3881 -5148 3915
rect -5214 3847 -5198 3881
rect -5164 3847 -5148 3881
rect -5214 3813 -5148 3847
rect -5214 3779 -5198 3813
rect -5164 3779 -5148 3813
rect -5214 3745 -5148 3779
rect -5214 3711 -5198 3745
rect -5164 3711 -5148 3745
rect -5214 3677 -5148 3711
rect -5214 3643 -5198 3677
rect -5164 3643 -5148 3677
rect -5214 3609 -5148 3643
rect -5214 3575 -5198 3609
rect -5164 3575 -5148 3609
rect -5214 3541 -5148 3575
rect -5214 3507 -5198 3541
rect -5164 3507 -5148 3541
rect -5214 3466 -5148 3507
rect -5118 4425 -5052 4466
rect -5118 4391 -5102 4425
rect -5068 4391 -5052 4425
rect -5118 4357 -5052 4391
rect -5118 4323 -5102 4357
rect -5068 4323 -5052 4357
rect -5118 4289 -5052 4323
rect -5118 4255 -5102 4289
rect -5068 4255 -5052 4289
rect -5118 4221 -5052 4255
rect -5118 4187 -5102 4221
rect -5068 4187 -5052 4221
rect -5118 4153 -5052 4187
rect -5118 4119 -5102 4153
rect -5068 4119 -5052 4153
rect -5118 4085 -5052 4119
rect -5118 4051 -5102 4085
rect -5068 4051 -5052 4085
rect -5118 4017 -5052 4051
rect -5118 3983 -5102 4017
rect -5068 3983 -5052 4017
rect -5118 3949 -5052 3983
rect -5118 3915 -5102 3949
rect -5068 3915 -5052 3949
rect -5118 3881 -5052 3915
rect -5118 3847 -5102 3881
rect -5068 3847 -5052 3881
rect -5118 3813 -5052 3847
rect -5118 3779 -5102 3813
rect -5068 3779 -5052 3813
rect -5118 3745 -5052 3779
rect -5118 3711 -5102 3745
rect -5068 3711 -5052 3745
rect -5118 3677 -5052 3711
rect -5118 3643 -5102 3677
rect -5068 3643 -5052 3677
rect -5118 3609 -5052 3643
rect -5118 3575 -5102 3609
rect -5068 3575 -5052 3609
rect -5118 3541 -5052 3575
rect -5118 3507 -5102 3541
rect -5068 3507 -5052 3541
rect -5118 3466 -5052 3507
rect -5022 4425 -4956 4466
rect -5022 4391 -5006 4425
rect -4972 4391 -4956 4425
rect -5022 4357 -4956 4391
rect -5022 4323 -5006 4357
rect -4972 4323 -4956 4357
rect -5022 4289 -4956 4323
rect -5022 4255 -5006 4289
rect -4972 4255 -4956 4289
rect -5022 4221 -4956 4255
rect -5022 4187 -5006 4221
rect -4972 4187 -4956 4221
rect -5022 4153 -4956 4187
rect -5022 4119 -5006 4153
rect -4972 4119 -4956 4153
rect -5022 4085 -4956 4119
rect -5022 4051 -5006 4085
rect -4972 4051 -4956 4085
rect -5022 4017 -4956 4051
rect -5022 3983 -5006 4017
rect -4972 3983 -4956 4017
rect -5022 3949 -4956 3983
rect -5022 3915 -5006 3949
rect -4972 3915 -4956 3949
rect -5022 3881 -4956 3915
rect -5022 3847 -5006 3881
rect -4972 3847 -4956 3881
rect -5022 3813 -4956 3847
rect -5022 3779 -5006 3813
rect -4972 3779 -4956 3813
rect -5022 3745 -4956 3779
rect -5022 3711 -5006 3745
rect -4972 3711 -4956 3745
rect -5022 3677 -4956 3711
rect -5022 3643 -5006 3677
rect -4972 3643 -4956 3677
rect -5022 3609 -4956 3643
rect -5022 3575 -5006 3609
rect -4972 3575 -4956 3609
rect -5022 3541 -4956 3575
rect -5022 3507 -5006 3541
rect -4972 3507 -4956 3541
rect -5022 3466 -4956 3507
rect -4926 4425 -4860 4466
rect -4926 4391 -4910 4425
rect -4876 4391 -4860 4425
rect -4926 4357 -4860 4391
rect -4926 4323 -4910 4357
rect -4876 4323 -4860 4357
rect -4926 4289 -4860 4323
rect -4926 4255 -4910 4289
rect -4876 4255 -4860 4289
rect -4926 4221 -4860 4255
rect -4926 4187 -4910 4221
rect -4876 4187 -4860 4221
rect -4926 4153 -4860 4187
rect -4926 4119 -4910 4153
rect -4876 4119 -4860 4153
rect -4926 4085 -4860 4119
rect -4926 4051 -4910 4085
rect -4876 4051 -4860 4085
rect -4926 4017 -4860 4051
rect -4926 3983 -4910 4017
rect -4876 3983 -4860 4017
rect -4926 3949 -4860 3983
rect -4926 3915 -4910 3949
rect -4876 3915 -4860 3949
rect -4926 3881 -4860 3915
rect -4926 3847 -4910 3881
rect -4876 3847 -4860 3881
rect -4926 3813 -4860 3847
rect -4926 3779 -4910 3813
rect -4876 3779 -4860 3813
rect -4926 3745 -4860 3779
rect -4926 3711 -4910 3745
rect -4876 3711 -4860 3745
rect -4926 3677 -4860 3711
rect -4926 3643 -4910 3677
rect -4876 3643 -4860 3677
rect -4926 3609 -4860 3643
rect -4926 3575 -4910 3609
rect -4876 3575 -4860 3609
rect -4926 3541 -4860 3575
rect -4926 3507 -4910 3541
rect -4876 3507 -4860 3541
rect -4926 3466 -4860 3507
rect -4830 4425 -4768 4466
rect -4830 4391 -4814 4425
rect -4780 4391 -4768 4425
rect -4830 4357 -4768 4391
rect -4830 4323 -4814 4357
rect -4780 4323 -4768 4357
rect -4830 4289 -4768 4323
rect -4830 4255 -4814 4289
rect -4780 4255 -4768 4289
rect -4830 4221 -4768 4255
rect -4830 4187 -4814 4221
rect -4780 4187 -4768 4221
rect -4830 4153 -4768 4187
rect -4830 4119 -4814 4153
rect -4780 4119 -4768 4153
rect -4830 4085 -4768 4119
rect -4830 4051 -4814 4085
rect -4780 4051 -4768 4085
rect -4830 4017 -4768 4051
rect -4830 3983 -4814 4017
rect -4780 3983 -4768 4017
rect -4830 3949 -4768 3983
rect -4830 3915 -4814 3949
rect -4780 3915 -4768 3949
rect 1472 4461 1484 4495
rect 1518 4461 1534 4495
rect 1472 4427 1534 4461
rect 1472 4393 1484 4427
rect 1518 4393 1534 4427
rect 1472 4359 1534 4393
rect 1472 4325 1484 4359
rect 1518 4325 1534 4359
rect 1472 4291 1534 4325
rect 1472 4257 1484 4291
rect 1518 4257 1534 4291
rect 1472 4223 1534 4257
rect 1472 4189 1484 4223
rect 1518 4189 1534 4223
rect 1472 4155 1534 4189
rect 1472 4121 1484 4155
rect 1518 4121 1534 4155
rect 1472 4087 1534 4121
rect 1472 4053 1484 4087
rect 1518 4053 1534 4087
rect 1472 4019 1534 4053
rect 1472 3985 1484 4019
rect 1518 3985 1534 4019
rect 1472 3944 1534 3985
rect 1564 4903 1630 4944
rect 1564 4869 1580 4903
rect 1614 4869 1630 4903
rect 1564 4835 1630 4869
rect 1564 4801 1580 4835
rect 1614 4801 1630 4835
rect 1564 4767 1630 4801
rect 1564 4733 1580 4767
rect 1614 4733 1630 4767
rect 1564 4699 1630 4733
rect 1564 4665 1580 4699
rect 1614 4665 1630 4699
rect 1564 4631 1630 4665
rect 1564 4597 1580 4631
rect 1614 4597 1630 4631
rect 1564 4563 1630 4597
rect 1564 4529 1580 4563
rect 1614 4529 1630 4563
rect 1564 4495 1630 4529
rect 1564 4461 1580 4495
rect 1614 4461 1630 4495
rect 1564 4427 1630 4461
rect 1564 4393 1580 4427
rect 1614 4393 1630 4427
rect 1564 4359 1630 4393
rect 1564 4325 1580 4359
rect 1614 4325 1630 4359
rect 1564 4291 1630 4325
rect 1564 4257 1580 4291
rect 1614 4257 1630 4291
rect 1564 4223 1630 4257
rect 1564 4189 1580 4223
rect 1614 4189 1630 4223
rect 1564 4155 1630 4189
rect 1564 4121 1580 4155
rect 1614 4121 1630 4155
rect 1564 4087 1630 4121
rect 1564 4053 1580 4087
rect 1614 4053 1630 4087
rect 1564 4019 1630 4053
rect 1564 3985 1580 4019
rect 1614 3985 1630 4019
rect 1564 3944 1630 3985
rect 1660 4903 1726 4944
rect 1660 4869 1676 4903
rect 1710 4869 1726 4903
rect 1660 4835 1726 4869
rect 1660 4801 1676 4835
rect 1710 4801 1726 4835
rect 1660 4767 1726 4801
rect 1660 4733 1676 4767
rect 1710 4733 1726 4767
rect 1660 4699 1726 4733
rect 1660 4665 1676 4699
rect 1710 4665 1726 4699
rect 1660 4631 1726 4665
rect 1660 4597 1676 4631
rect 1710 4597 1726 4631
rect 1660 4563 1726 4597
rect 1660 4529 1676 4563
rect 1710 4529 1726 4563
rect 1660 4495 1726 4529
rect 1660 4461 1676 4495
rect 1710 4461 1726 4495
rect 1660 4427 1726 4461
rect 1660 4393 1676 4427
rect 1710 4393 1726 4427
rect 1660 4359 1726 4393
rect 1660 4325 1676 4359
rect 1710 4325 1726 4359
rect 1660 4291 1726 4325
rect 1660 4257 1676 4291
rect 1710 4257 1726 4291
rect 1660 4223 1726 4257
rect 1660 4189 1676 4223
rect 1710 4189 1726 4223
rect 1660 4155 1726 4189
rect 1660 4121 1676 4155
rect 1710 4121 1726 4155
rect 1660 4087 1726 4121
rect 1660 4053 1676 4087
rect 1710 4053 1726 4087
rect 1660 4019 1726 4053
rect 1660 3985 1676 4019
rect 1710 3985 1726 4019
rect 1660 3944 1726 3985
rect 1756 4903 1822 4944
rect 1756 4869 1772 4903
rect 1806 4869 1822 4903
rect 1756 4835 1822 4869
rect 1756 4801 1772 4835
rect 1806 4801 1822 4835
rect 1756 4767 1822 4801
rect 1756 4733 1772 4767
rect 1806 4733 1822 4767
rect 1756 4699 1822 4733
rect 1756 4665 1772 4699
rect 1806 4665 1822 4699
rect 1756 4631 1822 4665
rect 1756 4597 1772 4631
rect 1806 4597 1822 4631
rect 1756 4563 1822 4597
rect 1756 4529 1772 4563
rect 1806 4529 1822 4563
rect 1756 4495 1822 4529
rect 1756 4461 1772 4495
rect 1806 4461 1822 4495
rect 1756 4427 1822 4461
rect 1756 4393 1772 4427
rect 1806 4393 1822 4427
rect 1756 4359 1822 4393
rect 1756 4325 1772 4359
rect 1806 4325 1822 4359
rect 1756 4291 1822 4325
rect 1756 4257 1772 4291
rect 1806 4257 1822 4291
rect 1756 4223 1822 4257
rect 1756 4189 1772 4223
rect 1806 4189 1822 4223
rect 1756 4155 1822 4189
rect 1756 4121 1772 4155
rect 1806 4121 1822 4155
rect 1756 4087 1822 4121
rect 1756 4053 1772 4087
rect 1806 4053 1822 4087
rect 1756 4019 1822 4053
rect 1756 3985 1772 4019
rect 1806 3985 1822 4019
rect 1756 3944 1822 3985
rect 1852 4903 1914 4944
rect 15506 4977 15518 5011
rect 15552 4977 15568 5011
rect 1852 4869 1868 4903
rect 1902 4869 1914 4903
rect 1852 4835 1914 4869
rect 1852 4801 1868 4835
rect 1902 4801 1914 4835
rect 1852 4767 1914 4801
rect 1852 4733 1868 4767
rect 1902 4733 1914 4767
rect 1852 4699 1914 4733
rect 1852 4665 1868 4699
rect 1902 4665 1914 4699
rect 1852 4631 1914 4665
rect 1852 4597 1868 4631
rect 1902 4597 1914 4631
rect 1852 4563 1914 4597
rect 1852 4529 1868 4563
rect 1902 4529 1914 4563
rect 1852 4495 1914 4529
rect 1852 4461 1868 4495
rect 1902 4461 1914 4495
rect 1852 4427 1914 4461
rect 1852 4393 1868 4427
rect 1902 4393 1914 4427
rect 1852 4359 1914 4393
rect 1852 4325 1868 4359
rect 1902 4325 1914 4359
rect 1852 4291 1914 4325
rect 1852 4257 1868 4291
rect 1902 4257 1914 4291
rect 1852 4223 1914 4257
rect 1852 4189 1868 4223
rect 1902 4189 1914 4223
rect 1852 4155 1914 4189
rect 1852 4121 1868 4155
rect 1902 4121 1914 4155
rect 1852 4087 1914 4121
rect 1852 4053 1868 4087
rect 1902 4053 1914 4087
rect 1852 4019 1914 4053
rect 1852 3985 1868 4019
rect 1902 3985 1914 4019
rect 1852 3944 1914 3985
rect 4428 4887 4490 4928
rect 4428 4853 4440 4887
rect 4474 4853 4490 4887
rect 4428 4819 4490 4853
rect 4428 4785 4440 4819
rect 4474 4785 4490 4819
rect 4428 4751 4490 4785
rect 4428 4717 4440 4751
rect 4474 4717 4490 4751
rect 4428 4683 4490 4717
rect 4428 4649 4440 4683
rect 4474 4649 4490 4683
rect 4428 4615 4490 4649
rect 4428 4581 4440 4615
rect 4474 4581 4490 4615
rect 4428 4547 4490 4581
rect 4428 4513 4440 4547
rect 4474 4513 4490 4547
rect 4428 4479 4490 4513
rect 4428 4445 4440 4479
rect 4474 4445 4490 4479
rect 4428 4411 4490 4445
rect 4428 4377 4440 4411
rect 4474 4377 4490 4411
rect 4428 4343 4490 4377
rect 4428 4309 4440 4343
rect 4474 4309 4490 4343
rect 4428 4275 4490 4309
rect 4428 4241 4440 4275
rect 4474 4241 4490 4275
rect 4428 4207 4490 4241
rect 4428 4173 4440 4207
rect 4474 4173 4490 4207
rect 4428 4139 4490 4173
rect 4428 4105 4440 4139
rect 4474 4105 4490 4139
rect 4428 4071 4490 4105
rect 4428 4037 4440 4071
rect 4474 4037 4490 4071
rect 4428 4003 4490 4037
rect 4428 3969 4440 4003
rect 4474 3969 4490 4003
rect -4830 3881 -4768 3915
rect -4830 3847 -4814 3881
rect -4780 3847 -4768 3881
rect -4830 3813 -4768 3847
rect 4428 3928 4490 3969
rect 4520 4887 4586 4928
rect 4520 4853 4536 4887
rect 4570 4853 4586 4887
rect 4520 4819 4586 4853
rect 4520 4785 4536 4819
rect 4570 4785 4586 4819
rect 4520 4751 4586 4785
rect 4520 4717 4536 4751
rect 4570 4717 4586 4751
rect 4520 4683 4586 4717
rect 4520 4649 4536 4683
rect 4570 4649 4586 4683
rect 4520 4615 4586 4649
rect 4520 4581 4536 4615
rect 4570 4581 4586 4615
rect 4520 4547 4586 4581
rect 4520 4513 4536 4547
rect 4570 4513 4586 4547
rect 4520 4479 4586 4513
rect 4520 4445 4536 4479
rect 4570 4445 4586 4479
rect 4520 4411 4586 4445
rect 4520 4377 4536 4411
rect 4570 4377 4586 4411
rect 4520 4343 4586 4377
rect 4520 4309 4536 4343
rect 4570 4309 4586 4343
rect 4520 4275 4586 4309
rect 4520 4241 4536 4275
rect 4570 4241 4586 4275
rect 4520 4207 4586 4241
rect 4520 4173 4536 4207
rect 4570 4173 4586 4207
rect 4520 4139 4586 4173
rect 4520 4105 4536 4139
rect 4570 4105 4586 4139
rect 4520 4071 4586 4105
rect 4520 4037 4536 4071
rect 4570 4037 4586 4071
rect 4520 4003 4586 4037
rect 4520 3969 4536 4003
rect 4570 3969 4586 4003
rect 4520 3928 4586 3969
rect 4616 4887 4682 4928
rect 4616 4853 4632 4887
rect 4666 4853 4682 4887
rect 4616 4819 4682 4853
rect 4616 4785 4632 4819
rect 4666 4785 4682 4819
rect 4616 4751 4682 4785
rect 4616 4717 4632 4751
rect 4666 4717 4682 4751
rect 4616 4683 4682 4717
rect 4616 4649 4632 4683
rect 4666 4649 4682 4683
rect 4616 4615 4682 4649
rect 4616 4581 4632 4615
rect 4666 4581 4682 4615
rect 4616 4547 4682 4581
rect 4616 4513 4632 4547
rect 4666 4513 4682 4547
rect 4616 4479 4682 4513
rect 4616 4445 4632 4479
rect 4666 4445 4682 4479
rect 4616 4411 4682 4445
rect 4616 4377 4632 4411
rect 4666 4377 4682 4411
rect 4616 4343 4682 4377
rect 4616 4309 4632 4343
rect 4666 4309 4682 4343
rect 4616 4275 4682 4309
rect 4616 4241 4632 4275
rect 4666 4241 4682 4275
rect 4616 4207 4682 4241
rect 4616 4173 4632 4207
rect 4666 4173 4682 4207
rect 4616 4139 4682 4173
rect 4616 4105 4632 4139
rect 4666 4105 4682 4139
rect 4616 4071 4682 4105
rect 4616 4037 4632 4071
rect 4666 4037 4682 4071
rect 4616 4003 4682 4037
rect 4616 3969 4632 4003
rect 4666 3969 4682 4003
rect 4616 3928 4682 3969
rect 4712 4887 4778 4928
rect 4712 4853 4728 4887
rect 4762 4853 4778 4887
rect 4712 4819 4778 4853
rect 4712 4785 4728 4819
rect 4762 4785 4778 4819
rect 4712 4751 4778 4785
rect 4712 4717 4728 4751
rect 4762 4717 4778 4751
rect 4712 4683 4778 4717
rect 4712 4649 4728 4683
rect 4762 4649 4778 4683
rect 4712 4615 4778 4649
rect 4712 4581 4728 4615
rect 4762 4581 4778 4615
rect 4712 4547 4778 4581
rect 4712 4513 4728 4547
rect 4762 4513 4778 4547
rect 4712 4479 4778 4513
rect 4712 4445 4728 4479
rect 4762 4445 4778 4479
rect 4712 4411 4778 4445
rect 4712 4377 4728 4411
rect 4762 4377 4778 4411
rect 4712 4343 4778 4377
rect 4712 4309 4728 4343
rect 4762 4309 4778 4343
rect 4712 4275 4778 4309
rect 4712 4241 4728 4275
rect 4762 4241 4778 4275
rect 4712 4207 4778 4241
rect 4712 4173 4728 4207
rect 4762 4173 4778 4207
rect 4712 4139 4778 4173
rect 4712 4105 4728 4139
rect 4762 4105 4778 4139
rect 4712 4071 4778 4105
rect 4712 4037 4728 4071
rect 4762 4037 4778 4071
rect 4712 4003 4778 4037
rect 4712 3969 4728 4003
rect 4762 3969 4778 4003
rect 4712 3928 4778 3969
rect 4808 4887 4870 4928
rect 4808 4853 4824 4887
rect 4858 4853 4870 4887
rect 4808 4819 4870 4853
rect 4808 4785 4824 4819
rect 4858 4785 4870 4819
rect 4808 4751 4870 4785
rect 4808 4717 4824 4751
rect 4858 4717 4870 4751
rect 4808 4683 4870 4717
rect 4808 4649 4824 4683
rect 4858 4649 4870 4683
rect 4808 4615 4870 4649
rect 4808 4581 4824 4615
rect 4858 4581 4870 4615
rect 4808 4547 4870 4581
rect 4808 4513 4824 4547
rect 4858 4513 4870 4547
rect 4808 4479 4870 4513
rect 4808 4445 4824 4479
rect 4858 4445 4870 4479
rect 4808 4411 4870 4445
rect 4808 4377 4824 4411
rect 4858 4377 4870 4411
rect 4808 4343 4870 4377
rect 4808 4309 4824 4343
rect 4858 4309 4870 4343
rect 4808 4275 4870 4309
rect 4808 4241 4824 4275
rect 4858 4241 4870 4275
rect 4808 4207 4870 4241
rect 4808 4173 4824 4207
rect 4858 4173 4870 4207
rect 4808 4139 4870 4173
rect 4808 4105 4824 4139
rect 4858 4105 4870 4139
rect 4808 4071 4870 4105
rect 4808 4037 4824 4071
rect 4858 4037 4870 4071
rect 4808 4003 4870 4037
rect 4808 3969 4824 4003
rect 4858 3969 4870 4003
rect 4808 3928 4870 3969
rect 7458 4887 7520 4928
rect 7458 4853 7470 4887
rect 7504 4853 7520 4887
rect 7458 4819 7520 4853
rect 7458 4785 7470 4819
rect 7504 4785 7520 4819
rect 7458 4751 7520 4785
rect 7458 4717 7470 4751
rect 7504 4717 7520 4751
rect 7458 4683 7520 4717
rect 7458 4649 7470 4683
rect 7504 4649 7520 4683
rect 7458 4615 7520 4649
rect 7458 4581 7470 4615
rect 7504 4581 7520 4615
rect 7458 4547 7520 4581
rect 7458 4513 7470 4547
rect 7504 4513 7520 4547
rect 7458 4479 7520 4513
rect 7458 4445 7470 4479
rect 7504 4445 7520 4479
rect 7458 4411 7520 4445
rect 7458 4377 7470 4411
rect 7504 4377 7520 4411
rect 7458 4343 7520 4377
rect 7458 4309 7470 4343
rect 7504 4309 7520 4343
rect 7458 4275 7520 4309
rect 7458 4241 7470 4275
rect 7504 4241 7520 4275
rect 7458 4207 7520 4241
rect 7458 4173 7470 4207
rect 7504 4173 7520 4207
rect 7458 4139 7520 4173
rect 7458 4105 7470 4139
rect 7504 4105 7520 4139
rect 7458 4071 7520 4105
rect 7458 4037 7470 4071
rect 7504 4037 7520 4071
rect 7458 4003 7520 4037
rect 7458 3969 7470 4003
rect 7504 3969 7520 4003
rect 7458 3928 7520 3969
rect 7550 4887 7616 4928
rect 7550 4853 7566 4887
rect 7600 4853 7616 4887
rect 7550 4819 7616 4853
rect 7550 4785 7566 4819
rect 7600 4785 7616 4819
rect 7550 4751 7616 4785
rect 7550 4717 7566 4751
rect 7600 4717 7616 4751
rect 7550 4683 7616 4717
rect 7550 4649 7566 4683
rect 7600 4649 7616 4683
rect 7550 4615 7616 4649
rect 7550 4581 7566 4615
rect 7600 4581 7616 4615
rect 7550 4547 7616 4581
rect 7550 4513 7566 4547
rect 7600 4513 7616 4547
rect 7550 4479 7616 4513
rect 7550 4445 7566 4479
rect 7600 4445 7616 4479
rect 7550 4411 7616 4445
rect 7550 4377 7566 4411
rect 7600 4377 7616 4411
rect 7550 4343 7616 4377
rect 7550 4309 7566 4343
rect 7600 4309 7616 4343
rect 7550 4275 7616 4309
rect 7550 4241 7566 4275
rect 7600 4241 7616 4275
rect 7550 4207 7616 4241
rect 7550 4173 7566 4207
rect 7600 4173 7616 4207
rect 7550 4139 7616 4173
rect 7550 4105 7566 4139
rect 7600 4105 7616 4139
rect 7550 4071 7616 4105
rect 7550 4037 7566 4071
rect 7600 4037 7616 4071
rect 7550 4003 7616 4037
rect 7550 3969 7566 4003
rect 7600 3969 7616 4003
rect 7550 3928 7616 3969
rect 7646 4887 7712 4928
rect 7646 4853 7662 4887
rect 7696 4853 7712 4887
rect 7646 4819 7712 4853
rect 7646 4785 7662 4819
rect 7696 4785 7712 4819
rect 7646 4751 7712 4785
rect 7646 4717 7662 4751
rect 7696 4717 7712 4751
rect 7646 4683 7712 4717
rect 7646 4649 7662 4683
rect 7696 4649 7712 4683
rect 7646 4615 7712 4649
rect 7646 4581 7662 4615
rect 7696 4581 7712 4615
rect 7646 4547 7712 4581
rect 7646 4513 7662 4547
rect 7696 4513 7712 4547
rect 7646 4479 7712 4513
rect 7646 4445 7662 4479
rect 7696 4445 7712 4479
rect 7646 4411 7712 4445
rect 7646 4377 7662 4411
rect 7696 4377 7712 4411
rect 7646 4343 7712 4377
rect 7646 4309 7662 4343
rect 7696 4309 7712 4343
rect 7646 4275 7712 4309
rect 7646 4241 7662 4275
rect 7696 4241 7712 4275
rect 7646 4207 7712 4241
rect 7646 4173 7662 4207
rect 7696 4173 7712 4207
rect 7646 4139 7712 4173
rect 7646 4105 7662 4139
rect 7696 4105 7712 4139
rect 7646 4071 7712 4105
rect 7646 4037 7662 4071
rect 7696 4037 7712 4071
rect 7646 4003 7712 4037
rect 7646 3969 7662 4003
rect 7696 3969 7712 4003
rect 7646 3928 7712 3969
rect 7742 4887 7808 4928
rect 7742 4853 7758 4887
rect 7792 4853 7808 4887
rect 7742 4819 7808 4853
rect 7742 4785 7758 4819
rect 7792 4785 7808 4819
rect 7742 4751 7808 4785
rect 7742 4717 7758 4751
rect 7792 4717 7808 4751
rect 7742 4683 7808 4717
rect 7742 4649 7758 4683
rect 7792 4649 7808 4683
rect 7742 4615 7808 4649
rect 7742 4581 7758 4615
rect 7792 4581 7808 4615
rect 7742 4547 7808 4581
rect 7742 4513 7758 4547
rect 7792 4513 7808 4547
rect 7742 4479 7808 4513
rect 7742 4445 7758 4479
rect 7792 4445 7808 4479
rect 7742 4411 7808 4445
rect 7742 4377 7758 4411
rect 7792 4377 7808 4411
rect 7742 4343 7808 4377
rect 7742 4309 7758 4343
rect 7792 4309 7808 4343
rect 7742 4275 7808 4309
rect 7742 4241 7758 4275
rect 7792 4241 7808 4275
rect 7742 4207 7808 4241
rect 7742 4173 7758 4207
rect 7792 4173 7808 4207
rect 7742 4139 7808 4173
rect 7742 4105 7758 4139
rect 7792 4105 7808 4139
rect 7742 4071 7808 4105
rect 7742 4037 7758 4071
rect 7792 4037 7808 4071
rect 7742 4003 7808 4037
rect 7742 3969 7758 4003
rect 7792 3969 7808 4003
rect 7742 3928 7808 3969
rect 7838 4887 7900 4928
rect 7838 4853 7854 4887
rect 7888 4853 7900 4887
rect 7838 4819 7900 4853
rect 7838 4785 7854 4819
rect 7888 4785 7900 4819
rect 7838 4751 7900 4785
rect 7838 4717 7854 4751
rect 7888 4717 7900 4751
rect 7838 4683 7900 4717
rect 7838 4649 7854 4683
rect 7888 4649 7900 4683
rect 7838 4615 7900 4649
rect 7838 4581 7854 4615
rect 7888 4581 7900 4615
rect 7838 4547 7900 4581
rect 7838 4513 7854 4547
rect 7888 4513 7900 4547
rect 7838 4479 7900 4513
rect 7838 4445 7854 4479
rect 7888 4445 7900 4479
rect 7838 4411 7900 4445
rect 7838 4377 7854 4411
rect 7888 4377 7900 4411
rect 7838 4343 7900 4377
rect 7838 4309 7854 4343
rect 7888 4309 7900 4343
rect 7838 4275 7900 4309
rect 7838 4241 7854 4275
rect 7888 4241 7900 4275
rect 7838 4207 7900 4241
rect 7838 4173 7854 4207
rect 7888 4173 7900 4207
rect 7838 4139 7900 4173
rect 7838 4105 7854 4139
rect 7888 4105 7900 4139
rect 7838 4071 7900 4105
rect 7838 4037 7854 4071
rect 7888 4037 7900 4071
rect 7838 4003 7900 4037
rect 7838 3969 7854 4003
rect 7888 3969 7900 4003
rect 7838 3928 7900 3969
rect 10546 4885 10608 4926
rect 10546 4851 10558 4885
rect 10592 4851 10608 4885
rect 10546 4817 10608 4851
rect 10546 4783 10558 4817
rect 10592 4783 10608 4817
rect 10546 4749 10608 4783
rect 10546 4715 10558 4749
rect 10592 4715 10608 4749
rect 10546 4681 10608 4715
rect 10546 4647 10558 4681
rect 10592 4647 10608 4681
rect 10546 4613 10608 4647
rect 10546 4579 10558 4613
rect 10592 4579 10608 4613
rect 10546 4545 10608 4579
rect 10546 4511 10558 4545
rect 10592 4511 10608 4545
rect 10546 4477 10608 4511
rect 10546 4443 10558 4477
rect 10592 4443 10608 4477
rect 10546 4409 10608 4443
rect 10546 4375 10558 4409
rect 10592 4375 10608 4409
rect 10546 4341 10608 4375
rect 10546 4307 10558 4341
rect 10592 4307 10608 4341
rect 10546 4273 10608 4307
rect 10546 4239 10558 4273
rect 10592 4239 10608 4273
rect 10546 4205 10608 4239
rect 10546 4171 10558 4205
rect 10592 4171 10608 4205
rect 10546 4137 10608 4171
rect 10546 4103 10558 4137
rect 10592 4103 10608 4137
rect 10546 4069 10608 4103
rect 10546 4035 10558 4069
rect 10592 4035 10608 4069
rect 10546 4001 10608 4035
rect 10546 3967 10558 4001
rect 10592 3967 10608 4001
rect -4830 3779 -4814 3813
rect -4780 3779 -4768 3813
rect 10546 3926 10608 3967
rect 10638 4885 10704 4926
rect 10638 4851 10654 4885
rect 10688 4851 10704 4885
rect 10638 4817 10704 4851
rect 10638 4783 10654 4817
rect 10688 4783 10704 4817
rect 10638 4749 10704 4783
rect 10638 4715 10654 4749
rect 10688 4715 10704 4749
rect 10638 4681 10704 4715
rect 10638 4647 10654 4681
rect 10688 4647 10704 4681
rect 10638 4613 10704 4647
rect 10638 4579 10654 4613
rect 10688 4579 10704 4613
rect 10638 4545 10704 4579
rect 10638 4511 10654 4545
rect 10688 4511 10704 4545
rect 10638 4477 10704 4511
rect 10638 4443 10654 4477
rect 10688 4443 10704 4477
rect 10638 4409 10704 4443
rect 10638 4375 10654 4409
rect 10688 4375 10704 4409
rect 10638 4341 10704 4375
rect 10638 4307 10654 4341
rect 10688 4307 10704 4341
rect 10638 4273 10704 4307
rect 10638 4239 10654 4273
rect 10688 4239 10704 4273
rect 10638 4205 10704 4239
rect 10638 4171 10654 4205
rect 10688 4171 10704 4205
rect 10638 4137 10704 4171
rect 10638 4103 10654 4137
rect 10688 4103 10704 4137
rect 10638 4069 10704 4103
rect 10638 4035 10654 4069
rect 10688 4035 10704 4069
rect 10638 4001 10704 4035
rect 10638 3967 10654 4001
rect 10688 3967 10704 4001
rect 10638 3926 10704 3967
rect 10734 4885 10800 4926
rect 10734 4851 10750 4885
rect 10784 4851 10800 4885
rect 10734 4817 10800 4851
rect 10734 4783 10750 4817
rect 10784 4783 10800 4817
rect 10734 4749 10800 4783
rect 10734 4715 10750 4749
rect 10784 4715 10800 4749
rect 10734 4681 10800 4715
rect 10734 4647 10750 4681
rect 10784 4647 10800 4681
rect 10734 4613 10800 4647
rect 10734 4579 10750 4613
rect 10784 4579 10800 4613
rect 10734 4545 10800 4579
rect 10734 4511 10750 4545
rect 10784 4511 10800 4545
rect 10734 4477 10800 4511
rect 10734 4443 10750 4477
rect 10784 4443 10800 4477
rect 10734 4409 10800 4443
rect 10734 4375 10750 4409
rect 10784 4375 10800 4409
rect 10734 4341 10800 4375
rect 10734 4307 10750 4341
rect 10784 4307 10800 4341
rect 10734 4273 10800 4307
rect 10734 4239 10750 4273
rect 10784 4239 10800 4273
rect 10734 4205 10800 4239
rect 10734 4171 10750 4205
rect 10784 4171 10800 4205
rect 10734 4137 10800 4171
rect 10734 4103 10750 4137
rect 10784 4103 10800 4137
rect 10734 4069 10800 4103
rect 10734 4035 10750 4069
rect 10784 4035 10800 4069
rect 10734 4001 10800 4035
rect 10734 3967 10750 4001
rect 10784 3967 10800 4001
rect 10734 3926 10800 3967
rect 10830 4885 10896 4926
rect 10830 4851 10846 4885
rect 10880 4851 10896 4885
rect 10830 4817 10896 4851
rect 10830 4783 10846 4817
rect 10880 4783 10896 4817
rect 10830 4749 10896 4783
rect 10830 4715 10846 4749
rect 10880 4715 10896 4749
rect 10830 4681 10896 4715
rect 10830 4647 10846 4681
rect 10880 4647 10896 4681
rect 10830 4613 10896 4647
rect 10830 4579 10846 4613
rect 10880 4579 10896 4613
rect 10830 4545 10896 4579
rect 10830 4511 10846 4545
rect 10880 4511 10896 4545
rect 10830 4477 10896 4511
rect 10830 4443 10846 4477
rect 10880 4443 10896 4477
rect 10830 4409 10896 4443
rect 10830 4375 10846 4409
rect 10880 4375 10896 4409
rect 10830 4341 10896 4375
rect 10830 4307 10846 4341
rect 10880 4307 10896 4341
rect 10830 4273 10896 4307
rect 10830 4239 10846 4273
rect 10880 4239 10896 4273
rect 10830 4205 10896 4239
rect 10830 4171 10846 4205
rect 10880 4171 10896 4205
rect 10830 4137 10896 4171
rect 10830 4103 10846 4137
rect 10880 4103 10896 4137
rect 10830 4069 10896 4103
rect 10830 4035 10846 4069
rect 10880 4035 10896 4069
rect 10830 4001 10896 4035
rect 10830 3967 10846 4001
rect 10880 3967 10896 4001
rect 10830 3926 10896 3967
rect 10926 4885 10988 4926
rect 15506 4943 15568 4977
rect 15506 4909 15518 4943
rect 15552 4909 15568 4943
rect 10926 4851 10942 4885
rect 10976 4851 10988 4885
rect 10926 4817 10988 4851
rect 10926 4783 10942 4817
rect 10976 4783 10988 4817
rect 10926 4749 10988 4783
rect 10926 4715 10942 4749
rect 10976 4715 10988 4749
rect 10926 4681 10988 4715
rect 10926 4647 10942 4681
rect 10976 4647 10988 4681
rect 10926 4613 10988 4647
rect 10926 4579 10942 4613
rect 10976 4579 10988 4613
rect 10926 4545 10988 4579
rect 10926 4511 10942 4545
rect 10976 4511 10988 4545
rect 10926 4477 10988 4511
rect 10926 4443 10942 4477
rect 10976 4443 10988 4477
rect 10926 4409 10988 4443
rect 10926 4375 10942 4409
rect 10976 4375 10988 4409
rect 10926 4341 10988 4375
rect 10926 4307 10942 4341
rect 10976 4307 10988 4341
rect 10926 4273 10988 4307
rect 10926 4239 10942 4273
rect 10976 4239 10988 4273
rect 10926 4205 10988 4239
rect 10926 4171 10942 4205
rect 10976 4171 10988 4205
rect 10926 4137 10988 4171
rect 10926 4103 10942 4137
rect 10976 4103 10988 4137
rect 10926 4069 10988 4103
rect 10926 4035 10942 4069
rect 10976 4035 10988 4069
rect 10926 4001 10988 4035
rect 10926 3967 10942 4001
rect 10976 3967 10988 4001
rect 10926 3926 10988 3967
rect 13702 4859 13764 4900
rect 13702 4825 13714 4859
rect 13748 4825 13764 4859
rect 13702 4791 13764 4825
rect 13702 4757 13714 4791
rect 13748 4757 13764 4791
rect 13702 4723 13764 4757
rect 13702 4689 13714 4723
rect 13748 4689 13764 4723
rect 13702 4655 13764 4689
rect 13702 4621 13714 4655
rect 13748 4621 13764 4655
rect 13702 4587 13764 4621
rect 13702 4553 13714 4587
rect 13748 4553 13764 4587
rect 13702 4519 13764 4553
rect 13702 4485 13714 4519
rect 13748 4485 13764 4519
rect 13702 4451 13764 4485
rect 13702 4417 13714 4451
rect 13748 4417 13764 4451
rect 13702 4383 13764 4417
rect 13702 4349 13714 4383
rect 13748 4349 13764 4383
rect 13702 4315 13764 4349
rect 13702 4281 13714 4315
rect 13748 4281 13764 4315
rect 13702 4247 13764 4281
rect 13702 4213 13714 4247
rect 13748 4213 13764 4247
rect 13702 4179 13764 4213
rect 13702 4145 13714 4179
rect 13748 4145 13764 4179
rect 13702 4111 13764 4145
rect 13702 4077 13714 4111
rect 13748 4077 13764 4111
rect 13702 4043 13764 4077
rect 13702 4009 13714 4043
rect 13748 4009 13764 4043
rect 13702 3975 13764 4009
rect 13702 3941 13714 3975
rect 13748 3941 13764 3975
rect -4830 3745 -4768 3779
rect -4830 3711 -4814 3745
rect -4780 3711 -4768 3745
rect 13702 3900 13764 3941
rect 13794 4859 13860 4900
rect 13794 4825 13810 4859
rect 13844 4825 13860 4859
rect 13794 4791 13860 4825
rect 13794 4757 13810 4791
rect 13844 4757 13860 4791
rect 13794 4723 13860 4757
rect 13794 4689 13810 4723
rect 13844 4689 13860 4723
rect 13794 4655 13860 4689
rect 13794 4621 13810 4655
rect 13844 4621 13860 4655
rect 13794 4587 13860 4621
rect 13794 4553 13810 4587
rect 13844 4553 13860 4587
rect 13794 4519 13860 4553
rect 13794 4485 13810 4519
rect 13844 4485 13860 4519
rect 13794 4451 13860 4485
rect 13794 4417 13810 4451
rect 13844 4417 13860 4451
rect 13794 4383 13860 4417
rect 13794 4349 13810 4383
rect 13844 4349 13860 4383
rect 13794 4315 13860 4349
rect 13794 4281 13810 4315
rect 13844 4281 13860 4315
rect 13794 4247 13860 4281
rect 13794 4213 13810 4247
rect 13844 4213 13860 4247
rect 13794 4179 13860 4213
rect 13794 4145 13810 4179
rect 13844 4145 13860 4179
rect 13794 4111 13860 4145
rect 13794 4077 13810 4111
rect 13844 4077 13860 4111
rect 13794 4043 13860 4077
rect 13794 4009 13810 4043
rect 13844 4009 13860 4043
rect 13794 3975 13860 4009
rect 13794 3941 13810 3975
rect 13844 3941 13860 3975
rect 13794 3900 13860 3941
rect 13890 4859 13956 4900
rect 13890 4825 13906 4859
rect 13940 4825 13956 4859
rect 13890 4791 13956 4825
rect 13890 4757 13906 4791
rect 13940 4757 13956 4791
rect 13890 4723 13956 4757
rect 13890 4689 13906 4723
rect 13940 4689 13956 4723
rect 13890 4655 13956 4689
rect 13890 4621 13906 4655
rect 13940 4621 13956 4655
rect 13890 4587 13956 4621
rect 13890 4553 13906 4587
rect 13940 4553 13956 4587
rect 13890 4519 13956 4553
rect 13890 4485 13906 4519
rect 13940 4485 13956 4519
rect 13890 4451 13956 4485
rect 13890 4417 13906 4451
rect 13940 4417 13956 4451
rect 13890 4383 13956 4417
rect 13890 4349 13906 4383
rect 13940 4349 13956 4383
rect 13890 4315 13956 4349
rect 13890 4281 13906 4315
rect 13940 4281 13956 4315
rect 13890 4247 13956 4281
rect 13890 4213 13906 4247
rect 13940 4213 13956 4247
rect 13890 4179 13956 4213
rect 13890 4145 13906 4179
rect 13940 4145 13956 4179
rect 13890 4111 13956 4145
rect 13890 4077 13906 4111
rect 13940 4077 13956 4111
rect 13890 4043 13956 4077
rect 13890 4009 13906 4043
rect 13940 4009 13956 4043
rect 13890 3975 13956 4009
rect 13890 3941 13906 3975
rect 13940 3941 13956 3975
rect 13890 3900 13956 3941
rect 13986 4859 14052 4900
rect 13986 4825 14002 4859
rect 14036 4825 14052 4859
rect 13986 4791 14052 4825
rect 13986 4757 14002 4791
rect 14036 4757 14052 4791
rect 13986 4723 14052 4757
rect 13986 4689 14002 4723
rect 14036 4689 14052 4723
rect 13986 4655 14052 4689
rect 13986 4621 14002 4655
rect 14036 4621 14052 4655
rect 13986 4587 14052 4621
rect 13986 4553 14002 4587
rect 14036 4553 14052 4587
rect 13986 4519 14052 4553
rect 13986 4485 14002 4519
rect 14036 4485 14052 4519
rect 13986 4451 14052 4485
rect 13986 4417 14002 4451
rect 14036 4417 14052 4451
rect 13986 4383 14052 4417
rect 13986 4349 14002 4383
rect 14036 4349 14052 4383
rect 13986 4315 14052 4349
rect 13986 4281 14002 4315
rect 14036 4281 14052 4315
rect 13986 4247 14052 4281
rect 13986 4213 14002 4247
rect 14036 4213 14052 4247
rect 13986 4179 14052 4213
rect 13986 4145 14002 4179
rect 14036 4145 14052 4179
rect 13986 4111 14052 4145
rect 13986 4077 14002 4111
rect 14036 4077 14052 4111
rect 13986 4043 14052 4077
rect 13986 4009 14002 4043
rect 14036 4009 14052 4043
rect 13986 3975 14052 4009
rect 13986 3941 14002 3975
rect 14036 3941 14052 3975
rect 13986 3900 14052 3941
rect 14082 4859 14144 4900
rect 14082 4825 14098 4859
rect 14132 4825 14144 4859
rect 14082 4791 14144 4825
rect 14082 4757 14098 4791
rect 14132 4757 14144 4791
rect 14082 4723 14144 4757
rect 14082 4689 14098 4723
rect 14132 4689 14144 4723
rect 14082 4655 14144 4689
rect 14082 4621 14098 4655
rect 14132 4621 14144 4655
rect 14082 4587 14144 4621
rect 14082 4553 14098 4587
rect 14132 4553 14144 4587
rect 14082 4519 14144 4553
rect 14082 4485 14098 4519
rect 14132 4485 14144 4519
rect 14082 4451 14144 4485
rect 14082 4417 14098 4451
rect 14132 4417 14144 4451
rect 14082 4383 14144 4417
rect 14082 4349 14098 4383
rect 14132 4349 14144 4383
rect 14082 4315 14144 4349
rect 14082 4281 14098 4315
rect 14132 4281 14144 4315
rect 14082 4247 14144 4281
rect 14082 4213 14098 4247
rect 14132 4213 14144 4247
rect 14082 4179 14144 4213
rect 14082 4145 14098 4179
rect 14132 4145 14144 4179
rect 14082 4111 14144 4145
rect 14082 4077 14098 4111
rect 14132 4077 14144 4111
rect 14082 4043 14144 4077
rect 14082 4009 14098 4043
rect 14132 4009 14144 4043
rect 14082 3975 14144 4009
rect 14082 3941 14098 3975
rect 14132 3941 14144 3975
rect 14082 3900 14144 3941
rect 15506 4875 15568 4909
rect 15506 4841 15518 4875
rect 15552 4841 15568 4875
rect 15506 4807 15568 4841
rect 15506 4773 15518 4807
rect 15552 4773 15568 4807
rect 15506 4739 15568 4773
rect 15506 4705 15518 4739
rect 15552 4705 15568 4739
rect 15506 4671 15568 4705
rect 15506 4637 15518 4671
rect 15552 4637 15568 4671
rect 15506 4603 15568 4637
rect 15506 4569 15518 4603
rect 15552 4569 15568 4603
rect 15506 4535 15568 4569
rect 15506 4501 15518 4535
rect 15552 4501 15568 4535
rect 15506 4467 15568 4501
rect 15506 4433 15518 4467
rect 15552 4433 15568 4467
rect 15506 4399 15568 4433
rect 15506 4365 15518 4399
rect 15552 4365 15568 4399
rect 15506 4331 15568 4365
rect 15506 4297 15518 4331
rect 15552 4297 15568 4331
rect 15506 4263 15568 4297
rect 15506 4229 15518 4263
rect 15552 4229 15568 4263
rect 15506 4195 15568 4229
rect 15506 4161 15518 4195
rect 15552 4161 15568 4195
rect 15506 4127 15568 4161
rect 15506 4093 15518 4127
rect 15552 4093 15568 4127
rect 15506 4059 15568 4093
rect 15506 4025 15518 4059
rect 15552 4025 15568 4059
rect 15506 3991 15568 4025
rect 15506 3957 15518 3991
rect 15552 3957 15568 3991
rect 15506 3926 15568 3957
rect 15598 5895 15664 5926
rect 15598 5861 15614 5895
rect 15648 5861 15664 5895
rect 15598 5827 15664 5861
rect 15598 5793 15614 5827
rect 15648 5793 15664 5827
rect 15598 5759 15664 5793
rect 15598 5725 15614 5759
rect 15648 5725 15664 5759
rect 15598 5691 15664 5725
rect 15598 5657 15614 5691
rect 15648 5657 15664 5691
rect 15598 5623 15664 5657
rect 15598 5589 15614 5623
rect 15648 5589 15664 5623
rect 15598 5555 15664 5589
rect 15598 5521 15614 5555
rect 15648 5521 15664 5555
rect 15598 5487 15664 5521
rect 15598 5453 15614 5487
rect 15648 5453 15664 5487
rect 15598 5419 15664 5453
rect 15598 5385 15614 5419
rect 15648 5385 15664 5419
rect 15598 5351 15664 5385
rect 15598 5317 15614 5351
rect 15648 5317 15664 5351
rect 15598 5283 15664 5317
rect 15598 5249 15614 5283
rect 15648 5249 15664 5283
rect 15598 5215 15664 5249
rect 15598 5181 15614 5215
rect 15648 5181 15664 5215
rect 15598 5147 15664 5181
rect 15598 5113 15614 5147
rect 15648 5113 15664 5147
rect 15598 5079 15664 5113
rect 15598 5045 15614 5079
rect 15648 5045 15664 5079
rect 15598 5011 15664 5045
rect 15598 4977 15614 5011
rect 15648 4977 15664 5011
rect 15598 4943 15664 4977
rect 15598 4909 15614 4943
rect 15648 4909 15664 4943
rect 15598 4875 15664 4909
rect 15598 4841 15614 4875
rect 15648 4841 15664 4875
rect 15598 4807 15664 4841
rect 15598 4773 15614 4807
rect 15648 4773 15664 4807
rect 15598 4739 15664 4773
rect 15598 4705 15614 4739
rect 15648 4705 15664 4739
rect 15598 4671 15664 4705
rect 15598 4637 15614 4671
rect 15648 4637 15664 4671
rect 15598 4603 15664 4637
rect 15598 4569 15614 4603
rect 15648 4569 15664 4603
rect 15598 4535 15664 4569
rect 15598 4501 15614 4535
rect 15648 4501 15664 4535
rect 15598 4467 15664 4501
rect 15598 4433 15614 4467
rect 15648 4433 15664 4467
rect 15598 4399 15664 4433
rect 15598 4365 15614 4399
rect 15648 4365 15664 4399
rect 15598 4331 15664 4365
rect 15598 4297 15614 4331
rect 15648 4297 15664 4331
rect 15598 4263 15664 4297
rect 15598 4229 15614 4263
rect 15648 4229 15664 4263
rect 15598 4195 15664 4229
rect 15598 4161 15614 4195
rect 15648 4161 15664 4195
rect 15598 4127 15664 4161
rect 15598 4093 15614 4127
rect 15648 4093 15664 4127
rect 15598 4059 15664 4093
rect 15598 4025 15614 4059
rect 15648 4025 15664 4059
rect 15598 3991 15664 4025
rect 15598 3957 15614 3991
rect 15648 3957 15664 3991
rect 15598 3926 15664 3957
rect 15694 5895 15756 5926
rect 15694 5861 15710 5895
rect 15744 5861 15756 5895
rect 15694 5827 15756 5861
rect 15694 5793 15710 5827
rect 15744 5793 15756 5827
rect 15694 5759 15756 5793
rect 15694 5725 15710 5759
rect 15744 5725 15756 5759
rect 15694 5691 15756 5725
rect 15694 5657 15710 5691
rect 15744 5657 15756 5691
rect 15694 5623 15756 5657
rect 15694 5589 15710 5623
rect 15744 5589 15756 5623
rect 15694 5555 15756 5589
rect 15694 5521 15710 5555
rect 15744 5521 15756 5555
rect 15694 5487 15756 5521
rect 15694 5453 15710 5487
rect 15744 5453 15756 5487
rect 15694 5419 15756 5453
rect 15694 5385 15710 5419
rect 15744 5385 15756 5419
rect 15694 5351 15756 5385
rect 15694 5317 15710 5351
rect 15744 5317 15756 5351
rect 15694 5283 15756 5317
rect 15694 5249 15710 5283
rect 15744 5249 15756 5283
rect 15694 5215 15756 5249
rect 15694 5181 15710 5215
rect 15744 5181 15756 5215
rect 15694 5147 15756 5181
rect 15694 5113 15710 5147
rect 15744 5113 15756 5147
rect 15694 5079 15756 5113
rect 15694 5045 15710 5079
rect 15744 5045 15756 5079
rect 15694 5011 15756 5045
rect 15694 4977 15710 5011
rect 15744 4977 15756 5011
rect 15694 4943 15756 4977
rect 15694 4909 15710 4943
rect 15744 4909 15756 4943
rect 15694 4875 15756 4909
rect 15694 4841 15710 4875
rect 15744 4841 15756 4875
rect 15694 4807 15756 4841
rect 15694 4773 15710 4807
rect 15744 4773 15756 4807
rect 15694 4739 15756 4773
rect 15694 4705 15710 4739
rect 15744 4705 15756 4739
rect 15694 4671 15756 4705
rect 15694 4637 15710 4671
rect 15744 4637 15756 4671
rect 15694 4603 15756 4637
rect 15694 4569 15710 4603
rect 15744 4569 15756 4603
rect 15694 4535 15756 4569
rect 15694 4501 15710 4535
rect 15744 4501 15756 4535
rect 15694 4467 15756 4501
rect 15694 4433 15710 4467
rect 15744 4433 15756 4467
rect 15694 4399 15756 4433
rect 15694 4365 15710 4399
rect 15744 4365 15756 4399
rect 15694 4331 15756 4365
rect 15694 4297 15710 4331
rect 15744 4297 15756 4331
rect 15694 4263 15756 4297
rect 15694 4229 15710 4263
rect 15744 4229 15756 4263
rect 15694 4195 15756 4229
rect 15694 4161 15710 4195
rect 15744 4161 15756 4195
rect 15694 4127 15756 4161
rect 16770 5089 16832 5130
rect 16770 5055 16782 5089
rect 16816 5055 16832 5089
rect 16770 5021 16832 5055
rect 16770 4987 16782 5021
rect 16816 4987 16832 5021
rect 16770 4953 16832 4987
rect 16770 4919 16782 4953
rect 16816 4919 16832 4953
rect 16770 4885 16832 4919
rect 16770 4851 16782 4885
rect 16816 4851 16832 4885
rect 16770 4817 16832 4851
rect 16770 4783 16782 4817
rect 16816 4783 16832 4817
rect 16770 4749 16832 4783
rect 16770 4715 16782 4749
rect 16816 4715 16832 4749
rect 16770 4681 16832 4715
rect 16770 4647 16782 4681
rect 16816 4647 16832 4681
rect 16770 4613 16832 4647
rect 16770 4579 16782 4613
rect 16816 4579 16832 4613
rect 16770 4545 16832 4579
rect 16770 4511 16782 4545
rect 16816 4511 16832 4545
rect 16770 4477 16832 4511
rect 16770 4443 16782 4477
rect 16816 4443 16832 4477
rect 16770 4409 16832 4443
rect 16770 4375 16782 4409
rect 16816 4375 16832 4409
rect 16770 4341 16832 4375
rect 16770 4307 16782 4341
rect 16816 4307 16832 4341
rect 16770 4273 16832 4307
rect 16770 4239 16782 4273
rect 16816 4239 16832 4273
rect 16770 4205 16832 4239
rect 16770 4171 16782 4205
rect 16816 4171 16832 4205
rect 16770 4130 16832 4171
rect 16862 5089 16928 5130
rect 16862 5055 16878 5089
rect 16912 5055 16928 5089
rect 16862 5021 16928 5055
rect 16862 4987 16878 5021
rect 16912 4987 16928 5021
rect 16862 4953 16928 4987
rect 16862 4919 16878 4953
rect 16912 4919 16928 4953
rect 16862 4885 16928 4919
rect 16862 4851 16878 4885
rect 16912 4851 16928 4885
rect 16862 4817 16928 4851
rect 16862 4783 16878 4817
rect 16912 4783 16928 4817
rect 16862 4749 16928 4783
rect 16862 4715 16878 4749
rect 16912 4715 16928 4749
rect 16862 4681 16928 4715
rect 16862 4647 16878 4681
rect 16912 4647 16928 4681
rect 16862 4613 16928 4647
rect 16862 4579 16878 4613
rect 16912 4579 16928 4613
rect 16862 4545 16928 4579
rect 16862 4511 16878 4545
rect 16912 4511 16928 4545
rect 16862 4477 16928 4511
rect 16862 4443 16878 4477
rect 16912 4443 16928 4477
rect 16862 4409 16928 4443
rect 16862 4375 16878 4409
rect 16912 4375 16928 4409
rect 16862 4341 16928 4375
rect 16862 4307 16878 4341
rect 16912 4307 16928 4341
rect 16862 4273 16928 4307
rect 16862 4239 16878 4273
rect 16912 4239 16928 4273
rect 16862 4205 16928 4239
rect 16862 4171 16878 4205
rect 16912 4171 16928 4205
rect 16862 4130 16928 4171
rect 16958 5089 17024 5130
rect 16958 5055 16974 5089
rect 17008 5055 17024 5089
rect 16958 5021 17024 5055
rect 16958 4987 16974 5021
rect 17008 4987 17024 5021
rect 16958 4953 17024 4987
rect 16958 4919 16974 4953
rect 17008 4919 17024 4953
rect 16958 4885 17024 4919
rect 16958 4851 16974 4885
rect 17008 4851 17024 4885
rect 16958 4817 17024 4851
rect 16958 4783 16974 4817
rect 17008 4783 17024 4817
rect 16958 4749 17024 4783
rect 16958 4715 16974 4749
rect 17008 4715 17024 4749
rect 16958 4681 17024 4715
rect 16958 4647 16974 4681
rect 17008 4647 17024 4681
rect 16958 4613 17024 4647
rect 16958 4579 16974 4613
rect 17008 4579 17024 4613
rect 16958 4545 17024 4579
rect 16958 4511 16974 4545
rect 17008 4511 17024 4545
rect 16958 4477 17024 4511
rect 16958 4443 16974 4477
rect 17008 4443 17024 4477
rect 16958 4409 17024 4443
rect 16958 4375 16974 4409
rect 17008 4375 17024 4409
rect 16958 4341 17024 4375
rect 16958 4307 16974 4341
rect 17008 4307 17024 4341
rect 16958 4273 17024 4307
rect 16958 4239 16974 4273
rect 17008 4239 17024 4273
rect 16958 4205 17024 4239
rect 16958 4171 16974 4205
rect 17008 4171 17024 4205
rect 16958 4130 17024 4171
rect 17054 5089 17120 5130
rect 17054 5055 17070 5089
rect 17104 5055 17120 5089
rect 17054 5021 17120 5055
rect 17054 4987 17070 5021
rect 17104 4987 17120 5021
rect 17054 4953 17120 4987
rect 17054 4919 17070 4953
rect 17104 4919 17120 4953
rect 17054 4885 17120 4919
rect 17054 4851 17070 4885
rect 17104 4851 17120 4885
rect 17054 4817 17120 4851
rect 17054 4783 17070 4817
rect 17104 4783 17120 4817
rect 17054 4749 17120 4783
rect 17054 4715 17070 4749
rect 17104 4715 17120 4749
rect 17054 4681 17120 4715
rect 17054 4647 17070 4681
rect 17104 4647 17120 4681
rect 17054 4613 17120 4647
rect 17054 4579 17070 4613
rect 17104 4579 17120 4613
rect 17054 4545 17120 4579
rect 17054 4511 17070 4545
rect 17104 4511 17120 4545
rect 17054 4477 17120 4511
rect 17054 4443 17070 4477
rect 17104 4443 17120 4477
rect 17054 4409 17120 4443
rect 17054 4375 17070 4409
rect 17104 4375 17120 4409
rect 17054 4341 17120 4375
rect 17054 4307 17070 4341
rect 17104 4307 17120 4341
rect 17054 4273 17120 4307
rect 17054 4239 17070 4273
rect 17104 4239 17120 4273
rect 17054 4205 17120 4239
rect 17054 4171 17070 4205
rect 17104 4171 17120 4205
rect 17054 4130 17120 4171
rect 17150 5089 17216 5130
rect 17150 5055 17166 5089
rect 17200 5055 17216 5089
rect 17150 5021 17216 5055
rect 17150 4987 17166 5021
rect 17200 4987 17216 5021
rect 17150 4953 17216 4987
rect 17150 4919 17166 4953
rect 17200 4919 17216 4953
rect 17150 4885 17216 4919
rect 17150 4851 17166 4885
rect 17200 4851 17216 4885
rect 17150 4817 17216 4851
rect 17150 4783 17166 4817
rect 17200 4783 17216 4817
rect 17150 4749 17216 4783
rect 17150 4715 17166 4749
rect 17200 4715 17216 4749
rect 17150 4681 17216 4715
rect 17150 4647 17166 4681
rect 17200 4647 17216 4681
rect 17150 4613 17216 4647
rect 17150 4579 17166 4613
rect 17200 4579 17216 4613
rect 17150 4545 17216 4579
rect 17150 4511 17166 4545
rect 17200 4511 17216 4545
rect 17150 4477 17216 4511
rect 17150 4443 17166 4477
rect 17200 4443 17216 4477
rect 17150 4409 17216 4443
rect 17150 4375 17166 4409
rect 17200 4375 17216 4409
rect 17150 4341 17216 4375
rect 17150 4307 17166 4341
rect 17200 4307 17216 4341
rect 17150 4273 17216 4307
rect 17150 4239 17166 4273
rect 17200 4239 17216 4273
rect 17150 4205 17216 4239
rect 17150 4171 17166 4205
rect 17200 4171 17216 4205
rect 17150 4130 17216 4171
rect 17246 5089 17308 5130
rect 17246 5055 17262 5089
rect 17296 5055 17308 5089
rect 17246 5021 17308 5055
rect 17246 4987 17262 5021
rect 17296 4987 17308 5021
rect 17246 4953 17308 4987
rect 17246 4919 17262 4953
rect 17296 4919 17308 4953
rect 17246 4885 17308 4919
rect 17246 4851 17262 4885
rect 17296 4851 17308 4885
rect 17246 4817 17308 4851
rect 17246 4783 17262 4817
rect 17296 4783 17308 4817
rect 17246 4749 17308 4783
rect 17246 4715 17262 4749
rect 17296 4715 17308 4749
rect 17246 4681 17308 4715
rect 17246 4647 17262 4681
rect 17296 4647 17308 4681
rect 17246 4613 17308 4647
rect 17246 4579 17262 4613
rect 17296 4579 17308 4613
rect 17246 4545 17308 4579
rect 17246 4511 17262 4545
rect 17296 4511 17308 4545
rect 17246 4477 17308 4511
rect 17246 4443 17262 4477
rect 17296 4443 17308 4477
rect 17246 4409 17308 4443
rect 17246 4375 17262 4409
rect 17296 4375 17308 4409
rect 17246 4341 17308 4375
rect 17246 4307 17262 4341
rect 17296 4307 17308 4341
rect 17246 4273 17308 4307
rect 17246 4239 17262 4273
rect 17296 4239 17308 4273
rect 17246 4205 17308 4239
rect 17246 4171 17262 4205
rect 17296 4171 17308 4205
rect 17246 4130 17308 4171
rect 17458 5087 17520 5128
rect 17458 5053 17470 5087
rect 17504 5053 17520 5087
rect 17458 5019 17520 5053
rect 17458 4985 17470 5019
rect 17504 4985 17520 5019
rect 17458 4951 17520 4985
rect 17458 4917 17470 4951
rect 17504 4917 17520 4951
rect 17458 4883 17520 4917
rect 17458 4849 17470 4883
rect 17504 4849 17520 4883
rect 17458 4815 17520 4849
rect 17458 4781 17470 4815
rect 17504 4781 17520 4815
rect 17458 4747 17520 4781
rect 17458 4713 17470 4747
rect 17504 4713 17520 4747
rect 17458 4679 17520 4713
rect 17458 4645 17470 4679
rect 17504 4645 17520 4679
rect 17458 4611 17520 4645
rect 17458 4577 17470 4611
rect 17504 4577 17520 4611
rect 17458 4543 17520 4577
rect 17458 4509 17470 4543
rect 17504 4509 17520 4543
rect 17458 4475 17520 4509
rect 17458 4441 17470 4475
rect 17504 4441 17520 4475
rect 17458 4407 17520 4441
rect 17458 4373 17470 4407
rect 17504 4373 17520 4407
rect 17458 4339 17520 4373
rect 17458 4305 17470 4339
rect 17504 4305 17520 4339
rect 17458 4271 17520 4305
rect 17458 4237 17470 4271
rect 17504 4237 17520 4271
rect 17458 4203 17520 4237
rect 17458 4169 17470 4203
rect 17504 4169 17520 4203
rect 15694 4093 15710 4127
rect 15744 4093 15756 4127
rect 15694 4059 15756 4093
rect 15694 4025 15710 4059
rect 15744 4025 15756 4059
rect 15694 3991 15756 4025
rect 15694 3957 15710 3991
rect 15744 3957 15756 3991
rect 17458 4128 17520 4169
rect 17550 5087 17616 5128
rect 17550 5053 17566 5087
rect 17600 5053 17616 5087
rect 17550 5019 17616 5053
rect 17550 4985 17566 5019
rect 17600 4985 17616 5019
rect 17550 4951 17616 4985
rect 17550 4917 17566 4951
rect 17600 4917 17616 4951
rect 17550 4883 17616 4917
rect 17550 4849 17566 4883
rect 17600 4849 17616 4883
rect 17550 4815 17616 4849
rect 17550 4781 17566 4815
rect 17600 4781 17616 4815
rect 17550 4747 17616 4781
rect 17550 4713 17566 4747
rect 17600 4713 17616 4747
rect 17550 4679 17616 4713
rect 17550 4645 17566 4679
rect 17600 4645 17616 4679
rect 17550 4611 17616 4645
rect 17550 4577 17566 4611
rect 17600 4577 17616 4611
rect 17550 4543 17616 4577
rect 17550 4509 17566 4543
rect 17600 4509 17616 4543
rect 17550 4475 17616 4509
rect 17550 4441 17566 4475
rect 17600 4441 17616 4475
rect 17550 4407 17616 4441
rect 17550 4373 17566 4407
rect 17600 4373 17616 4407
rect 17550 4339 17616 4373
rect 17550 4305 17566 4339
rect 17600 4305 17616 4339
rect 17550 4271 17616 4305
rect 17550 4237 17566 4271
rect 17600 4237 17616 4271
rect 17550 4203 17616 4237
rect 17550 4169 17566 4203
rect 17600 4169 17616 4203
rect 17550 4128 17616 4169
rect 17646 5087 17712 5128
rect 17646 5053 17662 5087
rect 17696 5053 17712 5087
rect 17646 5019 17712 5053
rect 17646 4985 17662 5019
rect 17696 4985 17712 5019
rect 17646 4951 17712 4985
rect 17646 4917 17662 4951
rect 17696 4917 17712 4951
rect 17646 4883 17712 4917
rect 17646 4849 17662 4883
rect 17696 4849 17712 4883
rect 17646 4815 17712 4849
rect 17646 4781 17662 4815
rect 17696 4781 17712 4815
rect 17646 4747 17712 4781
rect 17646 4713 17662 4747
rect 17696 4713 17712 4747
rect 17646 4679 17712 4713
rect 17646 4645 17662 4679
rect 17696 4645 17712 4679
rect 17646 4611 17712 4645
rect 17646 4577 17662 4611
rect 17696 4577 17712 4611
rect 17646 4543 17712 4577
rect 17646 4509 17662 4543
rect 17696 4509 17712 4543
rect 17646 4475 17712 4509
rect 17646 4441 17662 4475
rect 17696 4441 17712 4475
rect 17646 4407 17712 4441
rect 17646 4373 17662 4407
rect 17696 4373 17712 4407
rect 17646 4339 17712 4373
rect 17646 4305 17662 4339
rect 17696 4305 17712 4339
rect 17646 4271 17712 4305
rect 17646 4237 17662 4271
rect 17696 4237 17712 4271
rect 17646 4203 17712 4237
rect 17646 4169 17662 4203
rect 17696 4169 17712 4203
rect 17646 4128 17712 4169
rect 17742 5087 17808 5128
rect 17742 5053 17758 5087
rect 17792 5053 17808 5087
rect 17742 5019 17808 5053
rect 17742 4985 17758 5019
rect 17792 4985 17808 5019
rect 17742 4951 17808 4985
rect 17742 4917 17758 4951
rect 17792 4917 17808 4951
rect 17742 4883 17808 4917
rect 17742 4849 17758 4883
rect 17792 4849 17808 4883
rect 17742 4815 17808 4849
rect 17742 4781 17758 4815
rect 17792 4781 17808 4815
rect 17742 4747 17808 4781
rect 17742 4713 17758 4747
rect 17792 4713 17808 4747
rect 17742 4679 17808 4713
rect 17742 4645 17758 4679
rect 17792 4645 17808 4679
rect 17742 4611 17808 4645
rect 17742 4577 17758 4611
rect 17792 4577 17808 4611
rect 17742 4543 17808 4577
rect 17742 4509 17758 4543
rect 17792 4509 17808 4543
rect 17742 4475 17808 4509
rect 17742 4441 17758 4475
rect 17792 4441 17808 4475
rect 17742 4407 17808 4441
rect 17742 4373 17758 4407
rect 17792 4373 17808 4407
rect 17742 4339 17808 4373
rect 17742 4305 17758 4339
rect 17792 4305 17808 4339
rect 17742 4271 17808 4305
rect 17742 4237 17758 4271
rect 17792 4237 17808 4271
rect 17742 4203 17808 4237
rect 17742 4169 17758 4203
rect 17792 4169 17808 4203
rect 17742 4128 17808 4169
rect 17838 5087 17904 5128
rect 17838 5053 17854 5087
rect 17888 5053 17904 5087
rect 17838 5019 17904 5053
rect 17838 4985 17854 5019
rect 17888 4985 17904 5019
rect 17838 4951 17904 4985
rect 17838 4917 17854 4951
rect 17888 4917 17904 4951
rect 17838 4883 17904 4917
rect 17838 4849 17854 4883
rect 17888 4849 17904 4883
rect 17838 4815 17904 4849
rect 17838 4781 17854 4815
rect 17888 4781 17904 4815
rect 17838 4747 17904 4781
rect 17838 4713 17854 4747
rect 17888 4713 17904 4747
rect 17838 4679 17904 4713
rect 17838 4645 17854 4679
rect 17888 4645 17904 4679
rect 17838 4611 17904 4645
rect 17838 4577 17854 4611
rect 17888 4577 17904 4611
rect 17838 4543 17904 4577
rect 17838 4509 17854 4543
rect 17888 4509 17904 4543
rect 17838 4475 17904 4509
rect 17838 4441 17854 4475
rect 17888 4441 17904 4475
rect 17838 4407 17904 4441
rect 17838 4373 17854 4407
rect 17888 4373 17904 4407
rect 17838 4339 17904 4373
rect 17838 4305 17854 4339
rect 17888 4305 17904 4339
rect 17838 4271 17904 4305
rect 17838 4237 17854 4271
rect 17888 4237 17904 4271
rect 17838 4203 17904 4237
rect 17838 4169 17854 4203
rect 17888 4169 17904 4203
rect 17838 4128 17904 4169
rect 17934 5087 18000 5128
rect 17934 5053 17950 5087
rect 17984 5053 18000 5087
rect 17934 5019 18000 5053
rect 17934 4985 17950 5019
rect 17984 4985 18000 5019
rect 17934 4951 18000 4985
rect 17934 4917 17950 4951
rect 17984 4917 18000 4951
rect 17934 4883 18000 4917
rect 17934 4849 17950 4883
rect 17984 4849 18000 4883
rect 17934 4815 18000 4849
rect 17934 4781 17950 4815
rect 17984 4781 18000 4815
rect 17934 4747 18000 4781
rect 17934 4713 17950 4747
rect 17984 4713 18000 4747
rect 17934 4679 18000 4713
rect 17934 4645 17950 4679
rect 17984 4645 18000 4679
rect 17934 4611 18000 4645
rect 17934 4577 17950 4611
rect 17984 4577 18000 4611
rect 17934 4543 18000 4577
rect 17934 4509 17950 4543
rect 17984 4509 18000 4543
rect 17934 4475 18000 4509
rect 17934 4441 17950 4475
rect 17984 4441 18000 4475
rect 17934 4407 18000 4441
rect 17934 4373 17950 4407
rect 17984 4373 18000 4407
rect 17934 4339 18000 4373
rect 17934 4305 17950 4339
rect 17984 4305 18000 4339
rect 17934 4271 18000 4305
rect 17934 4237 17950 4271
rect 17984 4237 18000 4271
rect 17934 4203 18000 4237
rect 17934 4169 17950 4203
rect 17984 4169 18000 4203
rect 17934 4128 18000 4169
rect 18030 5087 18096 5128
rect 18030 5053 18046 5087
rect 18080 5053 18096 5087
rect 18030 5019 18096 5053
rect 18030 4985 18046 5019
rect 18080 4985 18096 5019
rect 18030 4951 18096 4985
rect 18030 4917 18046 4951
rect 18080 4917 18096 4951
rect 18030 4883 18096 4917
rect 18030 4849 18046 4883
rect 18080 4849 18096 4883
rect 18030 4815 18096 4849
rect 18030 4781 18046 4815
rect 18080 4781 18096 4815
rect 18030 4747 18096 4781
rect 18030 4713 18046 4747
rect 18080 4713 18096 4747
rect 18030 4679 18096 4713
rect 18030 4645 18046 4679
rect 18080 4645 18096 4679
rect 18030 4611 18096 4645
rect 18030 4577 18046 4611
rect 18080 4577 18096 4611
rect 18030 4543 18096 4577
rect 18030 4509 18046 4543
rect 18080 4509 18096 4543
rect 18030 4475 18096 4509
rect 18030 4441 18046 4475
rect 18080 4441 18096 4475
rect 18030 4407 18096 4441
rect 18030 4373 18046 4407
rect 18080 4373 18096 4407
rect 18030 4339 18096 4373
rect 18030 4305 18046 4339
rect 18080 4305 18096 4339
rect 18030 4271 18096 4305
rect 18030 4237 18046 4271
rect 18080 4237 18096 4271
rect 18030 4203 18096 4237
rect 18030 4169 18046 4203
rect 18080 4169 18096 4203
rect 18030 4128 18096 4169
rect 18126 5087 18192 5128
rect 18126 5053 18142 5087
rect 18176 5053 18192 5087
rect 18126 5019 18192 5053
rect 18126 4985 18142 5019
rect 18176 4985 18192 5019
rect 18126 4951 18192 4985
rect 18126 4917 18142 4951
rect 18176 4917 18192 4951
rect 18126 4883 18192 4917
rect 18126 4849 18142 4883
rect 18176 4849 18192 4883
rect 18126 4815 18192 4849
rect 18126 4781 18142 4815
rect 18176 4781 18192 4815
rect 18126 4747 18192 4781
rect 18126 4713 18142 4747
rect 18176 4713 18192 4747
rect 18126 4679 18192 4713
rect 18126 4645 18142 4679
rect 18176 4645 18192 4679
rect 18126 4611 18192 4645
rect 18126 4577 18142 4611
rect 18176 4577 18192 4611
rect 18126 4543 18192 4577
rect 18126 4509 18142 4543
rect 18176 4509 18192 4543
rect 18126 4475 18192 4509
rect 18126 4441 18142 4475
rect 18176 4441 18192 4475
rect 18126 4407 18192 4441
rect 18126 4373 18142 4407
rect 18176 4373 18192 4407
rect 18126 4339 18192 4373
rect 18126 4305 18142 4339
rect 18176 4305 18192 4339
rect 18126 4271 18192 4305
rect 18126 4237 18142 4271
rect 18176 4237 18192 4271
rect 18126 4203 18192 4237
rect 18126 4169 18142 4203
rect 18176 4169 18192 4203
rect 18126 4128 18192 4169
rect 18222 5087 18288 5128
rect 18222 5053 18238 5087
rect 18272 5053 18288 5087
rect 18222 5019 18288 5053
rect 18222 4985 18238 5019
rect 18272 4985 18288 5019
rect 18222 4951 18288 4985
rect 18222 4917 18238 4951
rect 18272 4917 18288 4951
rect 18222 4883 18288 4917
rect 18222 4849 18238 4883
rect 18272 4849 18288 4883
rect 18222 4815 18288 4849
rect 18222 4781 18238 4815
rect 18272 4781 18288 4815
rect 18222 4747 18288 4781
rect 18222 4713 18238 4747
rect 18272 4713 18288 4747
rect 18222 4679 18288 4713
rect 18222 4645 18238 4679
rect 18272 4645 18288 4679
rect 18222 4611 18288 4645
rect 18222 4577 18238 4611
rect 18272 4577 18288 4611
rect 18222 4543 18288 4577
rect 18222 4509 18238 4543
rect 18272 4509 18288 4543
rect 18222 4475 18288 4509
rect 18222 4441 18238 4475
rect 18272 4441 18288 4475
rect 18222 4407 18288 4441
rect 18222 4373 18238 4407
rect 18272 4373 18288 4407
rect 18222 4339 18288 4373
rect 18222 4305 18238 4339
rect 18272 4305 18288 4339
rect 18222 4271 18288 4305
rect 18222 4237 18238 4271
rect 18272 4237 18288 4271
rect 18222 4203 18288 4237
rect 18222 4169 18238 4203
rect 18272 4169 18288 4203
rect 18222 4128 18288 4169
rect 18318 5087 18384 5128
rect 18318 5053 18334 5087
rect 18368 5053 18384 5087
rect 18318 5019 18384 5053
rect 18318 4985 18334 5019
rect 18368 4985 18384 5019
rect 18318 4951 18384 4985
rect 18318 4917 18334 4951
rect 18368 4917 18384 4951
rect 18318 4883 18384 4917
rect 18318 4849 18334 4883
rect 18368 4849 18384 4883
rect 18318 4815 18384 4849
rect 18318 4781 18334 4815
rect 18368 4781 18384 4815
rect 18318 4747 18384 4781
rect 18318 4713 18334 4747
rect 18368 4713 18384 4747
rect 18318 4679 18384 4713
rect 18318 4645 18334 4679
rect 18368 4645 18384 4679
rect 18318 4611 18384 4645
rect 18318 4577 18334 4611
rect 18368 4577 18384 4611
rect 18318 4543 18384 4577
rect 18318 4509 18334 4543
rect 18368 4509 18384 4543
rect 18318 4475 18384 4509
rect 18318 4441 18334 4475
rect 18368 4441 18384 4475
rect 18318 4407 18384 4441
rect 18318 4373 18334 4407
rect 18368 4373 18384 4407
rect 18318 4339 18384 4373
rect 18318 4305 18334 4339
rect 18368 4305 18384 4339
rect 18318 4271 18384 4305
rect 18318 4237 18334 4271
rect 18368 4237 18384 4271
rect 18318 4203 18384 4237
rect 18318 4169 18334 4203
rect 18368 4169 18384 4203
rect 18318 4128 18384 4169
rect 18414 5087 18476 5128
rect 18414 5053 18430 5087
rect 18464 5053 18476 5087
rect 18414 5019 18476 5053
rect 18414 4985 18430 5019
rect 18464 4985 18476 5019
rect 18414 4951 18476 4985
rect 18414 4917 18430 4951
rect 18464 4917 18476 4951
rect 18414 4883 18476 4917
rect 18414 4849 18430 4883
rect 18464 4849 18476 4883
rect 18414 4815 18476 4849
rect 18414 4781 18430 4815
rect 18464 4781 18476 4815
rect 18414 4747 18476 4781
rect 18414 4713 18430 4747
rect 18464 4713 18476 4747
rect 18414 4679 18476 4713
rect 18414 4645 18430 4679
rect 18464 4645 18476 4679
rect 18414 4611 18476 4645
rect 18414 4577 18430 4611
rect 18464 4577 18476 4611
rect 18414 4543 18476 4577
rect 18414 4509 18430 4543
rect 18464 4509 18476 4543
rect 18414 4475 18476 4509
rect 18414 4441 18430 4475
rect 18464 4441 18476 4475
rect 18414 4407 18476 4441
rect 18414 4373 18430 4407
rect 18464 4373 18476 4407
rect 18414 4339 18476 4373
rect 18414 4305 18430 4339
rect 18464 4305 18476 4339
rect 18414 4271 18476 4305
rect 18414 4237 18430 4271
rect 18464 4237 18476 4271
rect 18414 4203 18476 4237
rect 18414 4169 18430 4203
rect 18464 4169 18476 4203
rect 18414 4128 18476 4169
rect 18662 5081 18724 5122
rect 18662 5047 18674 5081
rect 18708 5047 18724 5081
rect 18662 5013 18724 5047
rect 18662 4979 18674 5013
rect 18708 4979 18724 5013
rect 18662 4945 18724 4979
rect 18662 4911 18674 4945
rect 18708 4911 18724 4945
rect 18662 4877 18724 4911
rect 18662 4843 18674 4877
rect 18708 4843 18724 4877
rect 18662 4809 18724 4843
rect 18662 4775 18674 4809
rect 18708 4775 18724 4809
rect 18662 4741 18724 4775
rect 18662 4707 18674 4741
rect 18708 4707 18724 4741
rect 18662 4673 18724 4707
rect 18662 4639 18674 4673
rect 18708 4639 18724 4673
rect 18662 4605 18724 4639
rect 18662 4571 18674 4605
rect 18708 4571 18724 4605
rect 18662 4537 18724 4571
rect 18662 4503 18674 4537
rect 18708 4503 18724 4537
rect 18662 4469 18724 4503
rect 18662 4435 18674 4469
rect 18708 4435 18724 4469
rect 18662 4401 18724 4435
rect 18662 4367 18674 4401
rect 18708 4367 18724 4401
rect 18662 4333 18724 4367
rect 18662 4299 18674 4333
rect 18708 4299 18724 4333
rect 18662 4265 18724 4299
rect 18662 4231 18674 4265
rect 18708 4231 18724 4265
rect 18662 4197 18724 4231
rect 18662 4163 18674 4197
rect 18708 4163 18724 4197
rect 18662 4122 18724 4163
rect 18754 5081 18820 5122
rect 18754 5047 18770 5081
rect 18804 5047 18820 5081
rect 18754 5013 18820 5047
rect 18754 4979 18770 5013
rect 18804 4979 18820 5013
rect 18754 4945 18820 4979
rect 18754 4911 18770 4945
rect 18804 4911 18820 4945
rect 18754 4877 18820 4911
rect 18754 4843 18770 4877
rect 18804 4843 18820 4877
rect 18754 4809 18820 4843
rect 18754 4775 18770 4809
rect 18804 4775 18820 4809
rect 18754 4741 18820 4775
rect 18754 4707 18770 4741
rect 18804 4707 18820 4741
rect 18754 4673 18820 4707
rect 18754 4639 18770 4673
rect 18804 4639 18820 4673
rect 18754 4605 18820 4639
rect 18754 4571 18770 4605
rect 18804 4571 18820 4605
rect 18754 4537 18820 4571
rect 18754 4503 18770 4537
rect 18804 4503 18820 4537
rect 18754 4469 18820 4503
rect 18754 4435 18770 4469
rect 18804 4435 18820 4469
rect 18754 4401 18820 4435
rect 18754 4367 18770 4401
rect 18804 4367 18820 4401
rect 18754 4333 18820 4367
rect 18754 4299 18770 4333
rect 18804 4299 18820 4333
rect 18754 4265 18820 4299
rect 18754 4231 18770 4265
rect 18804 4231 18820 4265
rect 18754 4197 18820 4231
rect 18754 4163 18770 4197
rect 18804 4163 18820 4197
rect 18754 4122 18820 4163
rect 18850 5081 18916 5122
rect 18850 5047 18866 5081
rect 18900 5047 18916 5081
rect 18850 5013 18916 5047
rect 18850 4979 18866 5013
rect 18900 4979 18916 5013
rect 18850 4945 18916 4979
rect 18850 4911 18866 4945
rect 18900 4911 18916 4945
rect 18850 4877 18916 4911
rect 18850 4843 18866 4877
rect 18900 4843 18916 4877
rect 18850 4809 18916 4843
rect 18850 4775 18866 4809
rect 18900 4775 18916 4809
rect 18850 4741 18916 4775
rect 18850 4707 18866 4741
rect 18900 4707 18916 4741
rect 18850 4673 18916 4707
rect 18850 4639 18866 4673
rect 18900 4639 18916 4673
rect 18850 4605 18916 4639
rect 18850 4571 18866 4605
rect 18900 4571 18916 4605
rect 18850 4537 18916 4571
rect 18850 4503 18866 4537
rect 18900 4503 18916 4537
rect 18850 4469 18916 4503
rect 18850 4435 18866 4469
rect 18900 4435 18916 4469
rect 18850 4401 18916 4435
rect 18850 4367 18866 4401
rect 18900 4367 18916 4401
rect 18850 4333 18916 4367
rect 18850 4299 18866 4333
rect 18900 4299 18916 4333
rect 18850 4265 18916 4299
rect 18850 4231 18866 4265
rect 18900 4231 18916 4265
rect 18850 4197 18916 4231
rect 18850 4163 18866 4197
rect 18900 4163 18916 4197
rect 18850 4122 18916 4163
rect 18946 5081 19012 5122
rect 18946 5047 18962 5081
rect 18996 5047 19012 5081
rect 18946 5013 19012 5047
rect 18946 4979 18962 5013
rect 18996 4979 19012 5013
rect 18946 4945 19012 4979
rect 18946 4911 18962 4945
rect 18996 4911 19012 4945
rect 18946 4877 19012 4911
rect 18946 4843 18962 4877
rect 18996 4843 19012 4877
rect 18946 4809 19012 4843
rect 18946 4775 18962 4809
rect 18996 4775 19012 4809
rect 18946 4741 19012 4775
rect 18946 4707 18962 4741
rect 18996 4707 19012 4741
rect 18946 4673 19012 4707
rect 18946 4639 18962 4673
rect 18996 4639 19012 4673
rect 18946 4605 19012 4639
rect 18946 4571 18962 4605
rect 18996 4571 19012 4605
rect 18946 4537 19012 4571
rect 18946 4503 18962 4537
rect 18996 4503 19012 4537
rect 18946 4469 19012 4503
rect 18946 4435 18962 4469
rect 18996 4435 19012 4469
rect 18946 4401 19012 4435
rect 18946 4367 18962 4401
rect 18996 4367 19012 4401
rect 18946 4333 19012 4367
rect 18946 4299 18962 4333
rect 18996 4299 19012 4333
rect 18946 4265 19012 4299
rect 18946 4231 18962 4265
rect 18996 4231 19012 4265
rect 18946 4197 19012 4231
rect 18946 4163 18962 4197
rect 18996 4163 19012 4197
rect 18946 4122 19012 4163
rect 19042 5081 19108 5122
rect 19042 5047 19058 5081
rect 19092 5047 19108 5081
rect 19042 5013 19108 5047
rect 19042 4979 19058 5013
rect 19092 4979 19108 5013
rect 19042 4945 19108 4979
rect 19042 4911 19058 4945
rect 19092 4911 19108 4945
rect 19042 4877 19108 4911
rect 19042 4843 19058 4877
rect 19092 4843 19108 4877
rect 19042 4809 19108 4843
rect 19042 4775 19058 4809
rect 19092 4775 19108 4809
rect 19042 4741 19108 4775
rect 19042 4707 19058 4741
rect 19092 4707 19108 4741
rect 19042 4673 19108 4707
rect 19042 4639 19058 4673
rect 19092 4639 19108 4673
rect 19042 4605 19108 4639
rect 19042 4571 19058 4605
rect 19092 4571 19108 4605
rect 19042 4537 19108 4571
rect 19042 4503 19058 4537
rect 19092 4503 19108 4537
rect 19042 4469 19108 4503
rect 19042 4435 19058 4469
rect 19092 4435 19108 4469
rect 19042 4401 19108 4435
rect 19042 4367 19058 4401
rect 19092 4367 19108 4401
rect 19042 4333 19108 4367
rect 19042 4299 19058 4333
rect 19092 4299 19108 4333
rect 19042 4265 19108 4299
rect 19042 4231 19058 4265
rect 19092 4231 19108 4265
rect 19042 4197 19108 4231
rect 19042 4163 19058 4197
rect 19092 4163 19108 4197
rect 19042 4122 19108 4163
rect 19138 5081 19204 5122
rect 19138 5047 19154 5081
rect 19188 5047 19204 5081
rect 19138 5013 19204 5047
rect 19138 4979 19154 5013
rect 19188 4979 19204 5013
rect 19138 4945 19204 4979
rect 19138 4911 19154 4945
rect 19188 4911 19204 4945
rect 19138 4877 19204 4911
rect 19138 4843 19154 4877
rect 19188 4843 19204 4877
rect 19138 4809 19204 4843
rect 19138 4775 19154 4809
rect 19188 4775 19204 4809
rect 19138 4741 19204 4775
rect 19138 4707 19154 4741
rect 19188 4707 19204 4741
rect 19138 4673 19204 4707
rect 19138 4639 19154 4673
rect 19188 4639 19204 4673
rect 19138 4605 19204 4639
rect 19138 4571 19154 4605
rect 19188 4571 19204 4605
rect 19138 4537 19204 4571
rect 19138 4503 19154 4537
rect 19188 4503 19204 4537
rect 19138 4469 19204 4503
rect 19138 4435 19154 4469
rect 19188 4435 19204 4469
rect 19138 4401 19204 4435
rect 19138 4367 19154 4401
rect 19188 4367 19204 4401
rect 19138 4333 19204 4367
rect 19138 4299 19154 4333
rect 19188 4299 19204 4333
rect 19138 4265 19204 4299
rect 19138 4231 19154 4265
rect 19188 4231 19204 4265
rect 19138 4197 19204 4231
rect 19138 4163 19154 4197
rect 19188 4163 19204 4197
rect 19138 4122 19204 4163
rect 19234 5081 19300 5122
rect 19234 5047 19250 5081
rect 19284 5047 19300 5081
rect 19234 5013 19300 5047
rect 19234 4979 19250 5013
rect 19284 4979 19300 5013
rect 19234 4945 19300 4979
rect 19234 4911 19250 4945
rect 19284 4911 19300 4945
rect 19234 4877 19300 4911
rect 19234 4843 19250 4877
rect 19284 4843 19300 4877
rect 19234 4809 19300 4843
rect 19234 4775 19250 4809
rect 19284 4775 19300 4809
rect 19234 4741 19300 4775
rect 19234 4707 19250 4741
rect 19284 4707 19300 4741
rect 19234 4673 19300 4707
rect 19234 4639 19250 4673
rect 19284 4639 19300 4673
rect 19234 4605 19300 4639
rect 19234 4571 19250 4605
rect 19284 4571 19300 4605
rect 19234 4537 19300 4571
rect 19234 4503 19250 4537
rect 19284 4503 19300 4537
rect 19234 4469 19300 4503
rect 19234 4435 19250 4469
rect 19284 4435 19300 4469
rect 19234 4401 19300 4435
rect 19234 4367 19250 4401
rect 19284 4367 19300 4401
rect 19234 4333 19300 4367
rect 19234 4299 19250 4333
rect 19284 4299 19300 4333
rect 19234 4265 19300 4299
rect 19234 4231 19250 4265
rect 19284 4231 19300 4265
rect 19234 4197 19300 4231
rect 19234 4163 19250 4197
rect 19284 4163 19300 4197
rect 19234 4122 19300 4163
rect 19330 5081 19396 5122
rect 19330 5047 19346 5081
rect 19380 5047 19396 5081
rect 19330 5013 19396 5047
rect 19330 4979 19346 5013
rect 19380 4979 19396 5013
rect 19330 4945 19396 4979
rect 19330 4911 19346 4945
rect 19380 4911 19396 4945
rect 19330 4877 19396 4911
rect 19330 4843 19346 4877
rect 19380 4843 19396 4877
rect 19330 4809 19396 4843
rect 19330 4775 19346 4809
rect 19380 4775 19396 4809
rect 19330 4741 19396 4775
rect 19330 4707 19346 4741
rect 19380 4707 19396 4741
rect 19330 4673 19396 4707
rect 19330 4639 19346 4673
rect 19380 4639 19396 4673
rect 19330 4605 19396 4639
rect 19330 4571 19346 4605
rect 19380 4571 19396 4605
rect 19330 4537 19396 4571
rect 19330 4503 19346 4537
rect 19380 4503 19396 4537
rect 19330 4469 19396 4503
rect 19330 4435 19346 4469
rect 19380 4435 19396 4469
rect 19330 4401 19396 4435
rect 19330 4367 19346 4401
rect 19380 4367 19396 4401
rect 19330 4333 19396 4367
rect 19330 4299 19346 4333
rect 19380 4299 19396 4333
rect 19330 4265 19396 4299
rect 19330 4231 19346 4265
rect 19380 4231 19396 4265
rect 19330 4197 19396 4231
rect 19330 4163 19346 4197
rect 19380 4163 19396 4197
rect 19330 4122 19396 4163
rect 19426 5081 19492 5122
rect 19426 5047 19442 5081
rect 19476 5047 19492 5081
rect 19426 5013 19492 5047
rect 19426 4979 19442 5013
rect 19476 4979 19492 5013
rect 19426 4945 19492 4979
rect 19426 4911 19442 4945
rect 19476 4911 19492 4945
rect 19426 4877 19492 4911
rect 19426 4843 19442 4877
rect 19476 4843 19492 4877
rect 19426 4809 19492 4843
rect 19426 4775 19442 4809
rect 19476 4775 19492 4809
rect 19426 4741 19492 4775
rect 19426 4707 19442 4741
rect 19476 4707 19492 4741
rect 19426 4673 19492 4707
rect 19426 4639 19442 4673
rect 19476 4639 19492 4673
rect 19426 4605 19492 4639
rect 19426 4571 19442 4605
rect 19476 4571 19492 4605
rect 19426 4537 19492 4571
rect 19426 4503 19442 4537
rect 19476 4503 19492 4537
rect 19426 4469 19492 4503
rect 19426 4435 19442 4469
rect 19476 4435 19492 4469
rect 19426 4401 19492 4435
rect 19426 4367 19442 4401
rect 19476 4367 19492 4401
rect 19426 4333 19492 4367
rect 19426 4299 19442 4333
rect 19476 4299 19492 4333
rect 19426 4265 19492 4299
rect 19426 4231 19442 4265
rect 19476 4231 19492 4265
rect 19426 4197 19492 4231
rect 19426 4163 19442 4197
rect 19476 4163 19492 4197
rect 19426 4122 19492 4163
rect 19522 5081 19588 5122
rect 19522 5047 19538 5081
rect 19572 5047 19588 5081
rect 19522 5013 19588 5047
rect 19522 4979 19538 5013
rect 19572 4979 19588 5013
rect 19522 4945 19588 4979
rect 19522 4911 19538 4945
rect 19572 4911 19588 4945
rect 19522 4877 19588 4911
rect 19522 4843 19538 4877
rect 19572 4843 19588 4877
rect 19522 4809 19588 4843
rect 19522 4775 19538 4809
rect 19572 4775 19588 4809
rect 19522 4741 19588 4775
rect 19522 4707 19538 4741
rect 19572 4707 19588 4741
rect 19522 4673 19588 4707
rect 19522 4639 19538 4673
rect 19572 4639 19588 4673
rect 19522 4605 19588 4639
rect 19522 4571 19538 4605
rect 19572 4571 19588 4605
rect 19522 4537 19588 4571
rect 19522 4503 19538 4537
rect 19572 4503 19588 4537
rect 19522 4469 19588 4503
rect 19522 4435 19538 4469
rect 19572 4435 19588 4469
rect 19522 4401 19588 4435
rect 19522 4367 19538 4401
rect 19572 4367 19588 4401
rect 19522 4333 19588 4367
rect 19522 4299 19538 4333
rect 19572 4299 19588 4333
rect 19522 4265 19588 4299
rect 19522 4231 19538 4265
rect 19572 4231 19588 4265
rect 19522 4197 19588 4231
rect 19522 4163 19538 4197
rect 19572 4163 19588 4197
rect 19522 4122 19588 4163
rect 19618 5081 19684 5122
rect 19618 5047 19634 5081
rect 19668 5047 19684 5081
rect 19618 5013 19684 5047
rect 19618 4979 19634 5013
rect 19668 4979 19684 5013
rect 19618 4945 19684 4979
rect 19618 4911 19634 4945
rect 19668 4911 19684 4945
rect 19618 4877 19684 4911
rect 19618 4843 19634 4877
rect 19668 4843 19684 4877
rect 19618 4809 19684 4843
rect 19618 4775 19634 4809
rect 19668 4775 19684 4809
rect 19618 4741 19684 4775
rect 19618 4707 19634 4741
rect 19668 4707 19684 4741
rect 19618 4673 19684 4707
rect 19618 4639 19634 4673
rect 19668 4639 19684 4673
rect 19618 4605 19684 4639
rect 19618 4571 19634 4605
rect 19668 4571 19684 4605
rect 19618 4537 19684 4571
rect 19618 4503 19634 4537
rect 19668 4503 19684 4537
rect 19618 4469 19684 4503
rect 19618 4435 19634 4469
rect 19668 4435 19684 4469
rect 19618 4401 19684 4435
rect 19618 4367 19634 4401
rect 19668 4367 19684 4401
rect 19618 4333 19684 4367
rect 19618 4299 19634 4333
rect 19668 4299 19684 4333
rect 19618 4265 19684 4299
rect 19618 4231 19634 4265
rect 19668 4231 19684 4265
rect 19618 4197 19684 4231
rect 19618 4163 19634 4197
rect 19668 4163 19684 4197
rect 19618 4122 19684 4163
rect 19714 5081 19780 5122
rect 19714 5047 19730 5081
rect 19764 5047 19780 5081
rect 19714 5013 19780 5047
rect 19714 4979 19730 5013
rect 19764 4979 19780 5013
rect 19714 4945 19780 4979
rect 19714 4911 19730 4945
rect 19764 4911 19780 4945
rect 19714 4877 19780 4911
rect 19714 4843 19730 4877
rect 19764 4843 19780 4877
rect 19714 4809 19780 4843
rect 19714 4775 19730 4809
rect 19764 4775 19780 4809
rect 19714 4741 19780 4775
rect 19714 4707 19730 4741
rect 19764 4707 19780 4741
rect 19714 4673 19780 4707
rect 19714 4639 19730 4673
rect 19764 4639 19780 4673
rect 19714 4605 19780 4639
rect 19714 4571 19730 4605
rect 19764 4571 19780 4605
rect 19714 4537 19780 4571
rect 19714 4503 19730 4537
rect 19764 4503 19780 4537
rect 19714 4469 19780 4503
rect 19714 4435 19730 4469
rect 19764 4435 19780 4469
rect 19714 4401 19780 4435
rect 19714 4367 19730 4401
rect 19764 4367 19780 4401
rect 19714 4333 19780 4367
rect 19714 4299 19730 4333
rect 19764 4299 19780 4333
rect 19714 4265 19780 4299
rect 19714 4231 19730 4265
rect 19764 4231 19780 4265
rect 19714 4197 19780 4231
rect 19714 4163 19730 4197
rect 19764 4163 19780 4197
rect 19714 4122 19780 4163
rect 19810 5081 19876 5122
rect 19810 5047 19826 5081
rect 19860 5047 19876 5081
rect 19810 5013 19876 5047
rect 19810 4979 19826 5013
rect 19860 4979 19876 5013
rect 19810 4945 19876 4979
rect 19810 4911 19826 4945
rect 19860 4911 19876 4945
rect 19810 4877 19876 4911
rect 19810 4843 19826 4877
rect 19860 4843 19876 4877
rect 19810 4809 19876 4843
rect 19810 4775 19826 4809
rect 19860 4775 19876 4809
rect 19810 4741 19876 4775
rect 19810 4707 19826 4741
rect 19860 4707 19876 4741
rect 19810 4673 19876 4707
rect 19810 4639 19826 4673
rect 19860 4639 19876 4673
rect 19810 4605 19876 4639
rect 19810 4571 19826 4605
rect 19860 4571 19876 4605
rect 19810 4537 19876 4571
rect 19810 4503 19826 4537
rect 19860 4503 19876 4537
rect 19810 4469 19876 4503
rect 19810 4435 19826 4469
rect 19860 4435 19876 4469
rect 19810 4401 19876 4435
rect 19810 4367 19826 4401
rect 19860 4367 19876 4401
rect 19810 4333 19876 4367
rect 19810 4299 19826 4333
rect 19860 4299 19876 4333
rect 19810 4265 19876 4299
rect 19810 4231 19826 4265
rect 19860 4231 19876 4265
rect 19810 4197 19876 4231
rect 19810 4163 19826 4197
rect 19860 4163 19876 4197
rect 19810 4122 19876 4163
rect 19906 5081 19972 5122
rect 19906 5047 19922 5081
rect 19956 5047 19972 5081
rect 19906 5013 19972 5047
rect 19906 4979 19922 5013
rect 19956 4979 19972 5013
rect 19906 4945 19972 4979
rect 19906 4911 19922 4945
rect 19956 4911 19972 4945
rect 19906 4877 19972 4911
rect 19906 4843 19922 4877
rect 19956 4843 19972 4877
rect 19906 4809 19972 4843
rect 19906 4775 19922 4809
rect 19956 4775 19972 4809
rect 19906 4741 19972 4775
rect 19906 4707 19922 4741
rect 19956 4707 19972 4741
rect 19906 4673 19972 4707
rect 19906 4639 19922 4673
rect 19956 4639 19972 4673
rect 19906 4605 19972 4639
rect 19906 4571 19922 4605
rect 19956 4571 19972 4605
rect 19906 4537 19972 4571
rect 19906 4503 19922 4537
rect 19956 4503 19972 4537
rect 19906 4469 19972 4503
rect 19906 4435 19922 4469
rect 19956 4435 19972 4469
rect 19906 4401 19972 4435
rect 19906 4367 19922 4401
rect 19956 4367 19972 4401
rect 19906 4333 19972 4367
rect 19906 4299 19922 4333
rect 19956 4299 19972 4333
rect 19906 4265 19972 4299
rect 19906 4231 19922 4265
rect 19956 4231 19972 4265
rect 19906 4197 19972 4231
rect 19906 4163 19922 4197
rect 19956 4163 19972 4197
rect 19906 4122 19972 4163
rect 20002 5081 20068 5122
rect 20002 5047 20018 5081
rect 20052 5047 20068 5081
rect 20002 5013 20068 5047
rect 20002 4979 20018 5013
rect 20052 4979 20068 5013
rect 20002 4945 20068 4979
rect 20002 4911 20018 4945
rect 20052 4911 20068 4945
rect 20002 4877 20068 4911
rect 20002 4843 20018 4877
rect 20052 4843 20068 4877
rect 20002 4809 20068 4843
rect 20002 4775 20018 4809
rect 20052 4775 20068 4809
rect 20002 4741 20068 4775
rect 20002 4707 20018 4741
rect 20052 4707 20068 4741
rect 20002 4673 20068 4707
rect 20002 4639 20018 4673
rect 20052 4639 20068 4673
rect 20002 4605 20068 4639
rect 20002 4571 20018 4605
rect 20052 4571 20068 4605
rect 20002 4537 20068 4571
rect 20002 4503 20018 4537
rect 20052 4503 20068 4537
rect 20002 4469 20068 4503
rect 20002 4435 20018 4469
rect 20052 4435 20068 4469
rect 20002 4401 20068 4435
rect 20002 4367 20018 4401
rect 20052 4367 20068 4401
rect 20002 4333 20068 4367
rect 20002 4299 20018 4333
rect 20052 4299 20068 4333
rect 20002 4265 20068 4299
rect 20002 4231 20018 4265
rect 20052 4231 20068 4265
rect 20002 4197 20068 4231
rect 20002 4163 20018 4197
rect 20052 4163 20068 4197
rect 20002 4122 20068 4163
rect 20098 5081 20160 5122
rect 20098 5047 20114 5081
rect 20148 5047 20160 5081
rect 20098 5013 20160 5047
rect 20098 4979 20114 5013
rect 20148 4979 20160 5013
rect 20098 4945 20160 4979
rect 20098 4911 20114 4945
rect 20148 4911 20160 4945
rect 20098 4877 20160 4911
rect 20098 4843 20114 4877
rect 20148 4843 20160 4877
rect 20098 4809 20160 4843
rect 20098 4775 20114 4809
rect 20148 4775 20160 4809
rect 20098 4741 20160 4775
rect 20098 4707 20114 4741
rect 20148 4707 20160 4741
rect 20098 4673 20160 4707
rect 20098 4639 20114 4673
rect 20148 4639 20160 4673
rect 20098 4605 20160 4639
rect 20098 4571 20114 4605
rect 20148 4571 20160 4605
rect 20098 4537 20160 4571
rect 20098 4503 20114 4537
rect 20148 4503 20160 4537
rect 20098 4469 20160 4503
rect 20098 4435 20114 4469
rect 20148 4435 20160 4469
rect 20098 4401 20160 4435
rect 20098 4367 20114 4401
rect 20148 4367 20160 4401
rect 20098 4333 20160 4367
rect 20098 4299 20114 4333
rect 20148 4299 20160 4333
rect 20098 4265 20160 4299
rect 20098 4231 20114 4265
rect 20148 4231 20160 4265
rect 20098 4197 20160 4231
rect 20098 4163 20114 4197
rect 20148 4163 20160 4197
rect 20098 4122 20160 4163
rect 20326 5075 20388 5116
rect 20326 5041 20338 5075
rect 20372 5041 20388 5075
rect 20326 5007 20388 5041
rect 20326 4973 20338 5007
rect 20372 4973 20388 5007
rect 20326 4939 20388 4973
rect 20326 4905 20338 4939
rect 20372 4905 20388 4939
rect 20326 4871 20388 4905
rect 20326 4837 20338 4871
rect 20372 4837 20388 4871
rect 20326 4803 20388 4837
rect 20326 4769 20338 4803
rect 20372 4769 20388 4803
rect 20326 4735 20388 4769
rect 20326 4701 20338 4735
rect 20372 4701 20388 4735
rect 20326 4667 20388 4701
rect 20326 4633 20338 4667
rect 20372 4633 20388 4667
rect 20326 4599 20388 4633
rect 20326 4565 20338 4599
rect 20372 4565 20388 4599
rect 20326 4531 20388 4565
rect 20326 4497 20338 4531
rect 20372 4497 20388 4531
rect 20326 4463 20388 4497
rect 20326 4429 20338 4463
rect 20372 4429 20388 4463
rect 20326 4395 20388 4429
rect 20326 4361 20338 4395
rect 20372 4361 20388 4395
rect 20326 4327 20388 4361
rect 20326 4293 20338 4327
rect 20372 4293 20388 4327
rect 20326 4259 20388 4293
rect 20326 4225 20338 4259
rect 20372 4225 20388 4259
rect 20326 4191 20388 4225
rect 20326 4157 20338 4191
rect 20372 4157 20388 4191
rect 20326 4116 20388 4157
rect 20418 5075 20484 5116
rect 20418 5041 20434 5075
rect 20468 5041 20484 5075
rect 20418 5007 20484 5041
rect 20418 4973 20434 5007
rect 20468 4973 20484 5007
rect 20418 4939 20484 4973
rect 20418 4905 20434 4939
rect 20468 4905 20484 4939
rect 20418 4871 20484 4905
rect 20418 4837 20434 4871
rect 20468 4837 20484 4871
rect 20418 4803 20484 4837
rect 20418 4769 20434 4803
rect 20468 4769 20484 4803
rect 20418 4735 20484 4769
rect 20418 4701 20434 4735
rect 20468 4701 20484 4735
rect 20418 4667 20484 4701
rect 20418 4633 20434 4667
rect 20468 4633 20484 4667
rect 20418 4599 20484 4633
rect 20418 4565 20434 4599
rect 20468 4565 20484 4599
rect 20418 4531 20484 4565
rect 20418 4497 20434 4531
rect 20468 4497 20484 4531
rect 20418 4463 20484 4497
rect 20418 4429 20434 4463
rect 20468 4429 20484 4463
rect 20418 4395 20484 4429
rect 20418 4361 20434 4395
rect 20468 4361 20484 4395
rect 20418 4327 20484 4361
rect 20418 4293 20434 4327
rect 20468 4293 20484 4327
rect 20418 4259 20484 4293
rect 20418 4225 20434 4259
rect 20468 4225 20484 4259
rect 20418 4191 20484 4225
rect 20418 4157 20434 4191
rect 20468 4157 20484 4191
rect 20418 4116 20484 4157
rect 20514 5075 20580 5116
rect 20514 5041 20530 5075
rect 20564 5041 20580 5075
rect 20514 5007 20580 5041
rect 20514 4973 20530 5007
rect 20564 4973 20580 5007
rect 20514 4939 20580 4973
rect 20514 4905 20530 4939
rect 20564 4905 20580 4939
rect 20514 4871 20580 4905
rect 20514 4837 20530 4871
rect 20564 4837 20580 4871
rect 20514 4803 20580 4837
rect 20514 4769 20530 4803
rect 20564 4769 20580 4803
rect 20514 4735 20580 4769
rect 20514 4701 20530 4735
rect 20564 4701 20580 4735
rect 20514 4667 20580 4701
rect 20514 4633 20530 4667
rect 20564 4633 20580 4667
rect 20514 4599 20580 4633
rect 20514 4565 20530 4599
rect 20564 4565 20580 4599
rect 20514 4531 20580 4565
rect 20514 4497 20530 4531
rect 20564 4497 20580 4531
rect 20514 4463 20580 4497
rect 20514 4429 20530 4463
rect 20564 4429 20580 4463
rect 20514 4395 20580 4429
rect 20514 4361 20530 4395
rect 20564 4361 20580 4395
rect 20514 4327 20580 4361
rect 20514 4293 20530 4327
rect 20564 4293 20580 4327
rect 20514 4259 20580 4293
rect 20514 4225 20530 4259
rect 20564 4225 20580 4259
rect 20514 4191 20580 4225
rect 20514 4157 20530 4191
rect 20564 4157 20580 4191
rect 20514 4116 20580 4157
rect 20610 5075 20676 5116
rect 20610 5041 20626 5075
rect 20660 5041 20676 5075
rect 20610 5007 20676 5041
rect 20610 4973 20626 5007
rect 20660 4973 20676 5007
rect 20610 4939 20676 4973
rect 20610 4905 20626 4939
rect 20660 4905 20676 4939
rect 20610 4871 20676 4905
rect 20610 4837 20626 4871
rect 20660 4837 20676 4871
rect 20610 4803 20676 4837
rect 20610 4769 20626 4803
rect 20660 4769 20676 4803
rect 20610 4735 20676 4769
rect 20610 4701 20626 4735
rect 20660 4701 20676 4735
rect 20610 4667 20676 4701
rect 20610 4633 20626 4667
rect 20660 4633 20676 4667
rect 20610 4599 20676 4633
rect 20610 4565 20626 4599
rect 20660 4565 20676 4599
rect 20610 4531 20676 4565
rect 20610 4497 20626 4531
rect 20660 4497 20676 4531
rect 20610 4463 20676 4497
rect 20610 4429 20626 4463
rect 20660 4429 20676 4463
rect 20610 4395 20676 4429
rect 20610 4361 20626 4395
rect 20660 4361 20676 4395
rect 20610 4327 20676 4361
rect 20610 4293 20626 4327
rect 20660 4293 20676 4327
rect 20610 4259 20676 4293
rect 20610 4225 20626 4259
rect 20660 4225 20676 4259
rect 20610 4191 20676 4225
rect 20610 4157 20626 4191
rect 20660 4157 20676 4191
rect 20610 4116 20676 4157
rect 20706 5075 20772 5116
rect 20706 5041 20722 5075
rect 20756 5041 20772 5075
rect 20706 5007 20772 5041
rect 20706 4973 20722 5007
rect 20756 4973 20772 5007
rect 20706 4939 20772 4973
rect 20706 4905 20722 4939
rect 20756 4905 20772 4939
rect 20706 4871 20772 4905
rect 20706 4837 20722 4871
rect 20756 4837 20772 4871
rect 20706 4803 20772 4837
rect 20706 4769 20722 4803
rect 20756 4769 20772 4803
rect 20706 4735 20772 4769
rect 20706 4701 20722 4735
rect 20756 4701 20772 4735
rect 20706 4667 20772 4701
rect 20706 4633 20722 4667
rect 20756 4633 20772 4667
rect 20706 4599 20772 4633
rect 20706 4565 20722 4599
rect 20756 4565 20772 4599
rect 20706 4531 20772 4565
rect 20706 4497 20722 4531
rect 20756 4497 20772 4531
rect 20706 4463 20772 4497
rect 20706 4429 20722 4463
rect 20756 4429 20772 4463
rect 20706 4395 20772 4429
rect 20706 4361 20722 4395
rect 20756 4361 20772 4395
rect 20706 4327 20772 4361
rect 20706 4293 20722 4327
rect 20756 4293 20772 4327
rect 20706 4259 20772 4293
rect 20706 4225 20722 4259
rect 20756 4225 20772 4259
rect 20706 4191 20772 4225
rect 20706 4157 20722 4191
rect 20756 4157 20772 4191
rect 20706 4116 20772 4157
rect 20802 5075 20868 5116
rect 20802 5041 20818 5075
rect 20852 5041 20868 5075
rect 20802 5007 20868 5041
rect 20802 4973 20818 5007
rect 20852 4973 20868 5007
rect 20802 4939 20868 4973
rect 20802 4905 20818 4939
rect 20852 4905 20868 4939
rect 20802 4871 20868 4905
rect 20802 4837 20818 4871
rect 20852 4837 20868 4871
rect 20802 4803 20868 4837
rect 20802 4769 20818 4803
rect 20852 4769 20868 4803
rect 20802 4735 20868 4769
rect 20802 4701 20818 4735
rect 20852 4701 20868 4735
rect 20802 4667 20868 4701
rect 20802 4633 20818 4667
rect 20852 4633 20868 4667
rect 20802 4599 20868 4633
rect 20802 4565 20818 4599
rect 20852 4565 20868 4599
rect 20802 4531 20868 4565
rect 20802 4497 20818 4531
rect 20852 4497 20868 4531
rect 20802 4463 20868 4497
rect 20802 4429 20818 4463
rect 20852 4429 20868 4463
rect 20802 4395 20868 4429
rect 20802 4361 20818 4395
rect 20852 4361 20868 4395
rect 20802 4327 20868 4361
rect 20802 4293 20818 4327
rect 20852 4293 20868 4327
rect 20802 4259 20868 4293
rect 20802 4225 20818 4259
rect 20852 4225 20868 4259
rect 20802 4191 20868 4225
rect 20802 4157 20818 4191
rect 20852 4157 20868 4191
rect 20802 4116 20868 4157
rect 20898 5075 20964 5116
rect 20898 5041 20914 5075
rect 20948 5041 20964 5075
rect 20898 5007 20964 5041
rect 20898 4973 20914 5007
rect 20948 4973 20964 5007
rect 20898 4939 20964 4973
rect 20898 4905 20914 4939
rect 20948 4905 20964 4939
rect 20898 4871 20964 4905
rect 20898 4837 20914 4871
rect 20948 4837 20964 4871
rect 20898 4803 20964 4837
rect 20898 4769 20914 4803
rect 20948 4769 20964 4803
rect 20898 4735 20964 4769
rect 20898 4701 20914 4735
rect 20948 4701 20964 4735
rect 20898 4667 20964 4701
rect 20898 4633 20914 4667
rect 20948 4633 20964 4667
rect 20898 4599 20964 4633
rect 20898 4565 20914 4599
rect 20948 4565 20964 4599
rect 20898 4531 20964 4565
rect 20898 4497 20914 4531
rect 20948 4497 20964 4531
rect 20898 4463 20964 4497
rect 20898 4429 20914 4463
rect 20948 4429 20964 4463
rect 20898 4395 20964 4429
rect 20898 4361 20914 4395
rect 20948 4361 20964 4395
rect 20898 4327 20964 4361
rect 20898 4293 20914 4327
rect 20948 4293 20964 4327
rect 20898 4259 20964 4293
rect 20898 4225 20914 4259
rect 20948 4225 20964 4259
rect 20898 4191 20964 4225
rect 20898 4157 20914 4191
rect 20948 4157 20964 4191
rect 20898 4116 20964 4157
rect 20994 5075 21060 5116
rect 20994 5041 21010 5075
rect 21044 5041 21060 5075
rect 20994 5007 21060 5041
rect 20994 4973 21010 5007
rect 21044 4973 21060 5007
rect 20994 4939 21060 4973
rect 20994 4905 21010 4939
rect 21044 4905 21060 4939
rect 20994 4871 21060 4905
rect 20994 4837 21010 4871
rect 21044 4837 21060 4871
rect 20994 4803 21060 4837
rect 20994 4769 21010 4803
rect 21044 4769 21060 4803
rect 20994 4735 21060 4769
rect 20994 4701 21010 4735
rect 21044 4701 21060 4735
rect 20994 4667 21060 4701
rect 20994 4633 21010 4667
rect 21044 4633 21060 4667
rect 20994 4599 21060 4633
rect 20994 4565 21010 4599
rect 21044 4565 21060 4599
rect 20994 4531 21060 4565
rect 20994 4497 21010 4531
rect 21044 4497 21060 4531
rect 20994 4463 21060 4497
rect 20994 4429 21010 4463
rect 21044 4429 21060 4463
rect 20994 4395 21060 4429
rect 20994 4361 21010 4395
rect 21044 4361 21060 4395
rect 20994 4327 21060 4361
rect 20994 4293 21010 4327
rect 21044 4293 21060 4327
rect 20994 4259 21060 4293
rect 20994 4225 21010 4259
rect 21044 4225 21060 4259
rect 20994 4191 21060 4225
rect 20994 4157 21010 4191
rect 21044 4157 21060 4191
rect 20994 4116 21060 4157
rect 21090 5075 21156 5116
rect 21090 5041 21106 5075
rect 21140 5041 21156 5075
rect 21090 5007 21156 5041
rect 21090 4973 21106 5007
rect 21140 4973 21156 5007
rect 21090 4939 21156 4973
rect 21090 4905 21106 4939
rect 21140 4905 21156 4939
rect 21090 4871 21156 4905
rect 21090 4837 21106 4871
rect 21140 4837 21156 4871
rect 21090 4803 21156 4837
rect 21090 4769 21106 4803
rect 21140 4769 21156 4803
rect 21090 4735 21156 4769
rect 21090 4701 21106 4735
rect 21140 4701 21156 4735
rect 21090 4667 21156 4701
rect 21090 4633 21106 4667
rect 21140 4633 21156 4667
rect 21090 4599 21156 4633
rect 21090 4565 21106 4599
rect 21140 4565 21156 4599
rect 21090 4531 21156 4565
rect 21090 4497 21106 4531
rect 21140 4497 21156 4531
rect 21090 4463 21156 4497
rect 21090 4429 21106 4463
rect 21140 4429 21156 4463
rect 21090 4395 21156 4429
rect 21090 4361 21106 4395
rect 21140 4361 21156 4395
rect 21090 4327 21156 4361
rect 21090 4293 21106 4327
rect 21140 4293 21156 4327
rect 21090 4259 21156 4293
rect 21090 4225 21106 4259
rect 21140 4225 21156 4259
rect 21090 4191 21156 4225
rect 21090 4157 21106 4191
rect 21140 4157 21156 4191
rect 21090 4116 21156 4157
rect 21186 5075 21252 5116
rect 21186 5041 21202 5075
rect 21236 5041 21252 5075
rect 21186 5007 21252 5041
rect 21186 4973 21202 5007
rect 21236 4973 21252 5007
rect 21186 4939 21252 4973
rect 21186 4905 21202 4939
rect 21236 4905 21252 4939
rect 21186 4871 21252 4905
rect 21186 4837 21202 4871
rect 21236 4837 21252 4871
rect 21186 4803 21252 4837
rect 21186 4769 21202 4803
rect 21236 4769 21252 4803
rect 21186 4735 21252 4769
rect 21186 4701 21202 4735
rect 21236 4701 21252 4735
rect 21186 4667 21252 4701
rect 21186 4633 21202 4667
rect 21236 4633 21252 4667
rect 21186 4599 21252 4633
rect 21186 4565 21202 4599
rect 21236 4565 21252 4599
rect 21186 4531 21252 4565
rect 21186 4497 21202 4531
rect 21236 4497 21252 4531
rect 21186 4463 21252 4497
rect 21186 4429 21202 4463
rect 21236 4429 21252 4463
rect 21186 4395 21252 4429
rect 21186 4361 21202 4395
rect 21236 4361 21252 4395
rect 21186 4327 21252 4361
rect 21186 4293 21202 4327
rect 21236 4293 21252 4327
rect 21186 4259 21252 4293
rect 21186 4225 21202 4259
rect 21236 4225 21252 4259
rect 21186 4191 21252 4225
rect 21186 4157 21202 4191
rect 21236 4157 21252 4191
rect 21186 4116 21252 4157
rect 21282 5075 21348 5116
rect 21282 5041 21298 5075
rect 21332 5041 21348 5075
rect 21282 5007 21348 5041
rect 21282 4973 21298 5007
rect 21332 4973 21348 5007
rect 21282 4939 21348 4973
rect 21282 4905 21298 4939
rect 21332 4905 21348 4939
rect 21282 4871 21348 4905
rect 21282 4837 21298 4871
rect 21332 4837 21348 4871
rect 21282 4803 21348 4837
rect 21282 4769 21298 4803
rect 21332 4769 21348 4803
rect 21282 4735 21348 4769
rect 21282 4701 21298 4735
rect 21332 4701 21348 4735
rect 21282 4667 21348 4701
rect 21282 4633 21298 4667
rect 21332 4633 21348 4667
rect 21282 4599 21348 4633
rect 21282 4565 21298 4599
rect 21332 4565 21348 4599
rect 21282 4531 21348 4565
rect 21282 4497 21298 4531
rect 21332 4497 21348 4531
rect 21282 4463 21348 4497
rect 21282 4429 21298 4463
rect 21332 4429 21348 4463
rect 21282 4395 21348 4429
rect 21282 4361 21298 4395
rect 21332 4361 21348 4395
rect 21282 4327 21348 4361
rect 21282 4293 21298 4327
rect 21332 4293 21348 4327
rect 21282 4259 21348 4293
rect 21282 4225 21298 4259
rect 21332 4225 21348 4259
rect 21282 4191 21348 4225
rect 21282 4157 21298 4191
rect 21332 4157 21348 4191
rect 21282 4116 21348 4157
rect 21378 5075 21444 5116
rect 21378 5041 21394 5075
rect 21428 5041 21444 5075
rect 21378 5007 21444 5041
rect 21378 4973 21394 5007
rect 21428 4973 21444 5007
rect 21378 4939 21444 4973
rect 21378 4905 21394 4939
rect 21428 4905 21444 4939
rect 21378 4871 21444 4905
rect 21378 4837 21394 4871
rect 21428 4837 21444 4871
rect 21378 4803 21444 4837
rect 21378 4769 21394 4803
rect 21428 4769 21444 4803
rect 21378 4735 21444 4769
rect 21378 4701 21394 4735
rect 21428 4701 21444 4735
rect 21378 4667 21444 4701
rect 21378 4633 21394 4667
rect 21428 4633 21444 4667
rect 21378 4599 21444 4633
rect 21378 4565 21394 4599
rect 21428 4565 21444 4599
rect 21378 4531 21444 4565
rect 21378 4497 21394 4531
rect 21428 4497 21444 4531
rect 21378 4463 21444 4497
rect 21378 4429 21394 4463
rect 21428 4429 21444 4463
rect 21378 4395 21444 4429
rect 21378 4361 21394 4395
rect 21428 4361 21444 4395
rect 21378 4327 21444 4361
rect 21378 4293 21394 4327
rect 21428 4293 21444 4327
rect 21378 4259 21444 4293
rect 21378 4225 21394 4259
rect 21428 4225 21444 4259
rect 21378 4191 21444 4225
rect 21378 4157 21394 4191
rect 21428 4157 21444 4191
rect 21378 4116 21444 4157
rect 21474 5075 21540 5116
rect 21474 5041 21490 5075
rect 21524 5041 21540 5075
rect 21474 5007 21540 5041
rect 21474 4973 21490 5007
rect 21524 4973 21540 5007
rect 21474 4939 21540 4973
rect 21474 4905 21490 4939
rect 21524 4905 21540 4939
rect 21474 4871 21540 4905
rect 21474 4837 21490 4871
rect 21524 4837 21540 4871
rect 21474 4803 21540 4837
rect 21474 4769 21490 4803
rect 21524 4769 21540 4803
rect 21474 4735 21540 4769
rect 21474 4701 21490 4735
rect 21524 4701 21540 4735
rect 21474 4667 21540 4701
rect 21474 4633 21490 4667
rect 21524 4633 21540 4667
rect 21474 4599 21540 4633
rect 21474 4565 21490 4599
rect 21524 4565 21540 4599
rect 21474 4531 21540 4565
rect 21474 4497 21490 4531
rect 21524 4497 21540 4531
rect 21474 4463 21540 4497
rect 21474 4429 21490 4463
rect 21524 4429 21540 4463
rect 21474 4395 21540 4429
rect 21474 4361 21490 4395
rect 21524 4361 21540 4395
rect 21474 4327 21540 4361
rect 21474 4293 21490 4327
rect 21524 4293 21540 4327
rect 21474 4259 21540 4293
rect 21474 4225 21490 4259
rect 21524 4225 21540 4259
rect 21474 4191 21540 4225
rect 21474 4157 21490 4191
rect 21524 4157 21540 4191
rect 21474 4116 21540 4157
rect 21570 5075 21636 5116
rect 21570 5041 21586 5075
rect 21620 5041 21636 5075
rect 21570 5007 21636 5041
rect 21570 4973 21586 5007
rect 21620 4973 21636 5007
rect 21570 4939 21636 4973
rect 21570 4905 21586 4939
rect 21620 4905 21636 4939
rect 21570 4871 21636 4905
rect 21570 4837 21586 4871
rect 21620 4837 21636 4871
rect 21570 4803 21636 4837
rect 21570 4769 21586 4803
rect 21620 4769 21636 4803
rect 21570 4735 21636 4769
rect 21570 4701 21586 4735
rect 21620 4701 21636 4735
rect 21570 4667 21636 4701
rect 21570 4633 21586 4667
rect 21620 4633 21636 4667
rect 21570 4599 21636 4633
rect 21570 4565 21586 4599
rect 21620 4565 21636 4599
rect 21570 4531 21636 4565
rect 21570 4497 21586 4531
rect 21620 4497 21636 4531
rect 21570 4463 21636 4497
rect 21570 4429 21586 4463
rect 21620 4429 21636 4463
rect 21570 4395 21636 4429
rect 21570 4361 21586 4395
rect 21620 4361 21636 4395
rect 21570 4327 21636 4361
rect 21570 4293 21586 4327
rect 21620 4293 21636 4327
rect 21570 4259 21636 4293
rect 21570 4225 21586 4259
rect 21620 4225 21636 4259
rect 21570 4191 21636 4225
rect 21570 4157 21586 4191
rect 21620 4157 21636 4191
rect 21570 4116 21636 4157
rect 21666 5075 21732 5116
rect 21666 5041 21682 5075
rect 21716 5041 21732 5075
rect 21666 5007 21732 5041
rect 21666 4973 21682 5007
rect 21716 4973 21732 5007
rect 21666 4939 21732 4973
rect 21666 4905 21682 4939
rect 21716 4905 21732 4939
rect 21666 4871 21732 4905
rect 21666 4837 21682 4871
rect 21716 4837 21732 4871
rect 21666 4803 21732 4837
rect 21666 4769 21682 4803
rect 21716 4769 21732 4803
rect 21666 4735 21732 4769
rect 21666 4701 21682 4735
rect 21716 4701 21732 4735
rect 21666 4667 21732 4701
rect 21666 4633 21682 4667
rect 21716 4633 21732 4667
rect 21666 4599 21732 4633
rect 21666 4565 21682 4599
rect 21716 4565 21732 4599
rect 21666 4531 21732 4565
rect 21666 4497 21682 4531
rect 21716 4497 21732 4531
rect 21666 4463 21732 4497
rect 21666 4429 21682 4463
rect 21716 4429 21732 4463
rect 21666 4395 21732 4429
rect 21666 4361 21682 4395
rect 21716 4361 21732 4395
rect 21666 4327 21732 4361
rect 21666 4293 21682 4327
rect 21716 4293 21732 4327
rect 21666 4259 21732 4293
rect 21666 4225 21682 4259
rect 21716 4225 21732 4259
rect 21666 4191 21732 4225
rect 21666 4157 21682 4191
rect 21716 4157 21732 4191
rect 21666 4116 21732 4157
rect 21762 5075 21828 5116
rect 21762 5041 21778 5075
rect 21812 5041 21828 5075
rect 21762 5007 21828 5041
rect 21762 4973 21778 5007
rect 21812 4973 21828 5007
rect 21762 4939 21828 4973
rect 21762 4905 21778 4939
rect 21812 4905 21828 4939
rect 21762 4871 21828 4905
rect 21762 4837 21778 4871
rect 21812 4837 21828 4871
rect 21762 4803 21828 4837
rect 21762 4769 21778 4803
rect 21812 4769 21828 4803
rect 21762 4735 21828 4769
rect 21762 4701 21778 4735
rect 21812 4701 21828 4735
rect 21762 4667 21828 4701
rect 21762 4633 21778 4667
rect 21812 4633 21828 4667
rect 21762 4599 21828 4633
rect 21762 4565 21778 4599
rect 21812 4565 21828 4599
rect 21762 4531 21828 4565
rect 21762 4497 21778 4531
rect 21812 4497 21828 4531
rect 21762 4463 21828 4497
rect 21762 4429 21778 4463
rect 21812 4429 21828 4463
rect 21762 4395 21828 4429
rect 21762 4361 21778 4395
rect 21812 4361 21828 4395
rect 21762 4327 21828 4361
rect 21762 4293 21778 4327
rect 21812 4293 21828 4327
rect 21762 4259 21828 4293
rect 21762 4225 21778 4259
rect 21812 4225 21828 4259
rect 21762 4191 21828 4225
rect 21762 4157 21778 4191
rect 21812 4157 21828 4191
rect 21762 4116 21828 4157
rect 21858 5075 21924 5116
rect 21858 5041 21874 5075
rect 21908 5041 21924 5075
rect 21858 5007 21924 5041
rect 21858 4973 21874 5007
rect 21908 4973 21924 5007
rect 21858 4939 21924 4973
rect 21858 4905 21874 4939
rect 21908 4905 21924 4939
rect 21858 4871 21924 4905
rect 21858 4837 21874 4871
rect 21908 4837 21924 4871
rect 21858 4803 21924 4837
rect 21858 4769 21874 4803
rect 21908 4769 21924 4803
rect 21858 4735 21924 4769
rect 21858 4701 21874 4735
rect 21908 4701 21924 4735
rect 21858 4667 21924 4701
rect 21858 4633 21874 4667
rect 21908 4633 21924 4667
rect 21858 4599 21924 4633
rect 21858 4565 21874 4599
rect 21908 4565 21924 4599
rect 21858 4531 21924 4565
rect 21858 4497 21874 4531
rect 21908 4497 21924 4531
rect 21858 4463 21924 4497
rect 21858 4429 21874 4463
rect 21908 4429 21924 4463
rect 21858 4395 21924 4429
rect 21858 4361 21874 4395
rect 21908 4361 21924 4395
rect 21858 4327 21924 4361
rect 21858 4293 21874 4327
rect 21908 4293 21924 4327
rect 21858 4259 21924 4293
rect 21858 4225 21874 4259
rect 21908 4225 21924 4259
rect 21858 4191 21924 4225
rect 21858 4157 21874 4191
rect 21908 4157 21924 4191
rect 21858 4116 21924 4157
rect 21954 5075 22020 5116
rect 21954 5041 21970 5075
rect 22004 5041 22020 5075
rect 21954 5007 22020 5041
rect 21954 4973 21970 5007
rect 22004 4973 22020 5007
rect 21954 4939 22020 4973
rect 21954 4905 21970 4939
rect 22004 4905 22020 4939
rect 21954 4871 22020 4905
rect 21954 4837 21970 4871
rect 22004 4837 22020 4871
rect 21954 4803 22020 4837
rect 21954 4769 21970 4803
rect 22004 4769 22020 4803
rect 21954 4735 22020 4769
rect 21954 4701 21970 4735
rect 22004 4701 22020 4735
rect 21954 4667 22020 4701
rect 21954 4633 21970 4667
rect 22004 4633 22020 4667
rect 21954 4599 22020 4633
rect 21954 4565 21970 4599
rect 22004 4565 22020 4599
rect 21954 4531 22020 4565
rect 21954 4497 21970 4531
rect 22004 4497 22020 4531
rect 21954 4463 22020 4497
rect 21954 4429 21970 4463
rect 22004 4429 22020 4463
rect 21954 4395 22020 4429
rect 21954 4361 21970 4395
rect 22004 4361 22020 4395
rect 21954 4327 22020 4361
rect 21954 4293 21970 4327
rect 22004 4293 22020 4327
rect 21954 4259 22020 4293
rect 21954 4225 21970 4259
rect 22004 4225 22020 4259
rect 21954 4191 22020 4225
rect 21954 4157 21970 4191
rect 22004 4157 22020 4191
rect 21954 4116 22020 4157
rect 22050 5075 22116 5116
rect 22050 5041 22066 5075
rect 22100 5041 22116 5075
rect 22050 5007 22116 5041
rect 22050 4973 22066 5007
rect 22100 4973 22116 5007
rect 22050 4939 22116 4973
rect 22050 4905 22066 4939
rect 22100 4905 22116 4939
rect 22050 4871 22116 4905
rect 22050 4837 22066 4871
rect 22100 4837 22116 4871
rect 22050 4803 22116 4837
rect 22050 4769 22066 4803
rect 22100 4769 22116 4803
rect 22050 4735 22116 4769
rect 22050 4701 22066 4735
rect 22100 4701 22116 4735
rect 22050 4667 22116 4701
rect 22050 4633 22066 4667
rect 22100 4633 22116 4667
rect 22050 4599 22116 4633
rect 22050 4565 22066 4599
rect 22100 4565 22116 4599
rect 22050 4531 22116 4565
rect 22050 4497 22066 4531
rect 22100 4497 22116 4531
rect 22050 4463 22116 4497
rect 22050 4429 22066 4463
rect 22100 4429 22116 4463
rect 22050 4395 22116 4429
rect 22050 4361 22066 4395
rect 22100 4361 22116 4395
rect 22050 4327 22116 4361
rect 22050 4293 22066 4327
rect 22100 4293 22116 4327
rect 22050 4259 22116 4293
rect 22050 4225 22066 4259
rect 22100 4225 22116 4259
rect 22050 4191 22116 4225
rect 22050 4157 22066 4191
rect 22100 4157 22116 4191
rect 22050 4116 22116 4157
rect 22146 5075 22212 5116
rect 22146 5041 22162 5075
rect 22196 5041 22212 5075
rect 22146 5007 22212 5041
rect 22146 4973 22162 5007
rect 22196 4973 22212 5007
rect 22146 4939 22212 4973
rect 22146 4905 22162 4939
rect 22196 4905 22212 4939
rect 22146 4871 22212 4905
rect 22146 4837 22162 4871
rect 22196 4837 22212 4871
rect 22146 4803 22212 4837
rect 22146 4769 22162 4803
rect 22196 4769 22212 4803
rect 22146 4735 22212 4769
rect 22146 4701 22162 4735
rect 22196 4701 22212 4735
rect 22146 4667 22212 4701
rect 22146 4633 22162 4667
rect 22196 4633 22212 4667
rect 22146 4599 22212 4633
rect 22146 4565 22162 4599
rect 22196 4565 22212 4599
rect 22146 4531 22212 4565
rect 22146 4497 22162 4531
rect 22196 4497 22212 4531
rect 22146 4463 22212 4497
rect 22146 4429 22162 4463
rect 22196 4429 22212 4463
rect 22146 4395 22212 4429
rect 22146 4361 22162 4395
rect 22196 4361 22212 4395
rect 22146 4327 22212 4361
rect 22146 4293 22162 4327
rect 22196 4293 22212 4327
rect 22146 4259 22212 4293
rect 22146 4225 22162 4259
rect 22196 4225 22212 4259
rect 22146 4191 22212 4225
rect 22146 4157 22162 4191
rect 22196 4157 22212 4191
rect 22146 4116 22212 4157
rect 22242 5075 22304 5116
rect 22242 5041 22258 5075
rect 22292 5041 22304 5075
rect 22242 5007 22304 5041
rect 22242 4973 22258 5007
rect 22292 4973 22304 5007
rect 22242 4939 22304 4973
rect 22242 4905 22258 4939
rect 22292 4905 22304 4939
rect 22242 4871 22304 4905
rect 22242 4837 22258 4871
rect 22292 4837 22304 4871
rect 22242 4803 22304 4837
rect 22242 4769 22258 4803
rect 22292 4769 22304 4803
rect 22242 4735 22304 4769
rect 22242 4701 22258 4735
rect 22292 4701 22304 4735
rect 22242 4667 22304 4701
rect 22242 4633 22258 4667
rect 22292 4633 22304 4667
rect 22242 4599 22304 4633
rect 22242 4565 22258 4599
rect 22292 4565 22304 4599
rect 22242 4531 22304 4565
rect 22242 4497 22258 4531
rect 22292 4497 22304 4531
rect 22242 4463 22304 4497
rect 22242 4429 22258 4463
rect 22292 4429 22304 4463
rect 22242 4395 22304 4429
rect 22242 4361 22258 4395
rect 22292 4361 22304 4395
rect 22242 4327 22304 4361
rect 22242 4293 22258 4327
rect 22292 4293 22304 4327
rect 22242 4259 22304 4293
rect 22242 4225 22258 4259
rect 22292 4225 22304 4259
rect 22242 4191 22304 4225
rect 22242 4157 22258 4191
rect 22292 4157 22304 4191
rect 22242 4116 22304 4157
rect 23258 5087 23320 5128
rect 23258 5053 23270 5087
rect 23304 5053 23320 5087
rect 23258 5019 23320 5053
rect 23258 4985 23270 5019
rect 23304 4985 23320 5019
rect 23258 4951 23320 4985
rect 23258 4917 23270 4951
rect 23304 4917 23320 4951
rect 23258 4883 23320 4917
rect 23258 4849 23270 4883
rect 23304 4849 23320 4883
rect 23258 4815 23320 4849
rect 23258 4781 23270 4815
rect 23304 4781 23320 4815
rect 23258 4747 23320 4781
rect 23258 4713 23270 4747
rect 23304 4713 23320 4747
rect 23258 4679 23320 4713
rect 23258 4645 23270 4679
rect 23304 4645 23320 4679
rect 23258 4611 23320 4645
rect 23258 4577 23270 4611
rect 23304 4577 23320 4611
rect 23258 4543 23320 4577
rect 23258 4509 23270 4543
rect 23304 4509 23320 4543
rect 23258 4475 23320 4509
rect 23258 4441 23270 4475
rect 23304 4441 23320 4475
rect 23258 4407 23320 4441
rect 23258 4373 23270 4407
rect 23304 4373 23320 4407
rect 23258 4339 23320 4373
rect 23258 4305 23270 4339
rect 23304 4305 23320 4339
rect 23258 4271 23320 4305
rect 23258 4237 23270 4271
rect 23304 4237 23320 4271
rect 23258 4203 23320 4237
rect 23258 4169 23270 4203
rect 23304 4169 23320 4203
rect 23258 4128 23320 4169
rect 23350 5087 23416 5128
rect 23350 5053 23366 5087
rect 23400 5053 23416 5087
rect 23350 5019 23416 5053
rect 23350 4985 23366 5019
rect 23400 4985 23416 5019
rect 23350 4951 23416 4985
rect 23350 4917 23366 4951
rect 23400 4917 23416 4951
rect 23350 4883 23416 4917
rect 23350 4849 23366 4883
rect 23400 4849 23416 4883
rect 23350 4815 23416 4849
rect 23350 4781 23366 4815
rect 23400 4781 23416 4815
rect 23350 4747 23416 4781
rect 23350 4713 23366 4747
rect 23400 4713 23416 4747
rect 23350 4679 23416 4713
rect 23350 4645 23366 4679
rect 23400 4645 23416 4679
rect 23350 4611 23416 4645
rect 23350 4577 23366 4611
rect 23400 4577 23416 4611
rect 23350 4543 23416 4577
rect 23350 4509 23366 4543
rect 23400 4509 23416 4543
rect 23350 4475 23416 4509
rect 23350 4441 23366 4475
rect 23400 4441 23416 4475
rect 23350 4407 23416 4441
rect 23350 4373 23366 4407
rect 23400 4373 23416 4407
rect 23350 4339 23416 4373
rect 23350 4305 23366 4339
rect 23400 4305 23416 4339
rect 23350 4271 23416 4305
rect 23350 4237 23366 4271
rect 23400 4237 23416 4271
rect 23350 4203 23416 4237
rect 23350 4169 23366 4203
rect 23400 4169 23416 4203
rect 23350 4128 23416 4169
rect 23446 5087 23512 5128
rect 23446 5053 23462 5087
rect 23496 5053 23512 5087
rect 23446 5019 23512 5053
rect 23446 4985 23462 5019
rect 23496 4985 23512 5019
rect 23446 4951 23512 4985
rect 23446 4917 23462 4951
rect 23496 4917 23512 4951
rect 23446 4883 23512 4917
rect 23446 4849 23462 4883
rect 23496 4849 23512 4883
rect 23446 4815 23512 4849
rect 23446 4781 23462 4815
rect 23496 4781 23512 4815
rect 23446 4747 23512 4781
rect 23446 4713 23462 4747
rect 23496 4713 23512 4747
rect 23446 4679 23512 4713
rect 23446 4645 23462 4679
rect 23496 4645 23512 4679
rect 23446 4611 23512 4645
rect 23446 4577 23462 4611
rect 23496 4577 23512 4611
rect 23446 4543 23512 4577
rect 23446 4509 23462 4543
rect 23496 4509 23512 4543
rect 23446 4475 23512 4509
rect 23446 4441 23462 4475
rect 23496 4441 23512 4475
rect 23446 4407 23512 4441
rect 23446 4373 23462 4407
rect 23496 4373 23512 4407
rect 23446 4339 23512 4373
rect 23446 4305 23462 4339
rect 23496 4305 23512 4339
rect 23446 4271 23512 4305
rect 23446 4237 23462 4271
rect 23496 4237 23512 4271
rect 23446 4203 23512 4237
rect 23446 4169 23462 4203
rect 23496 4169 23512 4203
rect 23446 4128 23512 4169
rect 23542 5087 23608 5128
rect 23542 5053 23558 5087
rect 23592 5053 23608 5087
rect 23542 5019 23608 5053
rect 23542 4985 23558 5019
rect 23592 4985 23608 5019
rect 23542 4951 23608 4985
rect 23542 4917 23558 4951
rect 23592 4917 23608 4951
rect 23542 4883 23608 4917
rect 23542 4849 23558 4883
rect 23592 4849 23608 4883
rect 23542 4815 23608 4849
rect 23542 4781 23558 4815
rect 23592 4781 23608 4815
rect 23542 4747 23608 4781
rect 23542 4713 23558 4747
rect 23592 4713 23608 4747
rect 23542 4679 23608 4713
rect 23542 4645 23558 4679
rect 23592 4645 23608 4679
rect 23542 4611 23608 4645
rect 23542 4577 23558 4611
rect 23592 4577 23608 4611
rect 23542 4543 23608 4577
rect 23542 4509 23558 4543
rect 23592 4509 23608 4543
rect 23542 4475 23608 4509
rect 23542 4441 23558 4475
rect 23592 4441 23608 4475
rect 23542 4407 23608 4441
rect 23542 4373 23558 4407
rect 23592 4373 23608 4407
rect 23542 4339 23608 4373
rect 23542 4305 23558 4339
rect 23592 4305 23608 4339
rect 23542 4271 23608 4305
rect 23542 4237 23558 4271
rect 23592 4237 23608 4271
rect 23542 4203 23608 4237
rect 23542 4169 23558 4203
rect 23592 4169 23608 4203
rect 23542 4128 23608 4169
rect 23638 5087 23704 5128
rect 23638 5053 23654 5087
rect 23688 5053 23704 5087
rect 23638 5019 23704 5053
rect 23638 4985 23654 5019
rect 23688 4985 23704 5019
rect 23638 4951 23704 4985
rect 23638 4917 23654 4951
rect 23688 4917 23704 4951
rect 23638 4883 23704 4917
rect 23638 4849 23654 4883
rect 23688 4849 23704 4883
rect 23638 4815 23704 4849
rect 23638 4781 23654 4815
rect 23688 4781 23704 4815
rect 23638 4747 23704 4781
rect 23638 4713 23654 4747
rect 23688 4713 23704 4747
rect 23638 4679 23704 4713
rect 23638 4645 23654 4679
rect 23688 4645 23704 4679
rect 23638 4611 23704 4645
rect 23638 4577 23654 4611
rect 23688 4577 23704 4611
rect 23638 4543 23704 4577
rect 23638 4509 23654 4543
rect 23688 4509 23704 4543
rect 23638 4475 23704 4509
rect 23638 4441 23654 4475
rect 23688 4441 23704 4475
rect 23638 4407 23704 4441
rect 23638 4373 23654 4407
rect 23688 4373 23704 4407
rect 23638 4339 23704 4373
rect 23638 4305 23654 4339
rect 23688 4305 23704 4339
rect 23638 4271 23704 4305
rect 23638 4237 23654 4271
rect 23688 4237 23704 4271
rect 23638 4203 23704 4237
rect 23638 4169 23654 4203
rect 23688 4169 23704 4203
rect 23638 4128 23704 4169
rect 23734 5087 23796 5128
rect 23734 5053 23750 5087
rect 23784 5053 23796 5087
rect 23734 5019 23796 5053
rect 23734 4985 23750 5019
rect 23784 4985 23796 5019
rect 23734 4951 23796 4985
rect 23734 4917 23750 4951
rect 23784 4917 23796 4951
rect 23734 4883 23796 4917
rect 23734 4849 23750 4883
rect 23784 4849 23796 4883
rect 23734 4815 23796 4849
rect 23734 4781 23750 4815
rect 23784 4781 23796 4815
rect 23734 4747 23796 4781
rect 23734 4713 23750 4747
rect 23784 4713 23796 4747
rect 23734 4679 23796 4713
rect 23734 4645 23750 4679
rect 23784 4645 23796 4679
rect 23734 4611 23796 4645
rect 23734 4577 23750 4611
rect 23784 4577 23796 4611
rect 23734 4543 23796 4577
rect 23734 4509 23750 4543
rect 23784 4509 23796 4543
rect 23734 4475 23796 4509
rect 23734 4441 23750 4475
rect 23784 4441 23796 4475
rect 23734 4407 23796 4441
rect 23734 4373 23750 4407
rect 23784 4373 23796 4407
rect 23734 4339 23796 4373
rect 23734 4305 23750 4339
rect 23784 4305 23796 4339
rect 23734 4271 23796 4305
rect 23734 4237 23750 4271
rect 23784 4237 23796 4271
rect 23734 4203 23796 4237
rect 23734 4169 23750 4203
rect 23784 4169 23796 4203
rect 23734 4128 23796 4169
rect 23946 5085 24008 5126
rect 23946 5051 23958 5085
rect 23992 5051 24008 5085
rect 23946 5017 24008 5051
rect 23946 4983 23958 5017
rect 23992 4983 24008 5017
rect 23946 4949 24008 4983
rect 23946 4915 23958 4949
rect 23992 4915 24008 4949
rect 23946 4881 24008 4915
rect 23946 4847 23958 4881
rect 23992 4847 24008 4881
rect 23946 4813 24008 4847
rect 23946 4779 23958 4813
rect 23992 4779 24008 4813
rect 23946 4745 24008 4779
rect 23946 4711 23958 4745
rect 23992 4711 24008 4745
rect 23946 4677 24008 4711
rect 23946 4643 23958 4677
rect 23992 4643 24008 4677
rect 23946 4609 24008 4643
rect 23946 4575 23958 4609
rect 23992 4575 24008 4609
rect 23946 4541 24008 4575
rect 23946 4507 23958 4541
rect 23992 4507 24008 4541
rect 23946 4473 24008 4507
rect 23946 4439 23958 4473
rect 23992 4439 24008 4473
rect 23946 4405 24008 4439
rect 23946 4371 23958 4405
rect 23992 4371 24008 4405
rect 23946 4337 24008 4371
rect 23946 4303 23958 4337
rect 23992 4303 24008 4337
rect 23946 4269 24008 4303
rect 23946 4235 23958 4269
rect 23992 4235 24008 4269
rect 23946 4201 24008 4235
rect 23946 4167 23958 4201
rect 23992 4167 24008 4201
rect 23946 4126 24008 4167
rect 24038 5085 24104 5126
rect 24038 5051 24054 5085
rect 24088 5051 24104 5085
rect 24038 5017 24104 5051
rect 24038 4983 24054 5017
rect 24088 4983 24104 5017
rect 24038 4949 24104 4983
rect 24038 4915 24054 4949
rect 24088 4915 24104 4949
rect 24038 4881 24104 4915
rect 24038 4847 24054 4881
rect 24088 4847 24104 4881
rect 24038 4813 24104 4847
rect 24038 4779 24054 4813
rect 24088 4779 24104 4813
rect 24038 4745 24104 4779
rect 24038 4711 24054 4745
rect 24088 4711 24104 4745
rect 24038 4677 24104 4711
rect 24038 4643 24054 4677
rect 24088 4643 24104 4677
rect 24038 4609 24104 4643
rect 24038 4575 24054 4609
rect 24088 4575 24104 4609
rect 24038 4541 24104 4575
rect 24038 4507 24054 4541
rect 24088 4507 24104 4541
rect 24038 4473 24104 4507
rect 24038 4439 24054 4473
rect 24088 4439 24104 4473
rect 24038 4405 24104 4439
rect 24038 4371 24054 4405
rect 24088 4371 24104 4405
rect 24038 4337 24104 4371
rect 24038 4303 24054 4337
rect 24088 4303 24104 4337
rect 24038 4269 24104 4303
rect 24038 4235 24054 4269
rect 24088 4235 24104 4269
rect 24038 4201 24104 4235
rect 24038 4167 24054 4201
rect 24088 4167 24104 4201
rect 24038 4126 24104 4167
rect 24134 5085 24200 5126
rect 24134 5051 24150 5085
rect 24184 5051 24200 5085
rect 24134 5017 24200 5051
rect 24134 4983 24150 5017
rect 24184 4983 24200 5017
rect 24134 4949 24200 4983
rect 24134 4915 24150 4949
rect 24184 4915 24200 4949
rect 24134 4881 24200 4915
rect 24134 4847 24150 4881
rect 24184 4847 24200 4881
rect 24134 4813 24200 4847
rect 24134 4779 24150 4813
rect 24184 4779 24200 4813
rect 24134 4745 24200 4779
rect 24134 4711 24150 4745
rect 24184 4711 24200 4745
rect 24134 4677 24200 4711
rect 24134 4643 24150 4677
rect 24184 4643 24200 4677
rect 24134 4609 24200 4643
rect 24134 4575 24150 4609
rect 24184 4575 24200 4609
rect 24134 4541 24200 4575
rect 24134 4507 24150 4541
rect 24184 4507 24200 4541
rect 24134 4473 24200 4507
rect 24134 4439 24150 4473
rect 24184 4439 24200 4473
rect 24134 4405 24200 4439
rect 24134 4371 24150 4405
rect 24184 4371 24200 4405
rect 24134 4337 24200 4371
rect 24134 4303 24150 4337
rect 24184 4303 24200 4337
rect 24134 4269 24200 4303
rect 24134 4235 24150 4269
rect 24184 4235 24200 4269
rect 24134 4201 24200 4235
rect 24134 4167 24150 4201
rect 24184 4167 24200 4201
rect 24134 4126 24200 4167
rect 24230 5085 24296 5126
rect 24230 5051 24246 5085
rect 24280 5051 24296 5085
rect 24230 5017 24296 5051
rect 24230 4983 24246 5017
rect 24280 4983 24296 5017
rect 24230 4949 24296 4983
rect 24230 4915 24246 4949
rect 24280 4915 24296 4949
rect 24230 4881 24296 4915
rect 24230 4847 24246 4881
rect 24280 4847 24296 4881
rect 24230 4813 24296 4847
rect 24230 4779 24246 4813
rect 24280 4779 24296 4813
rect 24230 4745 24296 4779
rect 24230 4711 24246 4745
rect 24280 4711 24296 4745
rect 24230 4677 24296 4711
rect 24230 4643 24246 4677
rect 24280 4643 24296 4677
rect 24230 4609 24296 4643
rect 24230 4575 24246 4609
rect 24280 4575 24296 4609
rect 24230 4541 24296 4575
rect 24230 4507 24246 4541
rect 24280 4507 24296 4541
rect 24230 4473 24296 4507
rect 24230 4439 24246 4473
rect 24280 4439 24296 4473
rect 24230 4405 24296 4439
rect 24230 4371 24246 4405
rect 24280 4371 24296 4405
rect 24230 4337 24296 4371
rect 24230 4303 24246 4337
rect 24280 4303 24296 4337
rect 24230 4269 24296 4303
rect 24230 4235 24246 4269
rect 24280 4235 24296 4269
rect 24230 4201 24296 4235
rect 24230 4167 24246 4201
rect 24280 4167 24296 4201
rect 24230 4126 24296 4167
rect 24326 5085 24392 5126
rect 24326 5051 24342 5085
rect 24376 5051 24392 5085
rect 24326 5017 24392 5051
rect 24326 4983 24342 5017
rect 24376 4983 24392 5017
rect 24326 4949 24392 4983
rect 24326 4915 24342 4949
rect 24376 4915 24392 4949
rect 24326 4881 24392 4915
rect 24326 4847 24342 4881
rect 24376 4847 24392 4881
rect 24326 4813 24392 4847
rect 24326 4779 24342 4813
rect 24376 4779 24392 4813
rect 24326 4745 24392 4779
rect 24326 4711 24342 4745
rect 24376 4711 24392 4745
rect 24326 4677 24392 4711
rect 24326 4643 24342 4677
rect 24376 4643 24392 4677
rect 24326 4609 24392 4643
rect 24326 4575 24342 4609
rect 24376 4575 24392 4609
rect 24326 4541 24392 4575
rect 24326 4507 24342 4541
rect 24376 4507 24392 4541
rect 24326 4473 24392 4507
rect 24326 4439 24342 4473
rect 24376 4439 24392 4473
rect 24326 4405 24392 4439
rect 24326 4371 24342 4405
rect 24376 4371 24392 4405
rect 24326 4337 24392 4371
rect 24326 4303 24342 4337
rect 24376 4303 24392 4337
rect 24326 4269 24392 4303
rect 24326 4235 24342 4269
rect 24376 4235 24392 4269
rect 24326 4201 24392 4235
rect 24326 4167 24342 4201
rect 24376 4167 24392 4201
rect 24326 4126 24392 4167
rect 24422 5085 24488 5126
rect 24422 5051 24438 5085
rect 24472 5051 24488 5085
rect 24422 5017 24488 5051
rect 24422 4983 24438 5017
rect 24472 4983 24488 5017
rect 24422 4949 24488 4983
rect 24422 4915 24438 4949
rect 24472 4915 24488 4949
rect 24422 4881 24488 4915
rect 24422 4847 24438 4881
rect 24472 4847 24488 4881
rect 24422 4813 24488 4847
rect 24422 4779 24438 4813
rect 24472 4779 24488 4813
rect 24422 4745 24488 4779
rect 24422 4711 24438 4745
rect 24472 4711 24488 4745
rect 24422 4677 24488 4711
rect 24422 4643 24438 4677
rect 24472 4643 24488 4677
rect 24422 4609 24488 4643
rect 24422 4575 24438 4609
rect 24472 4575 24488 4609
rect 24422 4541 24488 4575
rect 24422 4507 24438 4541
rect 24472 4507 24488 4541
rect 24422 4473 24488 4507
rect 24422 4439 24438 4473
rect 24472 4439 24488 4473
rect 24422 4405 24488 4439
rect 24422 4371 24438 4405
rect 24472 4371 24488 4405
rect 24422 4337 24488 4371
rect 24422 4303 24438 4337
rect 24472 4303 24488 4337
rect 24422 4269 24488 4303
rect 24422 4235 24438 4269
rect 24472 4235 24488 4269
rect 24422 4201 24488 4235
rect 24422 4167 24438 4201
rect 24472 4167 24488 4201
rect 24422 4126 24488 4167
rect 24518 5085 24584 5126
rect 24518 5051 24534 5085
rect 24568 5051 24584 5085
rect 24518 5017 24584 5051
rect 24518 4983 24534 5017
rect 24568 4983 24584 5017
rect 24518 4949 24584 4983
rect 24518 4915 24534 4949
rect 24568 4915 24584 4949
rect 24518 4881 24584 4915
rect 24518 4847 24534 4881
rect 24568 4847 24584 4881
rect 24518 4813 24584 4847
rect 24518 4779 24534 4813
rect 24568 4779 24584 4813
rect 24518 4745 24584 4779
rect 24518 4711 24534 4745
rect 24568 4711 24584 4745
rect 24518 4677 24584 4711
rect 24518 4643 24534 4677
rect 24568 4643 24584 4677
rect 24518 4609 24584 4643
rect 24518 4575 24534 4609
rect 24568 4575 24584 4609
rect 24518 4541 24584 4575
rect 24518 4507 24534 4541
rect 24568 4507 24584 4541
rect 24518 4473 24584 4507
rect 24518 4439 24534 4473
rect 24568 4439 24584 4473
rect 24518 4405 24584 4439
rect 24518 4371 24534 4405
rect 24568 4371 24584 4405
rect 24518 4337 24584 4371
rect 24518 4303 24534 4337
rect 24568 4303 24584 4337
rect 24518 4269 24584 4303
rect 24518 4235 24534 4269
rect 24568 4235 24584 4269
rect 24518 4201 24584 4235
rect 24518 4167 24534 4201
rect 24568 4167 24584 4201
rect 24518 4126 24584 4167
rect 24614 5085 24680 5126
rect 24614 5051 24630 5085
rect 24664 5051 24680 5085
rect 24614 5017 24680 5051
rect 24614 4983 24630 5017
rect 24664 4983 24680 5017
rect 24614 4949 24680 4983
rect 24614 4915 24630 4949
rect 24664 4915 24680 4949
rect 24614 4881 24680 4915
rect 24614 4847 24630 4881
rect 24664 4847 24680 4881
rect 24614 4813 24680 4847
rect 24614 4779 24630 4813
rect 24664 4779 24680 4813
rect 24614 4745 24680 4779
rect 24614 4711 24630 4745
rect 24664 4711 24680 4745
rect 24614 4677 24680 4711
rect 24614 4643 24630 4677
rect 24664 4643 24680 4677
rect 24614 4609 24680 4643
rect 24614 4575 24630 4609
rect 24664 4575 24680 4609
rect 24614 4541 24680 4575
rect 24614 4507 24630 4541
rect 24664 4507 24680 4541
rect 24614 4473 24680 4507
rect 24614 4439 24630 4473
rect 24664 4439 24680 4473
rect 24614 4405 24680 4439
rect 24614 4371 24630 4405
rect 24664 4371 24680 4405
rect 24614 4337 24680 4371
rect 24614 4303 24630 4337
rect 24664 4303 24680 4337
rect 24614 4269 24680 4303
rect 24614 4235 24630 4269
rect 24664 4235 24680 4269
rect 24614 4201 24680 4235
rect 24614 4167 24630 4201
rect 24664 4167 24680 4201
rect 24614 4126 24680 4167
rect 24710 5085 24776 5126
rect 24710 5051 24726 5085
rect 24760 5051 24776 5085
rect 24710 5017 24776 5051
rect 24710 4983 24726 5017
rect 24760 4983 24776 5017
rect 24710 4949 24776 4983
rect 24710 4915 24726 4949
rect 24760 4915 24776 4949
rect 24710 4881 24776 4915
rect 24710 4847 24726 4881
rect 24760 4847 24776 4881
rect 24710 4813 24776 4847
rect 24710 4779 24726 4813
rect 24760 4779 24776 4813
rect 24710 4745 24776 4779
rect 24710 4711 24726 4745
rect 24760 4711 24776 4745
rect 24710 4677 24776 4711
rect 24710 4643 24726 4677
rect 24760 4643 24776 4677
rect 24710 4609 24776 4643
rect 24710 4575 24726 4609
rect 24760 4575 24776 4609
rect 24710 4541 24776 4575
rect 24710 4507 24726 4541
rect 24760 4507 24776 4541
rect 24710 4473 24776 4507
rect 24710 4439 24726 4473
rect 24760 4439 24776 4473
rect 24710 4405 24776 4439
rect 24710 4371 24726 4405
rect 24760 4371 24776 4405
rect 24710 4337 24776 4371
rect 24710 4303 24726 4337
rect 24760 4303 24776 4337
rect 24710 4269 24776 4303
rect 24710 4235 24726 4269
rect 24760 4235 24776 4269
rect 24710 4201 24776 4235
rect 24710 4167 24726 4201
rect 24760 4167 24776 4201
rect 24710 4126 24776 4167
rect 24806 5085 24872 5126
rect 24806 5051 24822 5085
rect 24856 5051 24872 5085
rect 24806 5017 24872 5051
rect 24806 4983 24822 5017
rect 24856 4983 24872 5017
rect 24806 4949 24872 4983
rect 24806 4915 24822 4949
rect 24856 4915 24872 4949
rect 24806 4881 24872 4915
rect 24806 4847 24822 4881
rect 24856 4847 24872 4881
rect 24806 4813 24872 4847
rect 24806 4779 24822 4813
rect 24856 4779 24872 4813
rect 24806 4745 24872 4779
rect 24806 4711 24822 4745
rect 24856 4711 24872 4745
rect 24806 4677 24872 4711
rect 24806 4643 24822 4677
rect 24856 4643 24872 4677
rect 24806 4609 24872 4643
rect 24806 4575 24822 4609
rect 24856 4575 24872 4609
rect 24806 4541 24872 4575
rect 24806 4507 24822 4541
rect 24856 4507 24872 4541
rect 24806 4473 24872 4507
rect 24806 4439 24822 4473
rect 24856 4439 24872 4473
rect 24806 4405 24872 4439
rect 24806 4371 24822 4405
rect 24856 4371 24872 4405
rect 24806 4337 24872 4371
rect 24806 4303 24822 4337
rect 24856 4303 24872 4337
rect 24806 4269 24872 4303
rect 24806 4235 24822 4269
rect 24856 4235 24872 4269
rect 24806 4201 24872 4235
rect 24806 4167 24822 4201
rect 24856 4167 24872 4201
rect 24806 4126 24872 4167
rect 24902 5085 24964 5126
rect 24902 5051 24918 5085
rect 24952 5051 24964 5085
rect 24902 5017 24964 5051
rect 24902 4983 24918 5017
rect 24952 4983 24964 5017
rect 24902 4949 24964 4983
rect 24902 4915 24918 4949
rect 24952 4915 24964 4949
rect 24902 4881 24964 4915
rect 24902 4847 24918 4881
rect 24952 4847 24964 4881
rect 24902 4813 24964 4847
rect 24902 4779 24918 4813
rect 24952 4779 24964 4813
rect 24902 4745 24964 4779
rect 24902 4711 24918 4745
rect 24952 4711 24964 4745
rect 24902 4677 24964 4711
rect 24902 4643 24918 4677
rect 24952 4643 24964 4677
rect 24902 4609 24964 4643
rect 24902 4575 24918 4609
rect 24952 4575 24964 4609
rect 24902 4541 24964 4575
rect 24902 4507 24918 4541
rect 24952 4507 24964 4541
rect 24902 4473 24964 4507
rect 24902 4439 24918 4473
rect 24952 4439 24964 4473
rect 24902 4405 24964 4439
rect 24902 4371 24918 4405
rect 24952 4371 24964 4405
rect 24902 4337 24964 4371
rect 24902 4303 24918 4337
rect 24952 4303 24964 4337
rect 24902 4269 24964 4303
rect 24902 4235 24918 4269
rect 24952 4235 24964 4269
rect 24902 4201 24964 4235
rect 24902 4167 24918 4201
rect 24952 4167 24964 4201
rect 24902 4126 24964 4167
rect 25150 5079 25212 5120
rect 25150 5045 25162 5079
rect 25196 5045 25212 5079
rect 25150 5011 25212 5045
rect 25150 4977 25162 5011
rect 25196 4977 25212 5011
rect 25150 4943 25212 4977
rect 25150 4909 25162 4943
rect 25196 4909 25212 4943
rect 25150 4875 25212 4909
rect 25150 4841 25162 4875
rect 25196 4841 25212 4875
rect 25150 4807 25212 4841
rect 25150 4773 25162 4807
rect 25196 4773 25212 4807
rect 25150 4739 25212 4773
rect 25150 4705 25162 4739
rect 25196 4705 25212 4739
rect 25150 4671 25212 4705
rect 25150 4637 25162 4671
rect 25196 4637 25212 4671
rect 25150 4603 25212 4637
rect 25150 4569 25162 4603
rect 25196 4569 25212 4603
rect 25150 4535 25212 4569
rect 25150 4501 25162 4535
rect 25196 4501 25212 4535
rect 25150 4467 25212 4501
rect 25150 4433 25162 4467
rect 25196 4433 25212 4467
rect 25150 4399 25212 4433
rect 25150 4365 25162 4399
rect 25196 4365 25212 4399
rect 25150 4331 25212 4365
rect 25150 4297 25162 4331
rect 25196 4297 25212 4331
rect 25150 4263 25212 4297
rect 25150 4229 25162 4263
rect 25196 4229 25212 4263
rect 25150 4195 25212 4229
rect 25150 4161 25162 4195
rect 25196 4161 25212 4195
rect 25150 4120 25212 4161
rect 25242 5079 25308 5120
rect 25242 5045 25258 5079
rect 25292 5045 25308 5079
rect 25242 5011 25308 5045
rect 25242 4977 25258 5011
rect 25292 4977 25308 5011
rect 25242 4943 25308 4977
rect 25242 4909 25258 4943
rect 25292 4909 25308 4943
rect 25242 4875 25308 4909
rect 25242 4841 25258 4875
rect 25292 4841 25308 4875
rect 25242 4807 25308 4841
rect 25242 4773 25258 4807
rect 25292 4773 25308 4807
rect 25242 4739 25308 4773
rect 25242 4705 25258 4739
rect 25292 4705 25308 4739
rect 25242 4671 25308 4705
rect 25242 4637 25258 4671
rect 25292 4637 25308 4671
rect 25242 4603 25308 4637
rect 25242 4569 25258 4603
rect 25292 4569 25308 4603
rect 25242 4535 25308 4569
rect 25242 4501 25258 4535
rect 25292 4501 25308 4535
rect 25242 4467 25308 4501
rect 25242 4433 25258 4467
rect 25292 4433 25308 4467
rect 25242 4399 25308 4433
rect 25242 4365 25258 4399
rect 25292 4365 25308 4399
rect 25242 4331 25308 4365
rect 25242 4297 25258 4331
rect 25292 4297 25308 4331
rect 25242 4263 25308 4297
rect 25242 4229 25258 4263
rect 25292 4229 25308 4263
rect 25242 4195 25308 4229
rect 25242 4161 25258 4195
rect 25292 4161 25308 4195
rect 25242 4120 25308 4161
rect 25338 5079 25404 5120
rect 25338 5045 25354 5079
rect 25388 5045 25404 5079
rect 25338 5011 25404 5045
rect 25338 4977 25354 5011
rect 25388 4977 25404 5011
rect 25338 4943 25404 4977
rect 25338 4909 25354 4943
rect 25388 4909 25404 4943
rect 25338 4875 25404 4909
rect 25338 4841 25354 4875
rect 25388 4841 25404 4875
rect 25338 4807 25404 4841
rect 25338 4773 25354 4807
rect 25388 4773 25404 4807
rect 25338 4739 25404 4773
rect 25338 4705 25354 4739
rect 25388 4705 25404 4739
rect 25338 4671 25404 4705
rect 25338 4637 25354 4671
rect 25388 4637 25404 4671
rect 25338 4603 25404 4637
rect 25338 4569 25354 4603
rect 25388 4569 25404 4603
rect 25338 4535 25404 4569
rect 25338 4501 25354 4535
rect 25388 4501 25404 4535
rect 25338 4467 25404 4501
rect 25338 4433 25354 4467
rect 25388 4433 25404 4467
rect 25338 4399 25404 4433
rect 25338 4365 25354 4399
rect 25388 4365 25404 4399
rect 25338 4331 25404 4365
rect 25338 4297 25354 4331
rect 25388 4297 25404 4331
rect 25338 4263 25404 4297
rect 25338 4229 25354 4263
rect 25388 4229 25404 4263
rect 25338 4195 25404 4229
rect 25338 4161 25354 4195
rect 25388 4161 25404 4195
rect 25338 4120 25404 4161
rect 25434 5079 25500 5120
rect 25434 5045 25450 5079
rect 25484 5045 25500 5079
rect 25434 5011 25500 5045
rect 25434 4977 25450 5011
rect 25484 4977 25500 5011
rect 25434 4943 25500 4977
rect 25434 4909 25450 4943
rect 25484 4909 25500 4943
rect 25434 4875 25500 4909
rect 25434 4841 25450 4875
rect 25484 4841 25500 4875
rect 25434 4807 25500 4841
rect 25434 4773 25450 4807
rect 25484 4773 25500 4807
rect 25434 4739 25500 4773
rect 25434 4705 25450 4739
rect 25484 4705 25500 4739
rect 25434 4671 25500 4705
rect 25434 4637 25450 4671
rect 25484 4637 25500 4671
rect 25434 4603 25500 4637
rect 25434 4569 25450 4603
rect 25484 4569 25500 4603
rect 25434 4535 25500 4569
rect 25434 4501 25450 4535
rect 25484 4501 25500 4535
rect 25434 4467 25500 4501
rect 25434 4433 25450 4467
rect 25484 4433 25500 4467
rect 25434 4399 25500 4433
rect 25434 4365 25450 4399
rect 25484 4365 25500 4399
rect 25434 4331 25500 4365
rect 25434 4297 25450 4331
rect 25484 4297 25500 4331
rect 25434 4263 25500 4297
rect 25434 4229 25450 4263
rect 25484 4229 25500 4263
rect 25434 4195 25500 4229
rect 25434 4161 25450 4195
rect 25484 4161 25500 4195
rect 25434 4120 25500 4161
rect 25530 5079 25596 5120
rect 25530 5045 25546 5079
rect 25580 5045 25596 5079
rect 25530 5011 25596 5045
rect 25530 4977 25546 5011
rect 25580 4977 25596 5011
rect 25530 4943 25596 4977
rect 25530 4909 25546 4943
rect 25580 4909 25596 4943
rect 25530 4875 25596 4909
rect 25530 4841 25546 4875
rect 25580 4841 25596 4875
rect 25530 4807 25596 4841
rect 25530 4773 25546 4807
rect 25580 4773 25596 4807
rect 25530 4739 25596 4773
rect 25530 4705 25546 4739
rect 25580 4705 25596 4739
rect 25530 4671 25596 4705
rect 25530 4637 25546 4671
rect 25580 4637 25596 4671
rect 25530 4603 25596 4637
rect 25530 4569 25546 4603
rect 25580 4569 25596 4603
rect 25530 4535 25596 4569
rect 25530 4501 25546 4535
rect 25580 4501 25596 4535
rect 25530 4467 25596 4501
rect 25530 4433 25546 4467
rect 25580 4433 25596 4467
rect 25530 4399 25596 4433
rect 25530 4365 25546 4399
rect 25580 4365 25596 4399
rect 25530 4331 25596 4365
rect 25530 4297 25546 4331
rect 25580 4297 25596 4331
rect 25530 4263 25596 4297
rect 25530 4229 25546 4263
rect 25580 4229 25596 4263
rect 25530 4195 25596 4229
rect 25530 4161 25546 4195
rect 25580 4161 25596 4195
rect 25530 4120 25596 4161
rect 25626 5079 25692 5120
rect 25626 5045 25642 5079
rect 25676 5045 25692 5079
rect 25626 5011 25692 5045
rect 25626 4977 25642 5011
rect 25676 4977 25692 5011
rect 25626 4943 25692 4977
rect 25626 4909 25642 4943
rect 25676 4909 25692 4943
rect 25626 4875 25692 4909
rect 25626 4841 25642 4875
rect 25676 4841 25692 4875
rect 25626 4807 25692 4841
rect 25626 4773 25642 4807
rect 25676 4773 25692 4807
rect 25626 4739 25692 4773
rect 25626 4705 25642 4739
rect 25676 4705 25692 4739
rect 25626 4671 25692 4705
rect 25626 4637 25642 4671
rect 25676 4637 25692 4671
rect 25626 4603 25692 4637
rect 25626 4569 25642 4603
rect 25676 4569 25692 4603
rect 25626 4535 25692 4569
rect 25626 4501 25642 4535
rect 25676 4501 25692 4535
rect 25626 4467 25692 4501
rect 25626 4433 25642 4467
rect 25676 4433 25692 4467
rect 25626 4399 25692 4433
rect 25626 4365 25642 4399
rect 25676 4365 25692 4399
rect 25626 4331 25692 4365
rect 25626 4297 25642 4331
rect 25676 4297 25692 4331
rect 25626 4263 25692 4297
rect 25626 4229 25642 4263
rect 25676 4229 25692 4263
rect 25626 4195 25692 4229
rect 25626 4161 25642 4195
rect 25676 4161 25692 4195
rect 25626 4120 25692 4161
rect 25722 5079 25788 5120
rect 25722 5045 25738 5079
rect 25772 5045 25788 5079
rect 25722 5011 25788 5045
rect 25722 4977 25738 5011
rect 25772 4977 25788 5011
rect 25722 4943 25788 4977
rect 25722 4909 25738 4943
rect 25772 4909 25788 4943
rect 25722 4875 25788 4909
rect 25722 4841 25738 4875
rect 25772 4841 25788 4875
rect 25722 4807 25788 4841
rect 25722 4773 25738 4807
rect 25772 4773 25788 4807
rect 25722 4739 25788 4773
rect 25722 4705 25738 4739
rect 25772 4705 25788 4739
rect 25722 4671 25788 4705
rect 25722 4637 25738 4671
rect 25772 4637 25788 4671
rect 25722 4603 25788 4637
rect 25722 4569 25738 4603
rect 25772 4569 25788 4603
rect 25722 4535 25788 4569
rect 25722 4501 25738 4535
rect 25772 4501 25788 4535
rect 25722 4467 25788 4501
rect 25722 4433 25738 4467
rect 25772 4433 25788 4467
rect 25722 4399 25788 4433
rect 25722 4365 25738 4399
rect 25772 4365 25788 4399
rect 25722 4331 25788 4365
rect 25722 4297 25738 4331
rect 25772 4297 25788 4331
rect 25722 4263 25788 4297
rect 25722 4229 25738 4263
rect 25772 4229 25788 4263
rect 25722 4195 25788 4229
rect 25722 4161 25738 4195
rect 25772 4161 25788 4195
rect 25722 4120 25788 4161
rect 25818 5079 25884 5120
rect 25818 5045 25834 5079
rect 25868 5045 25884 5079
rect 25818 5011 25884 5045
rect 25818 4977 25834 5011
rect 25868 4977 25884 5011
rect 25818 4943 25884 4977
rect 25818 4909 25834 4943
rect 25868 4909 25884 4943
rect 25818 4875 25884 4909
rect 25818 4841 25834 4875
rect 25868 4841 25884 4875
rect 25818 4807 25884 4841
rect 25818 4773 25834 4807
rect 25868 4773 25884 4807
rect 25818 4739 25884 4773
rect 25818 4705 25834 4739
rect 25868 4705 25884 4739
rect 25818 4671 25884 4705
rect 25818 4637 25834 4671
rect 25868 4637 25884 4671
rect 25818 4603 25884 4637
rect 25818 4569 25834 4603
rect 25868 4569 25884 4603
rect 25818 4535 25884 4569
rect 25818 4501 25834 4535
rect 25868 4501 25884 4535
rect 25818 4467 25884 4501
rect 25818 4433 25834 4467
rect 25868 4433 25884 4467
rect 25818 4399 25884 4433
rect 25818 4365 25834 4399
rect 25868 4365 25884 4399
rect 25818 4331 25884 4365
rect 25818 4297 25834 4331
rect 25868 4297 25884 4331
rect 25818 4263 25884 4297
rect 25818 4229 25834 4263
rect 25868 4229 25884 4263
rect 25818 4195 25884 4229
rect 25818 4161 25834 4195
rect 25868 4161 25884 4195
rect 25818 4120 25884 4161
rect 25914 5079 25980 5120
rect 25914 5045 25930 5079
rect 25964 5045 25980 5079
rect 25914 5011 25980 5045
rect 25914 4977 25930 5011
rect 25964 4977 25980 5011
rect 25914 4943 25980 4977
rect 25914 4909 25930 4943
rect 25964 4909 25980 4943
rect 25914 4875 25980 4909
rect 25914 4841 25930 4875
rect 25964 4841 25980 4875
rect 25914 4807 25980 4841
rect 25914 4773 25930 4807
rect 25964 4773 25980 4807
rect 25914 4739 25980 4773
rect 25914 4705 25930 4739
rect 25964 4705 25980 4739
rect 25914 4671 25980 4705
rect 25914 4637 25930 4671
rect 25964 4637 25980 4671
rect 25914 4603 25980 4637
rect 25914 4569 25930 4603
rect 25964 4569 25980 4603
rect 25914 4535 25980 4569
rect 25914 4501 25930 4535
rect 25964 4501 25980 4535
rect 25914 4467 25980 4501
rect 25914 4433 25930 4467
rect 25964 4433 25980 4467
rect 25914 4399 25980 4433
rect 25914 4365 25930 4399
rect 25964 4365 25980 4399
rect 25914 4331 25980 4365
rect 25914 4297 25930 4331
rect 25964 4297 25980 4331
rect 25914 4263 25980 4297
rect 25914 4229 25930 4263
rect 25964 4229 25980 4263
rect 25914 4195 25980 4229
rect 25914 4161 25930 4195
rect 25964 4161 25980 4195
rect 25914 4120 25980 4161
rect 26010 5079 26076 5120
rect 26010 5045 26026 5079
rect 26060 5045 26076 5079
rect 26010 5011 26076 5045
rect 26010 4977 26026 5011
rect 26060 4977 26076 5011
rect 26010 4943 26076 4977
rect 26010 4909 26026 4943
rect 26060 4909 26076 4943
rect 26010 4875 26076 4909
rect 26010 4841 26026 4875
rect 26060 4841 26076 4875
rect 26010 4807 26076 4841
rect 26010 4773 26026 4807
rect 26060 4773 26076 4807
rect 26010 4739 26076 4773
rect 26010 4705 26026 4739
rect 26060 4705 26076 4739
rect 26010 4671 26076 4705
rect 26010 4637 26026 4671
rect 26060 4637 26076 4671
rect 26010 4603 26076 4637
rect 26010 4569 26026 4603
rect 26060 4569 26076 4603
rect 26010 4535 26076 4569
rect 26010 4501 26026 4535
rect 26060 4501 26076 4535
rect 26010 4467 26076 4501
rect 26010 4433 26026 4467
rect 26060 4433 26076 4467
rect 26010 4399 26076 4433
rect 26010 4365 26026 4399
rect 26060 4365 26076 4399
rect 26010 4331 26076 4365
rect 26010 4297 26026 4331
rect 26060 4297 26076 4331
rect 26010 4263 26076 4297
rect 26010 4229 26026 4263
rect 26060 4229 26076 4263
rect 26010 4195 26076 4229
rect 26010 4161 26026 4195
rect 26060 4161 26076 4195
rect 26010 4120 26076 4161
rect 26106 5079 26172 5120
rect 26106 5045 26122 5079
rect 26156 5045 26172 5079
rect 26106 5011 26172 5045
rect 26106 4977 26122 5011
rect 26156 4977 26172 5011
rect 26106 4943 26172 4977
rect 26106 4909 26122 4943
rect 26156 4909 26172 4943
rect 26106 4875 26172 4909
rect 26106 4841 26122 4875
rect 26156 4841 26172 4875
rect 26106 4807 26172 4841
rect 26106 4773 26122 4807
rect 26156 4773 26172 4807
rect 26106 4739 26172 4773
rect 26106 4705 26122 4739
rect 26156 4705 26172 4739
rect 26106 4671 26172 4705
rect 26106 4637 26122 4671
rect 26156 4637 26172 4671
rect 26106 4603 26172 4637
rect 26106 4569 26122 4603
rect 26156 4569 26172 4603
rect 26106 4535 26172 4569
rect 26106 4501 26122 4535
rect 26156 4501 26172 4535
rect 26106 4467 26172 4501
rect 26106 4433 26122 4467
rect 26156 4433 26172 4467
rect 26106 4399 26172 4433
rect 26106 4365 26122 4399
rect 26156 4365 26172 4399
rect 26106 4331 26172 4365
rect 26106 4297 26122 4331
rect 26156 4297 26172 4331
rect 26106 4263 26172 4297
rect 26106 4229 26122 4263
rect 26156 4229 26172 4263
rect 26106 4195 26172 4229
rect 26106 4161 26122 4195
rect 26156 4161 26172 4195
rect 26106 4120 26172 4161
rect 26202 5079 26268 5120
rect 26202 5045 26218 5079
rect 26252 5045 26268 5079
rect 26202 5011 26268 5045
rect 26202 4977 26218 5011
rect 26252 4977 26268 5011
rect 26202 4943 26268 4977
rect 26202 4909 26218 4943
rect 26252 4909 26268 4943
rect 26202 4875 26268 4909
rect 26202 4841 26218 4875
rect 26252 4841 26268 4875
rect 26202 4807 26268 4841
rect 26202 4773 26218 4807
rect 26252 4773 26268 4807
rect 26202 4739 26268 4773
rect 26202 4705 26218 4739
rect 26252 4705 26268 4739
rect 26202 4671 26268 4705
rect 26202 4637 26218 4671
rect 26252 4637 26268 4671
rect 26202 4603 26268 4637
rect 26202 4569 26218 4603
rect 26252 4569 26268 4603
rect 26202 4535 26268 4569
rect 26202 4501 26218 4535
rect 26252 4501 26268 4535
rect 26202 4467 26268 4501
rect 26202 4433 26218 4467
rect 26252 4433 26268 4467
rect 26202 4399 26268 4433
rect 26202 4365 26218 4399
rect 26252 4365 26268 4399
rect 26202 4331 26268 4365
rect 26202 4297 26218 4331
rect 26252 4297 26268 4331
rect 26202 4263 26268 4297
rect 26202 4229 26218 4263
rect 26252 4229 26268 4263
rect 26202 4195 26268 4229
rect 26202 4161 26218 4195
rect 26252 4161 26268 4195
rect 26202 4120 26268 4161
rect 26298 5079 26364 5120
rect 26298 5045 26314 5079
rect 26348 5045 26364 5079
rect 26298 5011 26364 5045
rect 26298 4977 26314 5011
rect 26348 4977 26364 5011
rect 26298 4943 26364 4977
rect 26298 4909 26314 4943
rect 26348 4909 26364 4943
rect 26298 4875 26364 4909
rect 26298 4841 26314 4875
rect 26348 4841 26364 4875
rect 26298 4807 26364 4841
rect 26298 4773 26314 4807
rect 26348 4773 26364 4807
rect 26298 4739 26364 4773
rect 26298 4705 26314 4739
rect 26348 4705 26364 4739
rect 26298 4671 26364 4705
rect 26298 4637 26314 4671
rect 26348 4637 26364 4671
rect 26298 4603 26364 4637
rect 26298 4569 26314 4603
rect 26348 4569 26364 4603
rect 26298 4535 26364 4569
rect 26298 4501 26314 4535
rect 26348 4501 26364 4535
rect 26298 4467 26364 4501
rect 26298 4433 26314 4467
rect 26348 4433 26364 4467
rect 26298 4399 26364 4433
rect 26298 4365 26314 4399
rect 26348 4365 26364 4399
rect 26298 4331 26364 4365
rect 26298 4297 26314 4331
rect 26348 4297 26364 4331
rect 26298 4263 26364 4297
rect 26298 4229 26314 4263
rect 26348 4229 26364 4263
rect 26298 4195 26364 4229
rect 26298 4161 26314 4195
rect 26348 4161 26364 4195
rect 26298 4120 26364 4161
rect 26394 5079 26460 5120
rect 26394 5045 26410 5079
rect 26444 5045 26460 5079
rect 26394 5011 26460 5045
rect 26394 4977 26410 5011
rect 26444 4977 26460 5011
rect 26394 4943 26460 4977
rect 26394 4909 26410 4943
rect 26444 4909 26460 4943
rect 26394 4875 26460 4909
rect 26394 4841 26410 4875
rect 26444 4841 26460 4875
rect 26394 4807 26460 4841
rect 26394 4773 26410 4807
rect 26444 4773 26460 4807
rect 26394 4739 26460 4773
rect 26394 4705 26410 4739
rect 26444 4705 26460 4739
rect 26394 4671 26460 4705
rect 26394 4637 26410 4671
rect 26444 4637 26460 4671
rect 26394 4603 26460 4637
rect 26394 4569 26410 4603
rect 26444 4569 26460 4603
rect 26394 4535 26460 4569
rect 26394 4501 26410 4535
rect 26444 4501 26460 4535
rect 26394 4467 26460 4501
rect 26394 4433 26410 4467
rect 26444 4433 26460 4467
rect 26394 4399 26460 4433
rect 26394 4365 26410 4399
rect 26444 4365 26460 4399
rect 26394 4331 26460 4365
rect 26394 4297 26410 4331
rect 26444 4297 26460 4331
rect 26394 4263 26460 4297
rect 26394 4229 26410 4263
rect 26444 4229 26460 4263
rect 26394 4195 26460 4229
rect 26394 4161 26410 4195
rect 26444 4161 26460 4195
rect 26394 4120 26460 4161
rect 26490 5079 26556 5120
rect 26490 5045 26506 5079
rect 26540 5045 26556 5079
rect 26490 5011 26556 5045
rect 26490 4977 26506 5011
rect 26540 4977 26556 5011
rect 26490 4943 26556 4977
rect 26490 4909 26506 4943
rect 26540 4909 26556 4943
rect 26490 4875 26556 4909
rect 26490 4841 26506 4875
rect 26540 4841 26556 4875
rect 26490 4807 26556 4841
rect 26490 4773 26506 4807
rect 26540 4773 26556 4807
rect 26490 4739 26556 4773
rect 26490 4705 26506 4739
rect 26540 4705 26556 4739
rect 26490 4671 26556 4705
rect 26490 4637 26506 4671
rect 26540 4637 26556 4671
rect 26490 4603 26556 4637
rect 26490 4569 26506 4603
rect 26540 4569 26556 4603
rect 26490 4535 26556 4569
rect 26490 4501 26506 4535
rect 26540 4501 26556 4535
rect 26490 4467 26556 4501
rect 26490 4433 26506 4467
rect 26540 4433 26556 4467
rect 26490 4399 26556 4433
rect 26490 4365 26506 4399
rect 26540 4365 26556 4399
rect 26490 4331 26556 4365
rect 26490 4297 26506 4331
rect 26540 4297 26556 4331
rect 26490 4263 26556 4297
rect 26490 4229 26506 4263
rect 26540 4229 26556 4263
rect 26490 4195 26556 4229
rect 26490 4161 26506 4195
rect 26540 4161 26556 4195
rect 26490 4120 26556 4161
rect 26586 5079 26648 5120
rect 26586 5045 26602 5079
rect 26636 5045 26648 5079
rect 26586 5011 26648 5045
rect 26586 4977 26602 5011
rect 26636 4977 26648 5011
rect 26586 4943 26648 4977
rect 26586 4909 26602 4943
rect 26636 4909 26648 4943
rect 26586 4875 26648 4909
rect 26586 4841 26602 4875
rect 26636 4841 26648 4875
rect 26586 4807 26648 4841
rect 26586 4773 26602 4807
rect 26636 4773 26648 4807
rect 26586 4739 26648 4773
rect 26586 4705 26602 4739
rect 26636 4705 26648 4739
rect 26586 4671 26648 4705
rect 26586 4637 26602 4671
rect 26636 4637 26648 4671
rect 26586 4603 26648 4637
rect 26586 4569 26602 4603
rect 26636 4569 26648 4603
rect 26586 4535 26648 4569
rect 26586 4501 26602 4535
rect 26636 4501 26648 4535
rect 26586 4467 26648 4501
rect 26586 4433 26602 4467
rect 26636 4433 26648 4467
rect 26586 4399 26648 4433
rect 26586 4365 26602 4399
rect 26636 4365 26648 4399
rect 26586 4331 26648 4365
rect 26586 4297 26602 4331
rect 26636 4297 26648 4331
rect 26586 4263 26648 4297
rect 26586 4229 26602 4263
rect 26636 4229 26648 4263
rect 26586 4195 26648 4229
rect 26586 4161 26602 4195
rect 26636 4161 26648 4195
rect 26586 4120 26648 4161
rect 26814 5073 26876 5114
rect 26814 5039 26826 5073
rect 26860 5039 26876 5073
rect 26814 5005 26876 5039
rect 26814 4971 26826 5005
rect 26860 4971 26876 5005
rect 26814 4937 26876 4971
rect 26814 4903 26826 4937
rect 26860 4903 26876 4937
rect 26814 4869 26876 4903
rect 26814 4835 26826 4869
rect 26860 4835 26876 4869
rect 26814 4801 26876 4835
rect 26814 4767 26826 4801
rect 26860 4767 26876 4801
rect 26814 4733 26876 4767
rect 26814 4699 26826 4733
rect 26860 4699 26876 4733
rect 26814 4665 26876 4699
rect 26814 4631 26826 4665
rect 26860 4631 26876 4665
rect 26814 4597 26876 4631
rect 26814 4563 26826 4597
rect 26860 4563 26876 4597
rect 26814 4529 26876 4563
rect 26814 4495 26826 4529
rect 26860 4495 26876 4529
rect 26814 4461 26876 4495
rect 26814 4427 26826 4461
rect 26860 4427 26876 4461
rect 26814 4393 26876 4427
rect 26814 4359 26826 4393
rect 26860 4359 26876 4393
rect 26814 4325 26876 4359
rect 26814 4291 26826 4325
rect 26860 4291 26876 4325
rect 26814 4257 26876 4291
rect 26814 4223 26826 4257
rect 26860 4223 26876 4257
rect 26814 4189 26876 4223
rect 26814 4155 26826 4189
rect 26860 4155 26876 4189
rect 15694 3926 15756 3957
rect 26814 4114 26876 4155
rect 26906 5073 26972 5114
rect 26906 5039 26922 5073
rect 26956 5039 26972 5073
rect 26906 5005 26972 5039
rect 26906 4971 26922 5005
rect 26956 4971 26972 5005
rect 26906 4937 26972 4971
rect 26906 4903 26922 4937
rect 26956 4903 26972 4937
rect 26906 4869 26972 4903
rect 26906 4835 26922 4869
rect 26956 4835 26972 4869
rect 26906 4801 26972 4835
rect 26906 4767 26922 4801
rect 26956 4767 26972 4801
rect 26906 4733 26972 4767
rect 26906 4699 26922 4733
rect 26956 4699 26972 4733
rect 26906 4665 26972 4699
rect 26906 4631 26922 4665
rect 26956 4631 26972 4665
rect 26906 4597 26972 4631
rect 26906 4563 26922 4597
rect 26956 4563 26972 4597
rect 26906 4529 26972 4563
rect 26906 4495 26922 4529
rect 26956 4495 26972 4529
rect 26906 4461 26972 4495
rect 26906 4427 26922 4461
rect 26956 4427 26972 4461
rect 26906 4393 26972 4427
rect 26906 4359 26922 4393
rect 26956 4359 26972 4393
rect 26906 4325 26972 4359
rect 26906 4291 26922 4325
rect 26956 4291 26972 4325
rect 26906 4257 26972 4291
rect 26906 4223 26922 4257
rect 26956 4223 26972 4257
rect 26906 4189 26972 4223
rect 26906 4155 26922 4189
rect 26956 4155 26972 4189
rect 26906 4114 26972 4155
rect 27002 5073 27068 5114
rect 27002 5039 27018 5073
rect 27052 5039 27068 5073
rect 27002 5005 27068 5039
rect 27002 4971 27018 5005
rect 27052 4971 27068 5005
rect 27002 4937 27068 4971
rect 27002 4903 27018 4937
rect 27052 4903 27068 4937
rect 27002 4869 27068 4903
rect 27002 4835 27018 4869
rect 27052 4835 27068 4869
rect 27002 4801 27068 4835
rect 27002 4767 27018 4801
rect 27052 4767 27068 4801
rect 27002 4733 27068 4767
rect 27002 4699 27018 4733
rect 27052 4699 27068 4733
rect 27002 4665 27068 4699
rect 27002 4631 27018 4665
rect 27052 4631 27068 4665
rect 27002 4597 27068 4631
rect 27002 4563 27018 4597
rect 27052 4563 27068 4597
rect 27002 4529 27068 4563
rect 27002 4495 27018 4529
rect 27052 4495 27068 4529
rect 27002 4461 27068 4495
rect 27002 4427 27018 4461
rect 27052 4427 27068 4461
rect 27002 4393 27068 4427
rect 27002 4359 27018 4393
rect 27052 4359 27068 4393
rect 27002 4325 27068 4359
rect 27002 4291 27018 4325
rect 27052 4291 27068 4325
rect 27002 4257 27068 4291
rect 27002 4223 27018 4257
rect 27052 4223 27068 4257
rect 27002 4189 27068 4223
rect 27002 4155 27018 4189
rect 27052 4155 27068 4189
rect 27002 4114 27068 4155
rect 27098 5073 27164 5114
rect 27098 5039 27114 5073
rect 27148 5039 27164 5073
rect 27098 5005 27164 5039
rect 27098 4971 27114 5005
rect 27148 4971 27164 5005
rect 27098 4937 27164 4971
rect 27098 4903 27114 4937
rect 27148 4903 27164 4937
rect 27098 4869 27164 4903
rect 27098 4835 27114 4869
rect 27148 4835 27164 4869
rect 27098 4801 27164 4835
rect 27098 4767 27114 4801
rect 27148 4767 27164 4801
rect 27098 4733 27164 4767
rect 27098 4699 27114 4733
rect 27148 4699 27164 4733
rect 27098 4665 27164 4699
rect 27098 4631 27114 4665
rect 27148 4631 27164 4665
rect 27098 4597 27164 4631
rect 27098 4563 27114 4597
rect 27148 4563 27164 4597
rect 27098 4529 27164 4563
rect 27098 4495 27114 4529
rect 27148 4495 27164 4529
rect 27098 4461 27164 4495
rect 27098 4427 27114 4461
rect 27148 4427 27164 4461
rect 27098 4393 27164 4427
rect 27098 4359 27114 4393
rect 27148 4359 27164 4393
rect 27098 4325 27164 4359
rect 27098 4291 27114 4325
rect 27148 4291 27164 4325
rect 27098 4257 27164 4291
rect 27098 4223 27114 4257
rect 27148 4223 27164 4257
rect 27098 4189 27164 4223
rect 27098 4155 27114 4189
rect 27148 4155 27164 4189
rect 27098 4114 27164 4155
rect 27194 5073 27260 5114
rect 27194 5039 27210 5073
rect 27244 5039 27260 5073
rect 27194 5005 27260 5039
rect 27194 4971 27210 5005
rect 27244 4971 27260 5005
rect 27194 4937 27260 4971
rect 27194 4903 27210 4937
rect 27244 4903 27260 4937
rect 27194 4869 27260 4903
rect 27194 4835 27210 4869
rect 27244 4835 27260 4869
rect 27194 4801 27260 4835
rect 27194 4767 27210 4801
rect 27244 4767 27260 4801
rect 27194 4733 27260 4767
rect 27194 4699 27210 4733
rect 27244 4699 27260 4733
rect 27194 4665 27260 4699
rect 27194 4631 27210 4665
rect 27244 4631 27260 4665
rect 27194 4597 27260 4631
rect 27194 4563 27210 4597
rect 27244 4563 27260 4597
rect 27194 4529 27260 4563
rect 27194 4495 27210 4529
rect 27244 4495 27260 4529
rect 27194 4461 27260 4495
rect 27194 4427 27210 4461
rect 27244 4427 27260 4461
rect 27194 4393 27260 4427
rect 27194 4359 27210 4393
rect 27244 4359 27260 4393
rect 27194 4325 27260 4359
rect 27194 4291 27210 4325
rect 27244 4291 27260 4325
rect 27194 4257 27260 4291
rect 27194 4223 27210 4257
rect 27244 4223 27260 4257
rect 27194 4189 27260 4223
rect 27194 4155 27210 4189
rect 27244 4155 27260 4189
rect 27194 4114 27260 4155
rect 27290 5073 27356 5114
rect 27290 5039 27306 5073
rect 27340 5039 27356 5073
rect 27290 5005 27356 5039
rect 27290 4971 27306 5005
rect 27340 4971 27356 5005
rect 27290 4937 27356 4971
rect 27290 4903 27306 4937
rect 27340 4903 27356 4937
rect 27290 4869 27356 4903
rect 27290 4835 27306 4869
rect 27340 4835 27356 4869
rect 27290 4801 27356 4835
rect 27290 4767 27306 4801
rect 27340 4767 27356 4801
rect 27290 4733 27356 4767
rect 27290 4699 27306 4733
rect 27340 4699 27356 4733
rect 27290 4665 27356 4699
rect 27290 4631 27306 4665
rect 27340 4631 27356 4665
rect 27290 4597 27356 4631
rect 27290 4563 27306 4597
rect 27340 4563 27356 4597
rect 27290 4529 27356 4563
rect 27290 4495 27306 4529
rect 27340 4495 27356 4529
rect 27290 4461 27356 4495
rect 27290 4427 27306 4461
rect 27340 4427 27356 4461
rect 27290 4393 27356 4427
rect 27290 4359 27306 4393
rect 27340 4359 27356 4393
rect 27290 4325 27356 4359
rect 27290 4291 27306 4325
rect 27340 4291 27356 4325
rect 27290 4257 27356 4291
rect 27290 4223 27306 4257
rect 27340 4223 27356 4257
rect 27290 4189 27356 4223
rect 27290 4155 27306 4189
rect 27340 4155 27356 4189
rect 27290 4114 27356 4155
rect 27386 5073 27452 5114
rect 27386 5039 27402 5073
rect 27436 5039 27452 5073
rect 27386 5005 27452 5039
rect 27386 4971 27402 5005
rect 27436 4971 27452 5005
rect 27386 4937 27452 4971
rect 27386 4903 27402 4937
rect 27436 4903 27452 4937
rect 27386 4869 27452 4903
rect 27386 4835 27402 4869
rect 27436 4835 27452 4869
rect 27386 4801 27452 4835
rect 27386 4767 27402 4801
rect 27436 4767 27452 4801
rect 27386 4733 27452 4767
rect 27386 4699 27402 4733
rect 27436 4699 27452 4733
rect 27386 4665 27452 4699
rect 27386 4631 27402 4665
rect 27436 4631 27452 4665
rect 27386 4597 27452 4631
rect 27386 4563 27402 4597
rect 27436 4563 27452 4597
rect 27386 4529 27452 4563
rect 27386 4495 27402 4529
rect 27436 4495 27452 4529
rect 27386 4461 27452 4495
rect 27386 4427 27402 4461
rect 27436 4427 27452 4461
rect 27386 4393 27452 4427
rect 27386 4359 27402 4393
rect 27436 4359 27452 4393
rect 27386 4325 27452 4359
rect 27386 4291 27402 4325
rect 27436 4291 27452 4325
rect 27386 4257 27452 4291
rect 27386 4223 27402 4257
rect 27436 4223 27452 4257
rect 27386 4189 27452 4223
rect 27386 4155 27402 4189
rect 27436 4155 27452 4189
rect 27386 4114 27452 4155
rect 27482 5073 27548 5114
rect 27482 5039 27498 5073
rect 27532 5039 27548 5073
rect 27482 5005 27548 5039
rect 27482 4971 27498 5005
rect 27532 4971 27548 5005
rect 27482 4937 27548 4971
rect 27482 4903 27498 4937
rect 27532 4903 27548 4937
rect 27482 4869 27548 4903
rect 27482 4835 27498 4869
rect 27532 4835 27548 4869
rect 27482 4801 27548 4835
rect 27482 4767 27498 4801
rect 27532 4767 27548 4801
rect 27482 4733 27548 4767
rect 27482 4699 27498 4733
rect 27532 4699 27548 4733
rect 27482 4665 27548 4699
rect 27482 4631 27498 4665
rect 27532 4631 27548 4665
rect 27482 4597 27548 4631
rect 27482 4563 27498 4597
rect 27532 4563 27548 4597
rect 27482 4529 27548 4563
rect 27482 4495 27498 4529
rect 27532 4495 27548 4529
rect 27482 4461 27548 4495
rect 27482 4427 27498 4461
rect 27532 4427 27548 4461
rect 27482 4393 27548 4427
rect 27482 4359 27498 4393
rect 27532 4359 27548 4393
rect 27482 4325 27548 4359
rect 27482 4291 27498 4325
rect 27532 4291 27548 4325
rect 27482 4257 27548 4291
rect 27482 4223 27498 4257
rect 27532 4223 27548 4257
rect 27482 4189 27548 4223
rect 27482 4155 27498 4189
rect 27532 4155 27548 4189
rect 27482 4114 27548 4155
rect 27578 5073 27644 5114
rect 27578 5039 27594 5073
rect 27628 5039 27644 5073
rect 27578 5005 27644 5039
rect 27578 4971 27594 5005
rect 27628 4971 27644 5005
rect 27578 4937 27644 4971
rect 27578 4903 27594 4937
rect 27628 4903 27644 4937
rect 27578 4869 27644 4903
rect 27578 4835 27594 4869
rect 27628 4835 27644 4869
rect 27578 4801 27644 4835
rect 27578 4767 27594 4801
rect 27628 4767 27644 4801
rect 27578 4733 27644 4767
rect 27578 4699 27594 4733
rect 27628 4699 27644 4733
rect 27578 4665 27644 4699
rect 27578 4631 27594 4665
rect 27628 4631 27644 4665
rect 27578 4597 27644 4631
rect 27578 4563 27594 4597
rect 27628 4563 27644 4597
rect 27578 4529 27644 4563
rect 27578 4495 27594 4529
rect 27628 4495 27644 4529
rect 27578 4461 27644 4495
rect 27578 4427 27594 4461
rect 27628 4427 27644 4461
rect 27578 4393 27644 4427
rect 27578 4359 27594 4393
rect 27628 4359 27644 4393
rect 27578 4325 27644 4359
rect 27578 4291 27594 4325
rect 27628 4291 27644 4325
rect 27578 4257 27644 4291
rect 27578 4223 27594 4257
rect 27628 4223 27644 4257
rect 27578 4189 27644 4223
rect 27578 4155 27594 4189
rect 27628 4155 27644 4189
rect 27578 4114 27644 4155
rect 27674 5073 27740 5114
rect 27674 5039 27690 5073
rect 27724 5039 27740 5073
rect 27674 5005 27740 5039
rect 27674 4971 27690 5005
rect 27724 4971 27740 5005
rect 27674 4937 27740 4971
rect 27674 4903 27690 4937
rect 27724 4903 27740 4937
rect 27674 4869 27740 4903
rect 27674 4835 27690 4869
rect 27724 4835 27740 4869
rect 27674 4801 27740 4835
rect 27674 4767 27690 4801
rect 27724 4767 27740 4801
rect 27674 4733 27740 4767
rect 27674 4699 27690 4733
rect 27724 4699 27740 4733
rect 27674 4665 27740 4699
rect 27674 4631 27690 4665
rect 27724 4631 27740 4665
rect 27674 4597 27740 4631
rect 27674 4563 27690 4597
rect 27724 4563 27740 4597
rect 27674 4529 27740 4563
rect 27674 4495 27690 4529
rect 27724 4495 27740 4529
rect 27674 4461 27740 4495
rect 27674 4427 27690 4461
rect 27724 4427 27740 4461
rect 27674 4393 27740 4427
rect 27674 4359 27690 4393
rect 27724 4359 27740 4393
rect 27674 4325 27740 4359
rect 27674 4291 27690 4325
rect 27724 4291 27740 4325
rect 27674 4257 27740 4291
rect 27674 4223 27690 4257
rect 27724 4223 27740 4257
rect 27674 4189 27740 4223
rect 27674 4155 27690 4189
rect 27724 4155 27740 4189
rect 27674 4114 27740 4155
rect 27770 5073 27836 5114
rect 27770 5039 27786 5073
rect 27820 5039 27836 5073
rect 27770 5005 27836 5039
rect 27770 4971 27786 5005
rect 27820 4971 27836 5005
rect 27770 4937 27836 4971
rect 27770 4903 27786 4937
rect 27820 4903 27836 4937
rect 27770 4869 27836 4903
rect 27770 4835 27786 4869
rect 27820 4835 27836 4869
rect 27770 4801 27836 4835
rect 27770 4767 27786 4801
rect 27820 4767 27836 4801
rect 27770 4733 27836 4767
rect 27770 4699 27786 4733
rect 27820 4699 27836 4733
rect 27770 4665 27836 4699
rect 27770 4631 27786 4665
rect 27820 4631 27836 4665
rect 27770 4597 27836 4631
rect 27770 4563 27786 4597
rect 27820 4563 27836 4597
rect 27770 4529 27836 4563
rect 27770 4495 27786 4529
rect 27820 4495 27836 4529
rect 27770 4461 27836 4495
rect 27770 4427 27786 4461
rect 27820 4427 27836 4461
rect 27770 4393 27836 4427
rect 27770 4359 27786 4393
rect 27820 4359 27836 4393
rect 27770 4325 27836 4359
rect 27770 4291 27786 4325
rect 27820 4291 27836 4325
rect 27770 4257 27836 4291
rect 27770 4223 27786 4257
rect 27820 4223 27836 4257
rect 27770 4189 27836 4223
rect 27770 4155 27786 4189
rect 27820 4155 27836 4189
rect 27770 4114 27836 4155
rect 27866 5073 27932 5114
rect 27866 5039 27882 5073
rect 27916 5039 27932 5073
rect 27866 5005 27932 5039
rect 27866 4971 27882 5005
rect 27916 4971 27932 5005
rect 27866 4937 27932 4971
rect 27866 4903 27882 4937
rect 27916 4903 27932 4937
rect 27866 4869 27932 4903
rect 27866 4835 27882 4869
rect 27916 4835 27932 4869
rect 27866 4801 27932 4835
rect 27866 4767 27882 4801
rect 27916 4767 27932 4801
rect 27866 4733 27932 4767
rect 27866 4699 27882 4733
rect 27916 4699 27932 4733
rect 27866 4665 27932 4699
rect 27866 4631 27882 4665
rect 27916 4631 27932 4665
rect 27866 4597 27932 4631
rect 27866 4563 27882 4597
rect 27916 4563 27932 4597
rect 27866 4529 27932 4563
rect 27866 4495 27882 4529
rect 27916 4495 27932 4529
rect 27866 4461 27932 4495
rect 27866 4427 27882 4461
rect 27916 4427 27932 4461
rect 27866 4393 27932 4427
rect 27866 4359 27882 4393
rect 27916 4359 27932 4393
rect 27866 4325 27932 4359
rect 27866 4291 27882 4325
rect 27916 4291 27932 4325
rect 27866 4257 27932 4291
rect 27866 4223 27882 4257
rect 27916 4223 27932 4257
rect 27866 4189 27932 4223
rect 27866 4155 27882 4189
rect 27916 4155 27932 4189
rect 27866 4114 27932 4155
rect 27962 5073 28028 5114
rect 27962 5039 27978 5073
rect 28012 5039 28028 5073
rect 27962 5005 28028 5039
rect 27962 4971 27978 5005
rect 28012 4971 28028 5005
rect 27962 4937 28028 4971
rect 27962 4903 27978 4937
rect 28012 4903 28028 4937
rect 27962 4869 28028 4903
rect 27962 4835 27978 4869
rect 28012 4835 28028 4869
rect 27962 4801 28028 4835
rect 27962 4767 27978 4801
rect 28012 4767 28028 4801
rect 27962 4733 28028 4767
rect 27962 4699 27978 4733
rect 28012 4699 28028 4733
rect 27962 4665 28028 4699
rect 27962 4631 27978 4665
rect 28012 4631 28028 4665
rect 27962 4597 28028 4631
rect 27962 4563 27978 4597
rect 28012 4563 28028 4597
rect 27962 4529 28028 4563
rect 27962 4495 27978 4529
rect 28012 4495 28028 4529
rect 27962 4461 28028 4495
rect 27962 4427 27978 4461
rect 28012 4427 28028 4461
rect 27962 4393 28028 4427
rect 27962 4359 27978 4393
rect 28012 4359 28028 4393
rect 27962 4325 28028 4359
rect 27962 4291 27978 4325
rect 28012 4291 28028 4325
rect 27962 4257 28028 4291
rect 27962 4223 27978 4257
rect 28012 4223 28028 4257
rect 27962 4189 28028 4223
rect 27962 4155 27978 4189
rect 28012 4155 28028 4189
rect 27962 4114 28028 4155
rect 28058 5073 28124 5114
rect 28058 5039 28074 5073
rect 28108 5039 28124 5073
rect 28058 5005 28124 5039
rect 28058 4971 28074 5005
rect 28108 4971 28124 5005
rect 28058 4937 28124 4971
rect 28058 4903 28074 4937
rect 28108 4903 28124 4937
rect 28058 4869 28124 4903
rect 28058 4835 28074 4869
rect 28108 4835 28124 4869
rect 28058 4801 28124 4835
rect 28058 4767 28074 4801
rect 28108 4767 28124 4801
rect 28058 4733 28124 4767
rect 28058 4699 28074 4733
rect 28108 4699 28124 4733
rect 28058 4665 28124 4699
rect 28058 4631 28074 4665
rect 28108 4631 28124 4665
rect 28058 4597 28124 4631
rect 28058 4563 28074 4597
rect 28108 4563 28124 4597
rect 28058 4529 28124 4563
rect 28058 4495 28074 4529
rect 28108 4495 28124 4529
rect 28058 4461 28124 4495
rect 28058 4427 28074 4461
rect 28108 4427 28124 4461
rect 28058 4393 28124 4427
rect 28058 4359 28074 4393
rect 28108 4359 28124 4393
rect 28058 4325 28124 4359
rect 28058 4291 28074 4325
rect 28108 4291 28124 4325
rect 28058 4257 28124 4291
rect 28058 4223 28074 4257
rect 28108 4223 28124 4257
rect 28058 4189 28124 4223
rect 28058 4155 28074 4189
rect 28108 4155 28124 4189
rect 28058 4114 28124 4155
rect 28154 5073 28220 5114
rect 28154 5039 28170 5073
rect 28204 5039 28220 5073
rect 28154 5005 28220 5039
rect 28154 4971 28170 5005
rect 28204 4971 28220 5005
rect 28154 4937 28220 4971
rect 28154 4903 28170 4937
rect 28204 4903 28220 4937
rect 28154 4869 28220 4903
rect 28154 4835 28170 4869
rect 28204 4835 28220 4869
rect 28154 4801 28220 4835
rect 28154 4767 28170 4801
rect 28204 4767 28220 4801
rect 28154 4733 28220 4767
rect 28154 4699 28170 4733
rect 28204 4699 28220 4733
rect 28154 4665 28220 4699
rect 28154 4631 28170 4665
rect 28204 4631 28220 4665
rect 28154 4597 28220 4631
rect 28154 4563 28170 4597
rect 28204 4563 28220 4597
rect 28154 4529 28220 4563
rect 28154 4495 28170 4529
rect 28204 4495 28220 4529
rect 28154 4461 28220 4495
rect 28154 4427 28170 4461
rect 28204 4427 28220 4461
rect 28154 4393 28220 4427
rect 28154 4359 28170 4393
rect 28204 4359 28220 4393
rect 28154 4325 28220 4359
rect 28154 4291 28170 4325
rect 28204 4291 28220 4325
rect 28154 4257 28220 4291
rect 28154 4223 28170 4257
rect 28204 4223 28220 4257
rect 28154 4189 28220 4223
rect 28154 4155 28170 4189
rect 28204 4155 28220 4189
rect 28154 4114 28220 4155
rect 28250 5073 28316 5114
rect 28250 5039 28266 5073
rect 28300 5039 28316 5073
rect 28250 5005 28316 5039
rect 28250 4971 28266 5005
rect 28300 4971 28316 5005
rect 28250 4937 28316 4971
rect 28250 4903 28266 4937
rect 28300 4903 28316 4937
rect 28250 4869 28316 4903
rect 28250 4835 28266 4869
rect 28300 4835 28316 4869
rect 28250 4801 28316 4835
rect 28250 4767 28266 4801
rect 28300 4767 28316 4801
rect 28250 4733 28316 4767
rect 28250 4699 28266 4733
rect 28300 4699 28316 4733
rect 28250 4665 28316 4699
rect 28250 4631 28266 4665
rect 28300 4631 28316 4665
rect 28250 4597 28316 4631
rect 28250 4563 28266 4597
rect 28300 4563 28316 4597
rect 28250 4529 28316 4563
rect 28250 4495 28266 4529
rect 28300 4495 28316 4529
rect 28250 4461 28316 4495
rect 28250 4427 28266 4461
rect 28300 4427 28316 4461
rect 28250 4393 28316 4427
rect 28250 4359 28266 4393
rect 28300 4359 28316 4393
rect 28250 4325 28316 4359
rect 28250 4291 28266 4325
rect 28300 4291 28316 4325
rect 28250 4257 28316 4291
rect 28250 4223 28266 4257
rect 28300 4223 28316 4257
rect 28250 4189 28316 4223
rect 28250 4155 28266 4189
rect 28300 4155 28316 4189
rect 28250 4114 28316 4155
rect 28346 5073 28412 5114
rect 28346 5039 28362 5073
rect 28396 5039 28412 5073
rect 28346 5005 28412 5039
rect 28346 4971 28362 5005
rect 28396 4971 28412 5005
rect 28346 4937 28412 4971
rect 28346 4903 28362 4937
rect 28396 4903 28412 4937
rect 28346 4869 28412 4903
rect 28346 4835 28362 4869
rect 28396 4835 28412 4869
rect 28346 4801 28412 4835
rect 28346 4767 28362 4801
rect 28396 4767 28412 4801
rect 28346 4733 28412 4767
rect 28346 4699 28362 4733
rect 28396 4699 28412 4733
rect 28346 4665 28412 4699
rect 28346 4631 28362 4665
rect 28396 4631 28412 4665
rect 28346 4597 28412 4631
rect 28346 4563 28362 4597
rect 28396 4563 28412 4597
rect 28346 4529 28412 4563
rect 28346 4495 28362 4529
rect 28396 4495 28412 4529
rect 28346 4461 28412 4495
rect 28346 4427 28362 4461
rect 28396 4427 28412 4461
rect 28346 4393 28412 4427
rect 28346 4359 28362 4393
rect 28396 4359 28412 4393
rect 28346 4325 28412 4359
rect 28346 4291 28362 4325
rect 28396 4291 28412 4325
rect 28346 4257 28412 4291
rect 28346 4223 28362 4257
rect 28396 4223 28412 4257
rect 28346 4189 28412 4223
rect 28346 4155 28362 4189
rect 28396 4155 28412 4189
rect 28346 4114 28412 4155
rect 28442 5073 28508 5114
rect 28442 5039 28458 5073
rect 28492 5039 28508 5073
rect 28442 5005 28508 5039
rect 28442 4971 28458 5005
rect 28492 4971 28508 5005
rect 28442 4937 28508 4971
rect 28442 4903 28458 4937
rect 28492 4903 28508 4937
rect 28442 4869 28508 4903
rect 28442 4835 28458 4869
rect 28492 4835 28508 4869
rect 28442 4801 28508 4835
rect 28442 4767 28458 4801
rect 28492 4767 28508 4801
rect 28442 4733 28508 4767
rect 28442 4699 28458 4733
rect 28492 4699 28508 4733
rect 28442 4665 28508 4699
rect 28442 4631 28458 4665
rect 28492 4631 28508 4665
rect 28442 4597 28508 4631
rect 28442 4563 28458 4597
rect 28492 4563 28508 4597
rect 28442 4529 28508 4563
rect 28442 4495 28458 4529
rect 28492 4495 28508 4529
rect 28442 4461 28508 4495
rect 28442 4427 28458 4461
rect 28492 4427 28508 4461
rect 28442 4393 28508 4427
rect 28442 4359 28458 4393
rect 28492 4359 28508 4393
rect 28442 4325 28508 4359
rect 28442 4291 28458 4325
rect 28492 4291 28508 4325
rect 28442 4257 28508 4291
rect 28442 4223 28458 4257
rect 28492 4223 28508 4257
rect 28442 4189 28508 4223
rect 28442 4155 28458 4189
rect 28492 4155 28508 4189
rect 28442 4114 28508 4155
rect 28538 5073 28604 5114
rect 28538 5039 28554 5073
rect 28588 5039 28604 5073
rect 28538 5005 28604 5039
rect 28538 4971 28554 5005
rect 28588 4971 28604 5005
rect 28538 4937 28604 4971
rect 28538 4903 28554 4937
rect 28588 4903 28604 4937
rect 28538 4869 28604 4903
rect 28538 4835 28554 4869
rect 28588 4835 28604 4869
rect 28538 4801 28604 4835
rect 28538 4767 28554 4801
rect 28588 4767 28604 4801
rect 28538 4733 28604 4767
rect 28538 4699 28554 4733
rect 28588 4699 28604 4733
rect 28538 4665 28604 4699
rect 28538 4631 28554 4665
rect 28588 4631 28604 4665
rect 28538 4597 28604 4631
rect 28538 4563 28554 4597
rect 28588 4563 28604 4597
rect 28538 4529 28604 4563
rect 28538 4495 28554 4529
rect 28588 4495 28604 4529
rect 28538 4461 28604 4495
rect 28538 4427 28554 4461
rect 28588 4427 28604 4461
rect 28538 4393 28604 4427
rect 28538 4359 28554 4393
rect 28588 4359 28604 4393
rect 28538 4325 28604 4359
rect 28538 4291 28554 4325
rect 28588 4291 28604 4325
rect 28538 4257 28604 4291
rect 28538 4223 28554 4257
rect 28588 4223 28604 4257
rect 28538 4189 28604 4223
rect 28538 4155 28554 4189
rect 28588 4155 28604 4189
rect 28538 4114 28604 4155
rect 28634 5073 28700 5114
rect 28634 5039 28650 5073
rect 28684 5039 28700 5073
rect 28634 5005 28700 5039
rect 28634 4971 28650 5005
rect 28684 4971 28700 5005
rect 28634 4937 28700 4971
rect 28634 4903 28650 4937
rect 28684 4903 28700 4937
rect 28634 4869 28700 4903
rect 28634 4835 28650 4869
rect 28684 4835 28700 4869
rect 28634 4801 28700 4835
rect 28634 4767 28650 4801
rect 28684 4767 28700 4801
rect 28634 4733 28700 4767
rect 28634 4699 28650 4733
rect 28684 4699 28700 4733
rect 28634 4665 28700 4699
rect 28634 4631 28650 4665
rect 28684 4631 28700 4665
rect 28634 4597 28700 4631
rect 28634 4563 28650 4597
rect 28684 4563 28700 4597
rect 28634 4529 28700 4563
rect 28634 4495 28650 4529
rect 28684 4495 28700 4529
rect 28634 4461 28700 4495
rect 28634 4427 28650 4461
rect 28684 4427 28700 4461
rect 28634 4393 28700 4427
rect 28634 4359 28650 4393
rect 28684 4359 28700 4393
rect 28634 4325 28700 4359
rect 28634 4291 28650 4325
rect 28684 4291 28700 4325
rect 28634 4257 28700 4291
rect 28634 4223 28650 4257
rect 28684 4223 28700 4257
rect 28634 4189 28700 4223
rect 28634 4155 28650 4189
rect 28684 4155 28700 4189
rect 28634 4114 28700 4155
rect 28730 5073 28792 5114
rect 28730 5039 28746 5073
rect 28780 5039 28792 5073
rect 28730 5005 28792 5039
rect 28730 4971 28746 5005
rect 28780 4971 28792 5005
rect 28730 4937 28792 4971
rect 28730 4903 28746 4937
rect 28780 4903 28792 4937
rect 28730 4869 28792 4903
rect 28730 4835 28746 4869
rect 28780 4835 28792 4869
rect 28730 4801 28792 4835
rect 28730 4767 28746 4801
rect 28780 4767 28792 4801
rect 28730 4733 28792 4767
rect 28730 4699 28746 4733
rect 28780 4699 28792 4733
rect 28730 4665 28792 4699
rect 28730 4631 28746 4665
rect 28780 4631 28792 4665
rect 28730 4597 28792 4631
rect 28730 4563 28746 4597
rect 28780 4563 28792 4597
rect 28730 4529 28792 4563
rect 28730 4495 28746 4529
rect 28780 4495 28792 4529
rect 28730 4461 28792 4495
rect 28730 4427 28746 4461
rect 28780 4427 28792 4461
rect 28730 4393 28792 4427
rect 28730 4359 28746 4393
rect 28780 4359 28792 4393
rect 28730 4325 28792 4359
rect 28730 4291 28746 4325
rect 28780 4291 28792 4325
rect 28730 4257 28792 4291
rect 28730 4223 28746 4257
rect 28780 4223 28792 4257
rect 28730 4189 28792 4223
rect 28730 4155 28746 4189
rect 28780 4155 28792 4189
rect 28730 4114 28792 4155
rect -4830 3677 -4768 3711
rect -4830 3643 -4814 3677
rect -4780 3643 -4768 3677
rect -4830 3609 -4768 3643
rect -4830 3575 -4814 3609
rect -4780 3575 -4768 3609
rect -4830 3541 -4768 3575
rect -4830 3507 -4814 3541
rect -4780 3507 -4768 3541
rect -4830 3466 -4768 3507
<< ndiffc >>
rect 16686 3459 16720 3493
rect 16686 3391 16720 3425
rect 16686 3323 16720 3357
rect 16686 3255 16720 3289
rect -1686 3161 -1652 3195
rect -1686 3093 -1652 3127
rect -23492 2779 -23458 2813
rect -23492 2711 -23458 2745
rect -23492 2643 -23458 2677
rect -23492 2575 -23458 2609
rect -23492 2507 -23458 2541
rect -23492 2439 -23458 2473
rect -23492 2371 -23458 2405
rect -23492 2303 -23458 2337
rect -23492 2235 -23458 2269
rect -23492 2167 -23458 2201
rect -23492 2099 -23458 2133
rect -23492 2031 -23458 2065
rect -23492 1963 -23458 1997
rect -23492 1895 -23458 1929
rect -23396 2779 -23362 2813
rect -23396 2711 -23362 2745
rect -23396 2643 -23362 2677
rect -23396 2575 -23362 2609
rect -23396 2507 -23362 2541
rect -23396 2439 -23362 2473
rect -23396 2371 -23362 2405
rect -23396 2303 -23362 2337
rect -23396 2235 -23362 2269
rect -23396 2167 -23362 2201
rect -23396 2099 -23362 2133
rect -23396 2031 -23362 2065
rect -23396 1963 -23362 1997
rect -23396 1895 -23362 1929
rect -23300 2779 -23266 2813
rect -23300 2711 -23266 2745
rect -23300 2643 -23266 2677
rect -23300 2575 -23266 2609
rect -23300 2507 -23266 2541
rect -23300 2439 -23266 2473
rect -23300 2371 -23266 2405
rect -23300 2303 -23266 2337
rect -23300 2235 -23266 2269
rect -23300 2167 -23266 2201
rect -23300 2099 -23266 2133
rect -23300 2031 -23266 2065
rect -23300 1963 -23266 1997
rect -23300 1895 -23266 1929
rect -23204 2779 -23170 2813
rect -23204 2711 -23170 2745
rect -23204 2643 -23170 2677
rect -23204 2575 -23170 2609
rect -23204 2507 -23170 2541
rect -23204 2439 -23170 2473
rect -23204 2371 -23170 2405
rect -23204 2303 -23170 2337
rect -23204 2235 -23170 2269
rect -23204 2167 -23170 2201
rect -23204 2099 -23170 2133
rect -23204 2031 -23170 2065
rect -23204 1963 -23170 1997
rect -23204 1895 -23170 1929
rect -23108 2779 -23074 2813
rect -23108 2711 -23074 2745
rect -23108 2643 -23074 2677
rect -23108 2575 -23074 2609
rect -23108 2507 -23074 2541
rect -23108 2439 -23074 2473
rect -23108 2371 -23074 2405
rect -23108 2303 -23074 2337
rect -23108 2235 -23074 2269
rect -23108 2167 -23074 2201
rect -23108 2099 -23074 2133
rect -23108 2031 -23074 2065
rect -23108 1963 -23074 1997
rect -23108 1895 -23074 1929
rect -23012 2779 -22978 2813
rect -23012 2711 -22978 2745
rect -23012 2643 -22978 2677
rect -23012 2575 -22978 2609
rect -23012 2507 -22978 2541
rect -23012 2439 -22978 2473
rect -23012 2371 -22978 2405
rect -23012 2303 -22978 2337
rect -23012 2235 -22978 2269
rect -23012 2167 -22978 2201
rect -23012 2099 -22978 2133
rect -23012 2031 -22978 2065
rect -23012 1963 -22978 1997
rect -23012 1895 -22978 1929
rect -22916 2779 -22882 2813
rect -22916 2711 -22882 2745
rect -22916 2643 -22882 2677
rect -22916 2575 -22882 2609
rect -22916 2507 -22882 2541
rect -22916 2439 -22882 2473
rect -22916 2371 -22882 2405
rect -22916 2303 -22882 2337
rect -22916 2235 -22882 2269
rect -22916 2167 -22882 2201
rect -22916 2099 -22882 2133
rect -22916 2031 -22882 2065
rect -22916 1963 -22882 1997
rect -22916 1895 -22882 1929
rect -22820 2779 -22786 2813
rect -22820 2711 -22786 2745
rect -22820 2643 -22786 2677
rect -22820 2575 -22786 2609
rect -22820 2507 -22786 2541
rect -22820 2439 -22786 2473
rect -22820 2371 -22786 2405
rect -22820 2303 -22786 2337
rect -22820 2235 -22786 2269
rect -22820 2167 -22786 2201
rect -22820 2099 -22786 2133
rect -22820 2031 -22786 2065
rect -22820 1963 -22786 1997
rect -22820 1895 -22786 1929
rect -22724 2779 -22690 2813
rect -22724 2711 -22690 2745
rect -22724 2643 -22690 2677
rect -22724 2575 -22690 2609
rect -22724 2507 -22690 2541
rect -22724 2439 -22690 2473
rect -22724 2371 -22690 2405
rect -22724 2303 -22690 2337
rect -22724 2235 -22690 2269
rect -22724 2167 -22690 2201
rect -22724 2099 -22690 2133
rect -22724 2031 -22690 2065
rect -22724 1963 -22690 1997
rect -22724 1895 -22690 1929
rect -22628 2779 -22594 2813
rect -22628 2711 -22594 2745
rect -22628 2643 -22594 2677
rect -22628 2575 -22594 2609
rect -22628 2507 -22594 2541
rect -22628 2439 -22594 2473
rect -22628 2371 -22594 2405
rect -22628 2303 -22594 2337
rect -22628 2235 -22594 2269
rect -22628 2167 -22594 2201
rect -22628 2099 -22594 2133
rect -22628 2031 -22594 2065
rect -22628 1963 -22594 1997
rect -22628 1895 -22594 1929
rect -22532 2779 -22498 2813
rect -22532 2711 -22498 2745
rect -22532 2643 -22498 2677
rect -22532 2575 -22498 2609
rect -22532 2507 -22498 2541
rect -22532 2439 -22498 2473
rect -22532 2371 -22498 2405
rect -22532 2303 -22498 2337
rect -22532 2235 -22498 2269
rect -22532 2167 -22498 2201
rect -22532 2099 -22498 2133
rect -22532 2031 -22498 2065
rect -22532 1963 -22498 1997
rect -22532 1895 -22498 1929
rect -22436 2779 -22402 2813
rect -22436 2711 -22402 2745
rect -22436 2643 -22402 2677
rect -22436 2575 -22402 2609
rect -22436 2507 -22402 2541
rect -22436 2439 -22402 2473
rect -22436 2371 -22402 2405
rect -22436 2303 -22402 2337
rect -22436 2235 -22402 2269
rect -22436 2167 -22402 2201
rect -22436 2099 -22402 2133
rect -22436 2031 -22402 2065
rect -22436 1963 -22402 1997
rect -22436 1895 -22402 1929
rect -22340 2779 -22306 2813
rect -22340 2711 -22306 2745
rect -22340 2643 -22306 2677
rect -22340 2575 -22306 2609
rect -22340 2507 -22306 2541
rect -22340 2439 -22306 2473
rect -22340 2371 -22306 2405
rect -22340 2303 -22306 2337
rect -22340 2235 -22306 2269
rect -22340 2167 -22306 2201
rect -22340 2099 -22306 2133
rect -22340 2031 -22306 2065
rect -22340 1963 -22306 1997
rect -22340 1895 -22306 1929
rect -22244 2779 -22210 2813
rect -22244 2711 -22210 2745
rect -22244 2643 -22210 2677
rect -22244 2575 -22210 2609
rect -22244 2507 -22210 2541
rect -22244 2439 -22210 2473
rect -22244 2371 -22210 2405
rect -22244 2303 -22210 2337
rect -22244 2235 -22210 2269
rect -22244 2167 -22210 2201
rect -22244 2099 -22210 2133
rect -22244 2031 -22210 2065
rect -22244 1963 -22210 1997
rect -22244 1895 -22210 1929
rect -22148 2779 -22114 2813
rect -22148 2711 -22114 2745
rect -22148 2643 -22114 2677
rect -22148 2575 -22114 2609
rect -22148 2507 -22114 2541
rect -22148 2439 -22114 2473
rect -22148 2371 -22114 2405
rect -22148 2303 -22114 2337
rect -22148 2235 -22114 2269
rect -22148 2167 -22114 2201
rect -22148 2099 -22114 2133
rect -22148 2031 -22114 2065
rect -22148 1963 -22114 1997
rect -22148 1895 -22114 1929
rect -22052 2779 -22018 2813
rect -22052 2711 -22018 2745
rect -22052 2643 -22018 2677
rect -22052 2575 -22018 2609
rect -22052 2507 -22018 2541
rect -22052 2439 -22018 2473
rect -22052 2371 -22018 2405
rect -22052 2303 -22018 2337
rect -22052 2235 -22018 2269
rect -22052 2167 -22018 2201
rect -22052 2099 -22018 2133
rect -22052 2031 -22018 2065
rect -22052 1963 -22018 1997
rect -22052 1895 -22018 1929
rect -21956 2779 -21922 2813
rect -21956 2711 -21922 2745
rect -21956 2643 -21922 2677
rect -21956 2575 -21922 2609
rect -21956 2507 -21922 2541
rect -21956 2439 -21922 2473
rect -21956 2371 -21922 2405
rect -21956 2303 -21922 2337
rect -21956 2235 -21922 2269
rect -21956 2167 -21922 2201
rect -21956 2099 -21922 2133
rect -21956 2031 -21922 2065
rect -21956 1963 -21922 1997
rect -21956 1895 -21922 1929
rect -21860 2779 -21826 2813
rect -21860 2711 -21826 2745
rect -21860 2643 -21826 2677
rect -21860 2575 -21826 2609
rect -21860 2507 -21826 2541
rect -21860 2439 -21826 2473
rect -21860 2371 -21826 2405
rect -21860 2303 -21826 2337
rect -21860 2235 -21826 2269
rect -21860 2167 -21826 2201
rect -21860 2099 -21826 2133
rect -21860 2031 -21826 2065
rect -21860 1963 -21826 1997
rect -21860 1895 -21826 1929
rect -21764 2779 -21730 2813
rect -21764 2711 -21730 2745
rect -21764 2643 -21730 2677
rect -21764 2575 -21730 2609
rect -21764 2507 -21730 2541
rect -21764 2439 -21730 2473
rect -21764 2371 -21730 2405
rect -21764 2303 -21730 2337
rect -21764 2235 -21730 2269
rect -21764 2167 -21730 2201
rect -21764 2099 -21730 2133
rect -21764 2031 -21730 2065
rect -21764 1963 -21730 1997
rect -21764 1895 -21730 1929
rect -21668 2779 -21634 2813
rect -21668 2711 -21634 2745
rect -21668 2643 -21634 2677
rect -21668 2575 -21634 2609
rect -21668 2507 -21634 2541
rect -21668 2439 -21634 2473
rect -21668 2371 -21634 2405
rect -21668 2303 -21634 2337
rect -21668 2235 -21634 2269
rect -21668 2167 -21634 2201
rect -21668 2099 -21634 2133
rect -21668 2031 -21634 2065
rect -21668 1963 -21634 1997
rect -21668 1895 -21634 1929
rect -21572 2779 -21538 2813
rect -21572 2711 -21538 2745
rect -21572 2643 -21538 2677
rect -21572 2575 -21538 2609
rect -21572 2507 -21538 2541
rect -21572 2439 -21538 2473
rect -21572 2371 -21538 2405
rect -21572 2303 -21538 2337
rect -21572 2235 -21538 2269
rect -21572 2167 -21538 2201
rect -21572 2099 -21538 2133
rect -21572 2031 -21538 2065
rect -21572 1963 -21538 1997
rect -21572 1895 -21538 1929
rect -21344 2771 -21310 2805
rect -21344 2703 -21310 2737
rect -21344 2635 -21310 2669
rect -21344 2567 -21310 2601
rect -21344 2499 -21310 2533
rect -21344 2431 -21310 2465
rect -21344 2363 -21310 2397
rect -21344 2295 -21310 2329
rect -21344 2227 -21310 2261
rect -21344 2159 -21310 2193
rect -21344 2091 -21310 2125
rect -21344 2023 -21310 2057
rect -21344 1955 -21310 1989
rect -21344 1887 -21310 1921
rect -21248 2771 -21214 2805
rect -21248 2703 -21214 2737
rect -21248 2635 -21214 2669
rect -21248 2567 -21214 2601
rect -21248 2499 -21214 2533
rect -21248 2431 -21214 2465
rect -21248 2363 -21214 2397
rect -21248 2295 -21214 2329
rect -21248 2227 -21214 2261
rect -21248 2159 -21214 2193
rect -21248 2091 -21214 2125
rect -21248 2023 -21214 2057
rect -21248 1955 -21214 1989
rect -21248 1887 -21214 1921
rect -21152 2771 -21118 2805
rect -21152 2703 -21118 2737
rect -21152 2635 -21118 2669
rect -21152 2567 -21118 2601
rect -21152 2499 -21118 2533
rect -21152 2431 -21118 2465
rect -21152 2363 -21118 2397
rect -21152 2295 -21118 2329
rect -21152 2227 -21118 2261
rect -21152 2159 -21118 2193
rect -21152 2091 -21118 2125
rect -21152 2023 -21118 2057
rect -21152 1955 -21118 1989
rect -21152 1887 -21118 1921
rect -21056 2771 -21022 2805
rect -21056 2703 -21022 2737
rect -21056 2635 -21022 2669
rect -21056 2567 -21022 2601
rect -21056 2499 -21022 2533
rect -21056 2431 -21022 2465
rect -21056 2363 -21022 2397
rect -21056 2295 -21022 2329
rect -21056 2227 -21022 2261
rect -21056 2159 -21022 2193
rect -21056 2091 -21022 2125
rect -21056 2023 -21022 2057
rect -21056 1955 -21022 1989
rect -21056 1887 -21022 1921
rect -20960 2771 -20926 2805
rect -20960 2703 -20926 2737
rect -20960 2635 -20926 2669
rect -20960 2567 -20926 2601
rect -20960 2499 -20926 2533
rect -20960 2431 -20926 2465
rect -20960 2363 -20926 2397
rect -20960 2295 -20926 2329
rect -20960 2227 -20926 2261
rect -20960 2159 -20926 2193
rect -20960 2091 -20926 2125
rect -20960 2023 -20926 2057
rect -20960 1955 -20926 1989
rect -20960 1887 -20926 1921
rect -20864 2771 -20830 2805
rect -20864 2703 -20830 2737
rect -20864 2635 -20830 2669
rect -20864 2567 -20830 2601
rect -20864 2499 -20830 2533
rect -20864 2431 -20830 2465
rect -20864 2363 -20830 2397
rect -20864 2295 -20830 2329
rect -20864 2227 -20830 2261
rect -20864 2159 -20830 2193
rect -20864 2091 -20830 2125
rect -20864 2023 -20830 2057
rect -20864 1955 -20830 1989
rect -20864 1887 -20830 1921
rect -20768 2771 -20734 2805
rect -20768 2703 -20734 2737
rect -20768 2635 -20734 2669
rect -20768 2567 -20734 2601
rect -20768 2499 -20734 2533
rect -20768 2431 -20734 2465
rect -20768 2363 -20734 2397
rect -20768 2295 -20734 2329
rect -20768 2227 -20734 2261
rect -20768 2159 -20734 2193
rect -20768 2091 -20734 2125
rect -20768 2023 -20734 2057
rect -20768 1955 -20734 1989
rect -20768 1887 -20734 1921
rect -20672 2771 -20638 2805
rect -20672 2703 -20638 2737
rect -20672 2635 -20638 2669
rect -20672 2567 -20638 2601
rect -20672 2499 -20638 2533
rect -20672 2431 -20638 2465
rect -20672 2363 -20638 2397
rect -20672 2295 -20638 2329
rect -20672 2227 -20638 2261
rect -20672 2159 -20638 2193
rect -20672 2091 -20638 2125
rect -20672 2023 -20638 2057
rect -20672 1955 -20638 1989
rect -20672 1887 -20638 1921
rect -20576 2771 -20542 2805
rect -20576 2703 -20542 2737
rect -20576 2635 -20542 2669
rect -20576 2567 -20542 2601
rect -20576 2499 -20542 2533
rect -20576 2431 -20542 2465
rect -20576 2363 -20542 2397
rect -20576 2295 -20542 2329
rect -20576 2227 -20542 2261
rect -20576 2159 -20542 2193
rect -20576 2091 -20542 2125
rect -20576 2023 -20542 2057
rect -20576 1955 -20542 1989
rect -20576 1887 -20542 1921
rect -20480 2771 -20446 2805
rect -20480 2703 -20446 2737
rect -20480 2635 -20446 2669
rect -20480 2567 -20446 2601
rect -20480 2499 -20446 2533
rect -20480 2431 -20446 2465
rect -20480 2363 -20446 2397
rect -20480 2295 -20446 2329
rect -20480 2227 -20446 2261
rect -20480 2159 -20446 2193
rect -20480 2091 -20446 2125
rect -20480 2023 -20446 2057
rect -20480 1955 -20446 1989
rect -20480 1887 -20446 1921
rect -20384 2771 -20350 2805
rect -20384 2703 -20350 2737
rect -20384 2635 -20350 2669
rect -20384 2567 -20350 2601
rect -20384 2499 -20350 2533
rect -20384 2431 -20350 2465
rect -20384 2363 -20350 2397
rect -20384 2295 -20350 2329
rect -20384 2227 -20350 2261
rect -20384 2159 -20350 2193
rect -20384 2091 -20350 2125
rect -20384 2023 -20350 2057
rect -20384 1955 -20350 1989
rect -20384 1887 -20350 1921
rect -20288 2771 -20254 2805
rect -20288 2703 -20254 2737
rect -20288 2635 -20254 2669
rect -20288 2567 -20254 2601
rect -20288 2499 -20254 2533
rect -20288 2431 -20254 2465
rect -20288 2363 -20254 2397
rect -20288 2295 -20254 2329
rect -20288 2227 -20254 2261
rect -20288 2159 -20254 2193
rect -20288 2091 -20254 2125
rect -20288 2023 -20254 2057
rect -20288 1955 -20254 1989
rect -20288 1887 -20254 1921
rect -20192 2771 -20158 2805
rect -20192 2703 -20158 2737
rect -20192 2635 -20158 2669
rect -20192 2567 -20158 2601
rect -20192 2499 -20158 2533
rect -20192 2431 -20158 2465
rect -20192 2363 -20158 2397
rect -20192 2295 -20158 2329
rect -20192 2227 -20158 2261
rect -20192 2159 -20158 2193
rect -20192 2091 -20158 2125
rect -20192 2023 -20158 2057
rect -20192 1955 -20158 1989
rect -20192 1887 -20158 1921
rect -20096 2771 -20062 2805
rect -20096 2703 -20062 2737
rect -20096 2635 -20062 2669
rect -20096 2567 -20062 2601
rect -20096 2499 -20062 2533
rect -20096 2431 -20062 2465
rect -20096 2363 -20062 2397
rect -20096 2295 -20062 2329
rect -20096 2227 -20062 2261
rect -20096 2159 -20062 2193
rect -20096 2091 -20062 2125
rect -20096 2023 -20062 2057
rect -20096 1955 -20062 1989
rect -20096 1887 -20062 1921
rect -20000 2771 -19966 2805
rect -20000 2703 -19966 2737
rect -20000 2635 -19966 2669
rect -20000 2567 -19966 2601
rect -20000 2499 -19966 2533
rect -20000 2431 -19966 2465
rect -20000 2363 -19966 2397
rect -20000 2295 -19966 2329
rect -20000 2227 -19966 2261
rect -20000 2159 -19966 2193
rect -20000 2091 -19966 2125
rect -20000 2023 -19966 2057
rect -20000 1955 -19966 1989
rect -20000 1887 -19966 1921
rect -19904 2771 -19870 2805
rect -19904 2703 -19870 2737
rect -19904 2635 -19870 2669
rect -19904 2567 -19870 2601
rect -19904 2499 -19870 2533
rect -19904 2431 -19870 2465
rect -19904 2363 -19870 2397
rect -19904 2295 -19870 2329
rect -19904 2227 -19870 2261
rect -19904 2159 -19870 2193
rect -19904 2091 -19870 2125
rect -19904 2023 -19870 2057
rect -19904 1955 -19870 1989
rect -19904 1887 -19870 1921
rect -19666 2775 -19632 2809
rect -19666 2707 -19632 2741
rect -19666 2639 -19632 2673
rect -19666 2571 -19632 2605
rect -19666 2503 -19632 2537
rect -19666 2435 -19632 2469
rect -19666 2367 -19632 2401
rect -19666 2299 -19632 2333
rect -19666 2231 -19632 2265
rect -19666 2163 -19632 2197
rect -19666 2095 -19632 2129
rect -19666 2027 -19632 2061
rect -19666 1959 -19632 1993
rect -19666 1891 -19632 1925
rect -19570 2775 -19536 2809
rect -19570 2707 -19536 2741
rect -19570 2639 -19536 2673
rect -19570 2571 -19536 2605
rect -19570 2503 -19536 2537
rect -19570 2435 -19536 2469
rect -19570 2367 -19536 2401
rect -19570 2299 -19536 2333
rect -19570 2231 -19536 2265
rect -19570 2163 -19536 2197
rect -19570 2095 -19536 2129
rect -19570 2027 -19536 2061
rect -19570 1959 -19536 1993
rect -19570 1891 -19536 1925
rect -19474 2775 -19440 2809
rect -19474 2707 -19440 2741
rect -19474 2639 -19440 2673
rect -19474 2571 -19440 2605
rect -19474 2503 -19440 2537
rect -19474 2435 -19440 2469
rect -19474 2367 -19440 2401
rect -19474 2299 -19440 2333
rect -19474 2231 -19440 2265
rect -19474 2163 -19440 2197
rect -19474 2095 -19440 2129
rect -19474 2027 -19440 2061
rect -19474 1959 -19440 1993
rect -19474 1891 -19440 1925
rect -19378 2775 -19344 2809
rect -19378 2707 -19344 2741
rect -19378 2639 -19344 2673
rect -19378 2571 -19344 2605
rect -19378 2503 -19344 2537
rect -19378 2435 -19344 2469
rect -19378 2367 -19344 2401
rect -19378 2299 -19344 2333
rect -19378 2231 -19344 2265
rect -19378 2163 -19344 2197
rect -19378 2095 -19344 2129
rect -19378 2027 -19344 2061
rect -19378 1959 -19344 1993
rect -19378 1891 -19344 1925
rect -19282 2775 -19248 2809
rect -19282 2707 -19248 2741
rect -19282 2639 -19248 2673
rect -19282 2571 -19248 2605
rect -19282 2503 -19248 2537
rect -19282 2435 -19248 2469
rect -19282 2367 -19248 2401
rect -19282 2299 -19248 2333
rect -19282 2231 -19248 2265
rect -19282 2163 -19248 2197
rect -19282 2095 -19248 2129
rect -19282 2027 -19248 2061
rect -19282 1959 -19248 1993
rect -19282 1891 -19248 1925
rect -19186 2775 -19152 2809
rect -19186 2707 -19152 2741
rect -19186 2639 -19152 2673
rect -19186 2571 -19152 2605
rect -19186 2503 -19152 2537
rect -19186 2435 -19152 2469
rect -19186 2367 -19152 2401
rect -19186 2299 -19152 2333
rect -19186 2231 -19152 2265
rect -19186 2163 -19152 2197
rect -19186 2095 -19152 2129
rect -19186 2027 -19152 2061
rect -19186 1959 -19152 1993
rect -19186 1891 -19152 1925
rect -19090 2775 -19056 2809
rect -19090 2707 -19056 2741
rect -19090 2639 -19056 2673
rect -19090 2571 -19056 2605
rect -19090 2503 -19056 2537
rect -19090 2435 -19056 2469
rect -19090 2367 -19056 2401
rect -19090 2299 -19056 2333
rect -19090 2231 -19056 2265
rect -19090 2163 -19056 2197
rect -19090 2095 -19056 2129
rect -19090 2027 -19056 2061
rect -19090 1959 -19056 1993
rect -19090 1891 -19056 1925
rect -18994 2775 -18960 2809
rect -18994 2707 -18960 2741
rect -18994 2639 -18960 2673
rect -18994 2571 -18960 2605
rect -18994 2503 -18960 2537
rect -18994 2435 -18960 2469
rect -18994 2367 -18960 2401
rect -18994 2299 -18960 2333
rect -18994 2231 -18960 2265
rect -18994 2163 -18960 2197
rect -18994 2095 -18960 2129
rect -18994 2027 -18960 2061
rect -18994 1959 -18960 1993
rect -18994 1891 -18960 1925
rect -18898 2775 -18864 2809
rect -18898 2707 -18864 2741
rect -18898 2639 -18864 2673
rect -18898 2571 -18864 2605
rect -18898 2503 -18864 2537
rect -18898 2435 -18864 2469
rect -18898 2367 -18864 2401
rect -18898 2299 -18864 2333
rect -18898 2231 -18864 2265
rect -18898 2163 -18864 2197
rect -18898 2095 -18864 2129
rect -18898 2027 -18864 2061
rect -18898 1959 -18864 1993
rect -18898 1891 -18864 1925
rect -18802 2775 -18768 2809
rect -18802 2707 -18768 2741
rect -18802 2639 -18768 2673
rect -18802 2571 -18768 2605
rect -18802 2503 -18768 2537
rect -18802 2435 -18768 2469
rect -18802 2367 -18768 2401
rect -18802 2299 -18768 2333
rect -18802 2231 -18768 2265
rect -18802 2163 -18768 2197
rect -18802 2095 -18768 2129
rect -18802 2027 -18768 2061
rect -18802 1959 -18768 1993
rect -18802 1891 -18768 1925
rect -18706 2775 -18672 2809
rect -18706 2707 -18672 2741
rect -18706 2639 -18672 2673
rect -18706 2571 -18672 2605
rect -18706 2503 -18672 2537
rect -18706 2435 -18672 2469
rect -18706 2367 -18672 2401
rect -18706 2299 -18672 2333
rect -18706 2231 -18672 2265
rect -18706 2163 -18672 2197
rect -18706 2095 -18672 2129
rect -18706 2027 -18672 2061
rect -18706 1959 -18672 1993
rect -18706 1891 -18672 1925
rect -18494 2785 -18460 2819
rect -18494 2717 -18460 2751
rect -18494 2649 -18460 2683
rect -18494 2581 -18460 2615
rect -18494 2513 -18460 2547
rect -18494 2445 -18460 2479
rect -18494 2377 -18460 2411
rect -18494 2309 -18460 2343
rect -18494 2241 -18460 2275
rect -18494 2173 -18460 2207
rect -18494 2105 -18460 2139
rect -18494 2037 -18460 2071
rect -18494 1969 -18460 2003
rect -18494 1901 -18460 1935
rect -18398 2785 -18364 2819
rect -18398 2717 -18364 2751
rect -18398 2649 -18364 2683
rect -18398 2581 -18364 2615
rect -18398 2513 -18364 2547
rect -18398 2445 -18364 2479
rect -18398 2377 -18364 2411
rect -18398 2309 -18364 2343
rect -18398 2241 -18364 2275
rect -18398 2173 -18364 2207
rect -18398 2105 -18364 2139
rect -18398 2037 -18364 2071
rect -18398 1969 -18364 2003
rect -18398 1901 -18364 1935
rect -18302 2785 -18268 2819
rect -18302 2717 -18268 2751
rect -18302 2649 -18268 2683
rect -18302 2581 -18268 2615
rect -18302 2513 -18268 2547
rect -18302 2445 -18268 2479
rect -18302 2377 -18268 2411
rect -18302 2309 -18268 2343
rect -18302 2241 -18268 2275
rect -18302 2173 -18268 2207
rect -18302 2105 -18268 2139
rect -18302 2037 -18268 2071
rect -18302 1969 -18268 2003
rect -18302 1901 -18268 1935
rect -18206 2785 -18172 2819
rect -18206 2717 -18172 2751
rect -18206 2649 -18172 2683
rect -18206 2581 -18172 2615
rect -18206 2513 -18172 2547
rect -18206 2445 -18172 2479
rect -18206 2377 -18172 2411
rect -18206 2309 -18172 2343
rect -18206 2241 -18172 2275
rect -18206 2173 -18172 2207
rect -18206 2105 -18172 2139
rect -18206 2037 -18172 2071
rect -18206 1969 -18172 2003
rect -18206 1901 -18172 1935
rect -18110 2785 -18076 2819
rect -18110 2717 -18076 2751
rect -18110 2649 -18076 2683
rect -18110 2581 -18076 2615
rect -18110 2513 -18076 2547
rect -18110 2445 -18076 2479
rect -18110 2377 -18076 2411
rect -18110 2309 -18076 2343
rect -18110 2241 -18076 2275
rect -18110 2173 -18076 2207
rect -18110 2105 -18076 2139
rect -18110 2037 -18076 2071
rect -18110 1969 -18076 2003
rect -18110 1901 -18076 1935
rect -18014 2785 -17980 2819
rect -18014 2717 -17980 2751
rect -18014 2649 -17980 2683
rect -18014 2581 -17980 2615
rect -18014 2513 -17980 2547
rect -18014 2445 -17980 2479
rect -18014 2377 -17980 2411
rect -18014 2309 -17980 2343
rect -18014 2241 -17980 2275
rect -18014 2173 -17980 2207
rect -18014 2105 -17980 2139
rect -18014 2037 -17980 2071
rect -18014 1969 -17980 2003
rect -18014 1901 -17980 1935
rect -16662 2791 -16628 2825
rect -16662 2723 -16628 2757
rect -16662 2655 -16628 2689
rect -16662 2587 -16628 2621
rect -16662 2519 -16628 2553
rect -16662 2451 -16628 2485
rect -16662 2383 -16628 2417
rect -16662 2315 -16628 2349
rect -16662 2247 -16628 2281
rect -16662 2179 -16628 2213
rect -16662 2111 -16628 2145
rect -16662 2043 -16628 2077
rect -16662 1975 -16628 2009
rect -16662 1907 -16628 1941
rect -16566 2791 -16532 2825
rect -16566 2723 -16532 2757
rect -16566 2655 -16532 2689
rect -16566 2587 -16532 2621
rect -16566 2519 -16532 2553
rect -16566 2451 -16532 2485
rect -16566 2383 -16532 2417
rect -16566 2315 -16532 2349
rect -16566 2247 -16532 2281
rect -16566 2179 -16532 2213
rect -16566 2111 -16532 2145
rect -16566 2043 -16532 2077
rect -16566 1975 -16532 2009
rect -16566 1907 -16532 1941
rect -16470 2791 -16436 2825
rect -16470 2723 -16436 2757
rect -16470 2655 -16436 2689
rect -16470 2587 -16436 2621
rect -16470 2519 -16436 2553
rect -16470 2451 -16436 2485
rect -16470 2383 -16436 2417
rect -16470 2315 -16436 2349
rect -16470 2247 -16436 2281
rect -16470 2179 -16436 2213
rect -16470 2111 -16436 2145
rect -16470 2043 -16436 2077
rect -16470 1975 -16436 2009
rect -16470 1907 -16436 1941
rect -16374 2791 -16340 2825
rect -16374 2723 -16340 2757
rect -16374 2655 -16340 2689
rect -16374 2587 -16340 2621
rect -16374 2519 -16340 2553
rect -16374 2451 -16340 2485
rect -16374 2383 -16340 2417
rect -16374 2315 -16340 2349
rect -16374 2247 -16340 2281
rect -16374 2179 -16340 2213
rect -16374 2111 -16340 2145
rect -16374 2043 -16340 2077
rect -16374 1975 -16340 2009
rect -16374 1907 -16340 1941
rect -16278 2791 -16244 2825
rect -16278 2723 -16244 2757
rect -16278 2655 -16244 2689
rect -16278 2587 -16244 2621
rect -16278 2519 -16244 2553
rect -16278 2451 -16244 2485
rect -16278 2383 -16244 2417
rect -16278 2315 -16244 2349
rect -16278 2247 -16244 2281
rect -16278 2179 -16244 2213
rect -16278 2111 -16244 2145
rect -16278 2043 -16244 2077
rect -16278 1975 -16244 2009
rect -16278 1907 -16244 1941
rect -16182 2791 -16148 2825
rect -16182 2723 -16148 2757
rect -16182 2655 -16148 2689
rect -16182 2587 -16148 2621
rect -16182 2519 -16148 2553
rect -16182 2451 -16148 2485
rect -16182 2383 -16148 2417
rect -16182 2315 -16148 2349
rect -16182 2247 -16148 2281
rect -16182 2179 -16148 2213
rect -16182 2111 -16148 2145
rect -16182 2043 -16148 2077
rect -16182 1975 -16148 2009
rect -16182 1907 -16148 1941
rect -16086 2791 -16052 2825
rect -16086 2723 -16052 2757
rect -16086 2655 -16052 2689
rect -16086 2587 -16052 2621
rect -16086 2519 -16052 2553
rect -16086 2451 -16052 2485
rect -16086 2383 -16052 2417
rect -16086 2315 -16052 2349
rect -16086 2247 -16052 2281
rect -16086 2179 -16052 2213
rect -16086 2111 -16052 2145
rect -16086 2043 -16052 2077
rect -16086 1975 -16052 2009
rect -16086 1907 -16052 1941
rect -15990 2791 -15956 2825
rect -15990 2723 -15956 2757
rect -15990 2655 -15956 2689
rect -15990 2587 -15956 2621
rect -15990 2519 -15956 2553
rect -15990 2451 -15956 2485
rect -15990 2383 -15956 2417
rect -15990 2315 -15956 2349
rect -15990 2247 -15956 2281
rect -15990 2179 -15956 2213
rect -15990 2111 -15956 2145
rect -15990 2043 -15956 2077
rect -15990 1975 -15956 2009
rect -15990 1907 -15956 1941
rect -15894 2791 -15860 2825
rect -15894 2723 -15860 2757
rect -15894 2655 -15860 2689
rect -15894 2587 -15860 2621
rect -15894 2519 -15860 2553
rect -15894 2451 -15860 2485
rect -15894 2383 -15860 2417
rect -15894 2315 -15860 2349
rect -15894 2247 -15860 2281
rect -15894 2179 -15860 2213
rect -15894 2111 -15860 2145
rect -15894 2043 -15860 2077
rect -15894 1975 -15860 2009
rect -15894 1907 -15860 1941
rect -15798 2791 -15764 2825
rect -15798 2723 -15764 2757
rect -15798 2655 -15764 2689
rect -15798 2587 -15764 2621
rect -15798 2519 -15764 2553
rect -15798 2451 -15764 2485
rect -15798 2383 -15764 2417
rect -15798 2315 -15764 2349
rect -15798 2247 -15764 2281
rect -15798 2179 -15764 2213
rect -15798 2111 -15764 2145
rect -15798 2043 -15764 2077
rect -15798 1975 -15764 2009
rect -15798 1907 -15764 1941
rect -15702 2791 -15668 2825
rect -15702 2723 -15668 2757
rect -15702 2655 -15668 2689
rect -15702 2587 -15668 2621
rect -15702 2519 -15668 2553
rect -15702 2451 -15668 2485
rect -15702 2383 -15668 2417
rect -15702 2315 -15668 2349
rect -15702 2247 -15668 2281
rect -15702 2179 -15668 2213
rect -15702 2111 -15668 2145
rect -15702 2043 -15668 2077
rect -15702 1975 -15668 2009
rect -15702 1907 -15668 1941
rect -15606 2791 -15572 2825
rect -15606 2723 -15572 2757
rect -15606 2655 -15572 2689
rect -15606 2587 -15572 2621
rect -15606 2519 -15572 2553
rect -15606 2451 -15572 2485
rect -15606 2383 -15572 2417
rect -15606 2315 -15572 2349
rect -15606 2247 -15572 2281
rect -15606 2179 -15572 2213
rect -15606 2111 -15572 2145
rect -15606 2043 -15572 2077
rect -15606 1975 -15572 2009
rect -15606 1907 -15572 1941
rect -15510 2791 -15476 2825
rect -15510 2723 -15476 2757
rect -15510 2655 -15476 2689
rect -15510 2587 -15476 2621
rect -15510 2519 -15476 2553
rect -15510 2451 -15476 2485
rect -15510 2383 -15476 2417
rect -15510 2315 -15476 2349
rect -15510 2247 -15476 2281
rect -15510 2179 -15476 2213
rect -15510 2111 -15476 2145
rect -15510 2043 -15476 2077
rect -15510 1975 -15476 2009
rect -15510 1907 -15476 1941
rect -15414 2791 -15380 2825
rect -15414 2723 -15380 2757
rect -15414 2655 -15380 2689
rect -15414 2587 -15380 2621
rect -15414 2519 -15380 2553
rect -15414 2451 -15380 2485
rect -15414 2383 -15380 2417
rect -15414 2315 -15380 2349
rect -15414 2247 -15380 2281
rect -15414 2179 -15380 2213
rect -15414 2111 -15380 2145
rect -15414 2043 -15380 2077
rect -15414 1975 -15380 2009
rect -15414 1907 -15380 1941
rect -15318 2791 -15284 2825
rect -15318 2723 -15284 2757
rect -15318 2655 -15284 2689
rect -15318 2587 -15284 2621
rect -15318 2519 -15284 2553
rect -15318 2451 -15284 2485
rect -15318 2383 -15284 2417
rect -15318 2315 -15284 2349
rect -15318 2247 -15284 2281
rect -15318 2179 -15284 2213
rect -15318 2111 -15284 2145
rect -15318 2043 -15284 2077
rect -15318 1975 -15284 2009
rect -15318 1907 -15284 1941
rect -15222 2791 -15188 2825
rect -15222 2723 -15188 2757
rect -15222 2655 -15188 2689
rect -15222 2587 -15188 2621
rect -15222 2519 -15188 2553
rect -15222 2451 -15188 2485
rect -15222 2383 -15188 2417
rect -15222 2315 -15188 2349
rect -15222 2247 -15188 2281
rect -15222 2179 -15188 2213
rect -15222 2111 -15188 2145
rect -15222 2043 -15188 2077
rect -15222 1975 -15188 2009
rect -15222 1907 -15188 1941
rect -15126 2791 -15092 2825
rect -15126 2723 -15092 2757
rect -15126 2655 -15092 2689
rect -15126 2587 -15092 2621
rect -15126 2519 -15092 2553
rect -15126 2451 -15092 2485
rect -15126 2383 -15092 2417
rect -15126 2315 -15092 2349
rect -15126 2247 -15092 2281
rect -15126 2179 -15092 2213
rect -15126 2111 -15092 2145
rect -15126 2043 -15092 2077
rect -15126 1975 -15092 2009
rect -15126 1907 -15092 1941
rect -15030 2791 -14996 2825
rect -15030 2723 -14996 2757
rect -15030 2655 -14996 2689
rect -15030 2587 -14996 2621
rect -15030 2519 -14996 2553
rect -15030 2451 -14996 2485
rect -15030 2383 -14996 2417
rect -15030 2315 -14996 2349
rect -15030 2247 -14996 2281
rect -15030 2179 -14996 2213
rect -15030 2111 -14996 2145
rect -15030 2043 -14996 2077
rect -15030 1975 -14996 2009
rect -15030 1907 -14996 1941
rect -14934 2791 -14900 2825
rect -14934 2723 -14900 2757
rect -14934 2655 -14900 2689
rect -14934 2587 -14900 2621
rect -14934 2519 -14900 2553
rect -14934 2451 -14900 2485
rect -14934 2383 -14900 2417
rect -14934 2315 -14900 2349
rect -14934 2247 -14900 2281
rect -14934 2179 -14900 2213
rect -14934 2111 -14900 2145
rect -14934 2043 -14900 2077
rect -14934 1975 -14900 2009
rect -14934 1907 -14900 1941
rect -14838 2791 -14804 2825
rect -14838 2723 -14804 2757
rect -14838 2655 -14804 2689
rect -14838 2587 -14804 2621
rect -14838 2519 -14804 2553
rect -14838 2451 -14804 2485
rect -14838 2383 -14804 2417
rect -14838 2315 -14804 2349
rect -14838 2247 -14804 2281
rect -14838 2179 -14804 2213
rect -14838 2111 -14804 2145
rect -14838 2043 -14804 2077
rect -14838 1975 -14804 2009
rect -14838 1907 -14804 1941
rect -1686 3025 -1652 3059
rect -1686 2957 -1652 2991
rect -14742 2791 -14708 2825
rect -14742 2723 -14708 2757
rect -14742 2655 -14708 2689
rect -14742 2587 -14708 2621
rect -14742 2519 -14708 2553
rect -14742 2451 -14708 2485
rect -14742 2383 -14708 2417
rect -14742 2315 -14708 2349
rect -14742 2247 -14708 2281
rect -14742 2179 -14708 2213
rect -14742 2111 -14708 2145
rect -14742 2043 -14708 2077
rect -14742 1975 -14708 2009
rect -14742 1907 -14708 1941
rect -14514 2783 -14480 2817
rect -14514 2715 -14480 2749
rect -14514 2647 -14480 2681
rect -14514 2579 -14480 2613
rect -14514 2511 -14480 2545
rect -14514 2443 -14480 2477
rect -14514 2375 -14480 2409
rect -14514 2307 -14480 2341
rect -14514 2239 -14480 2273
rect -14514 2171 -14480 2205
rect -14514 2103 -14480 2137
rect -14514 2035 -14480 2069
rect -14514 1967 -14480 2001
rect -14514 1899 -14480 1933
rect -14418 2783 -14384 2817
rect -14418 2715 -14384 2749
rect -14418 2647 -14384 2681
rect -14418 2579 -14384 2613
rect -14418 2511 -14384 2545
rect -14418 2443 -14384 2477
rect -14418 2375 -14384 2409
rect -14418 2307 -14384 2341
rect -14418 2239 -14384 2273
rect -14418 2171 -14384 2205
rect -14418 2103 -14384 2137
rect -14418 2035 -14384 2069
rect -14418 1967 -14384 2001
rect -14418 1899 -14384 1933
rect -14322 2783 -14288 2817
rect -14322 2715 -14288 2749
rect -14322 2647 -14288 2681
rect -14322 2579 -14288 2613
rect -14322 2511 -14288 2545
rect -14322 2443 -14288 2477
rect -14322 2375 -14288 2409
rect -14322 2307 -14288 2341
rect -14322 2239 -14288 2273
rect -14322 2171 -14288 2205
rect -14322 2103 -14288 2137
rect -14322 2035 -14288 2069
rect -14322 1967 -14288 2001
rect -14322 1899 -14288 1933
rect -14226 2783 -14192 2817
rect -14226 2715 -14192 2749
rect -14226 2647 -14192 2681
rect -14226 2579 -14192 2613
rect -14226 2511 -14192 2545
rect -14226 2443 -14192 2477
rect -14226 2375 -14192 2409
rect -14226 2307 -14192 2341
rect -14226 2239 -14192 2273
rect -14226 2171 -14192 2205
rect -14226 2103 -14192 2137
rect -14226 2035 -14192 2069
rect -14226 1967 -14192 2001
rect -14226 1899 -14192 1933
rect -14130 2783 -14096 2817
rect -14130 2715 -14096 2749
rect -14130 2647 -14096 2681
rect -14130 2579 -14096 2613
rect -14130 2511 -14096 2545
rect -14130 2443 -14096 2477
rect -14130 2375 -14096 2409
rect -14130 2307 -14096 2341
rect -14130 2239 -14096 2273
rect -14130 2171 -14096 2205
rect -14130 2103 -14096 2137
rect -14130 2035 -14096 2069
rect -14130 1967 -14096 2001
rect -14130 1899 -14096 1933
rect -14034 2783 -14000 2817
rect -14034 2715 -14000 2749
rect -14034 2647 -14000 2681
rect -14034 2579 -14000 2613
rect -14034 2511 -14000 2545
rect -14034 2443 -14000 2477
rect -14034 2375 -14000 2409
rect -14034 2307 -14000 2341
rect -14034 2239 -14000 2273
rect -14034 2171 -14000 2205
rect -14034 2103 -14000 2137
rect -14034 2035 -14000 2069
rect -14034 1967 -14000 2001
rect -14034 1899 -14000 1933
rect -13938 2783 -13904 2817
rect -13938 2715 -13904 2749
rect -13938 2647 -13904 2681
rect -13938 2579 -13904 2613
rect -13938 2511 -13904 2545
rect -13938 2443 -13904 2477
rect -13938 2375 -13904 2409
rect -13938 2307 -13904 2341
rect -13938 2239 -13904 2273
rect -13938 2171 -13904 2205
rect -13938 2103 -13904 2137
rect -13938 2035 -13904 2069
rect -13938 1967 -13904 2001
rect -13938 1899 -13904 1933
rect -13842 2783 -13808 2817
rect -13842 2715 -13808 2749
rect -13842 2647 -13808 2681
rect -13842 2579 -13808 2613
rect -13842 2511 -13808 2545
rect -13842 2443 -13808 2477
rect -13842 2375 -13808 2409
rect -13842 2307 -13808 2341
rect -13842 2239 -13808 2273
rect -13842 2171 -13808 2205
rect -13842 2103 -13808 2137
rect -13842 2035 -13808 2069
rect -13842 1967 -13808 2001
rect -13842 1899 -13808 1933
rect -13746 2783 -13712 2817
rect -13746 2715 -13712 2749
rect -13746 2647 -13712 2681
rect -13746 2579 -13712 2613
rect -13746 2511 -13712 2545
rect -13746 2443 -13712 2477
rect -13746 2375 -13712 2409
rect -13746 2307 -13712 2341
rect -13746 2239 -13712 2273
rect -13746 2171 -13712 2205
rect -13746 2103 -13712 2137
rect -13746 2035 -13712 2069
rect -13746 1967 -13712 2001
rect -13746 1899 -13712 1933
rect -13650 2783 -13616 2817
rect -13650 2715 -13616 2749
rect -13650 2647 -13616 2681
rect -13650 2579 -13616 2613
rect -13650 2511 -13616 2545
rect -13650 2443 -13616 2477
rect -13650 2375 -13616 2409
rect -13650 2307 -13616 2341
rect -13650 2239 -13616 2273
rect -13650 2171 -13616 2205
rect -13650 2103 -13616 2137
rect -13650 2035 -13616 2069
rect -13650 1967 -13616 2001
rect -13650 1899 -13616 1933
rect -13554 2783 -13520 2817
rect -13554 2715 -13520 2749
rect -13554 2647 -13520 2681
rect -13554 2579 -13520 2613
rect -13554 2511 -13520 2545
rect -13554 2443 -13520 2477
rect -13554 2375 -13520 2409
rect -13554 2307 -13520 2341
rect -13554 2239 -13520 2273
rect -13554 2171 -13520 2205
rect -13554 2103 -13520 2137
rect -13554 2035 -13520 2069
rect -13554 1967 -13520 2001
rect -13554 1899 -13520 1933
rect -13458 2783 -13424 2817
rect -13458 2715 -13424 2749
rect -13458 2647 -13424 2681
rect -13458 2579 -13424 2613
rect -13458 2511 -13424 2545
rect -13458 2443 -13424 2477
rect -13458 2375 -13424 2409
rect -13458 2307 -13424 2341
rect -13458 2239 -13424 2273
rect -13458 2171 -13424 2205
rect -13458 2103 -13424 2137
rect -13458 2035 -13424 2069
rect -13458 1967 -13424 2001
rect -13458 1899 -13424 1933
rect -13362 2783 -13328 2817
rect -13362 2715 -13328 2749
rect -13362 2647 -13328 2681
rect -13362 2579 -13328 2613
rect -13362 2511 -13328 2545
rect -13362 2443 -13328 2477
rect -13362 2375 -13328 2409
rect -13362 2307 -13328 2341
rect -13362 2239 -13328 2273
rect -13362 2171 -13328 2205
rect -13362 2103 -13328 2137
rect -13362 2035 -13328 2069
rect -13362 1967 -13328 2001
rect -13362 1899 -13328 1933
rect -13266 2783 -13232 2817
rect -13266 2715 -13232 2749
rect -13266 2647 -13232 2681
rect -13266 2579 -13232 2613
rect -13266 2511 -13232 2545
rect -13266 2443 -13232 2477
rect -13266 2375 -13232 2409
rect -13266 2307 -13232 2341
rect -13266 2239 -13232 2273
rect -13266 2171 -13232 2205
rect -13266 2103 -13232 2137
rect -13266 2035 -13232 2069
rect -13266 1967 -13232 2001
rect -13266 1899 -13232 1933
rect -13170 2783 -13136 2817
rect -13170 2715 -13136 2749
rect -13170 2647 -13136 2681
rect -13170 2579 -13136 2613
rect -13170 2511 -13136 2545
rect -13170 2443 -13136 2477
rect -13170 2375 -13136 2409
rect -13170 2307 -13136 2341
rect -13170 2239 -13136 2273
rect -13170 2171 -13136 2205
rect -13170 2103 -13136 2137
rect -13170 2035 -13136 2069
rect -13170 1967 -13136 2001
rect -13170 1899 -13136 1933
rect -13074 2783 -13040 2817
rect -13074 2715 -13040 2749
rect -13074 2647 -13040 2681
rect -13074 2579 -13040 2613
rect -13074 2511 -13040 2545
rect -13074 2443 -13040 2477
rect -13074 2375 -13040 2409
rect -13074 2307 -13040 2341
rect -13074 2239 -13040 2273
rect -13074 2171 -13040 2205
rect -13074 2103 -13040 2137
rect -13074 2035 -13040 2069
rect -13074 1967 -13040 2001
rect -13074 1899 -13040 1933
rect -12836 2787 -12802 2821
rect -12836 2719 -12802 2753
rect -12836 2651 -12802 2685
rect -12836 2583 -12802 2617
rect -12836 2515 -12802 2549
rect -12836 2447 -12802 2481
rect -12836 2379 -12802 2413
rect -12836 2311 -12802 2345
rect -12836 2243 -12802 2277
rect -12836 2175 -12802 2209
rect -12836 2107 -12802 2141
rect -12836 2039 -12802 2073
rect -12836 1971 -12802 2005
rect -12836 1903 -12802 1937
rect -12740 2787 -12706 2821
rect -12740 2719 -12706 2753
rect -12740 2651 -12706 2685
rect -12740 2583 -12706 2617
rect -12740 2515 -12706 2549
rect -12740 2447 -12706 2481
rect -12740 2379 -12706 2413
rect -12740 2311 -12706 2345
rect -12740 2243 -12706 2277
rect -12740 2175 -12706 2209
rect -12740 2107 -12706 2141
rect -12740 2039 -12706 2073
rect -12740 1971 -12706 2005
rect -12740 1903 -12706 1937
rect -12644 2787 -12610 2821
rect -12644 2719 -12610 2753
rect -12644 2651 -12610 2685
rect -12644 2583 -12610 2617
rect -12644 2515 -12610 2549
rect -12644 2447 -12610 2481
rect -12644 2379 -12610 2413
rect -12644 2311 -12610 2345
rect -12644 2243 -12610 2277
rect -12644 2175 -12610 2209
rect -12644 2107 -12610 2141
rect -12644 2039 -12610 2073
rect -12644 1971 -12610 2005
rect -12644 1903 -12610 1937
rect -12548 2787 -12514 2821
rect -12548 2719 -12514 2753
rect -12548 2651 -12514 2685
rect -12548 2583 -12514 2617
rect -12548 2515 -12514 2549
rect -12548 2447 -12514 2481
rect -12548 2379 -12514 2413
rect -12548 2311 -12514 2345
rect -12548 2243 -12514 2277
rect -12548 2175 -12514 2209
rect -12548 2107 -12514 2141
rect -12548 2039 -12514 2073
rect -12548 1971 -12514 2005
rect -12548 1903 -12514 1937
rect -12452 2787 -12418 2821
rect -12452 2719 -12418 2753
rect -12452 2651 -12418 2685
rect -12452 2583 -12418 2617
rect -12452 2515 -12418 2549
rect -12452 2447 -12418 2481
rect -12452 2379 -12418 2413
rect -12452 2311 -12418 2345
rect -12452 2243 -12418 2277
rect -12452 2175 -12418 2209
rect -12452 2107 -12418 2141
rect -12452 2039 -12418 2073
rect -12452 1971 -12418 2005
rect -12452 1903 -12418 1937
rect -12356 2787 -12322 2821
rect -12356 2719 -12322 2753
rect -12356 2651 -12322 2685
rect -12356 2583 -12322 2617
rect -12356 2515 -12322 2549
rect -12356 2447 -12322 2481
rect -12356 2379 -12322 2413
rect -12356 2311 -12322 2345
rect -12356 2243 -12322 2277
rect -12356 2175 -12322 2209
rect -12356 2107 -12322 2141
rect -12356 2039 -12322 2073
rect -12356 1971 -12322 2005
rect -12356 1903 -12322 1937
rect -12260 2787 -12226 2821
rect -12260 2719 -12226 2753
rect -12260 2651 -12226 2685
rect -12260 2583 -12226 2617
rect -12260 2515 -12226 2549
rect -12260 2447 -12226 2481
rect -12260 2379 -12226 2413
rect -12260 2311 -12226 2345
rect -12260 2243 -12226 2277
rect -12260 2175 -12226 2209
rect -12260 2107 -12226 2141
rect -12260 2039 -12226 2073
rect -12260 1971 -12226 2005
rect -12260 1903 -12226 1937
rect -12164 2787 -12130 2821
rect -12164 2719 -12130 2753
rect -12164 2651 -12130 2685
rect -12164 2583 -12130 2617
rect -12164 2515 -12130 2549
rect -12164 2447 -12130 2481
rect -12164 2379 -12130 2413
rect -12164 2311 -12130 2345
rect -12164 2243 -12130 2277
rect -12164 2175 -12130 2209
rect -12164 2107 -12130 2141
rect -12164 2039 -12130 2073
rect -12164 1971 -12130 2005
rect -12164 1903 -12130 1937
rect -12068 2787 -12034 2821
rect -12068 2719 -12034 2753
rect -12068 2651 -12034 2685
rect -12068 2583 -12034 2617
rect -12068 2515 -12034 2549
rect -12068 2447 -12034 2481
rect -12068 2379 -12034 2413
rect -12068 2311 -12034 2345
rect -12068 2243 -12034 2277
rect -12068 2175 -12034 2209
rect -12068 2107 -12034 2141
rect -12068 2039 -12034 2073
rect -12068 1971 -12034 2005
rect -12068 1903 -12034 1937
rect -11972 2787 -11938 2821
rect -11972 2719 -11938 2753
rect -11972 2651 -11938 2685
rect -11972 2583 -11938 2617
rect -11972 2515 -11938 2549
rect -11972 2447 -11938 2481
rect -11972 2379 -11938 2413
rect -11972 2311 -11938 2345
rect -11972 2243 -11938 2277
rect -11972 2175 -11938 2209
rect -11972 2107 -11938 2141
rect -11972 2039 -11938 2073
rect -11972 1971 -11938 2005
rect -11972 1903 -11938 1937
rect -11876 2787 -11842 2821
rect -11876 2719 -11842 2753
rect -11876 2651 -11842 2685
rect -11876 2583 -11842 2617
rect -11876 2515 -11842 2549
rect -11876 2447 -11842 2481
rect -11876 2379 -11842 2413
rect -11876 2311 -11842 2345
rect -11876 2243 -11842 2277
rect -11876 2175 -11842 2209
rect -11876 2107 -11842 2141
rect -11876 2039 -11842 2073
rect -11876 1971 -11842 2005
rect -11876 1903 -11842 1937
rect -11664 2797 -11630 2831
rect -11664 2729 -11630 2763
rect -11664 2661 -11630 2695
rect -11664 2593 -11630 2627
rect -11664 2525 -11630 2559
rect -11664 2457 -11630 2491
rect -11664 2389 -11630 2423
rect -11664 2321 -11630 2355
rect -11664 2253 -11630 2287
rect -11664 2185 -11630 2219
rect -11664 2117 -11630 2151
rect -11664 2049 -11630 2083
rect -11664 1981 -11630 2015
rect -11664 1913 -11630 1947
rect -11568 2797 -11534 2831
rect -11568 2729 -11534 2763
rect -11568 2661 -11534 2695
rect -11568 2593 -11534 2627
rect -11568 2525 -11534 2559
rect -11568 2457 -11534 2491
rect -11568 2389 -11534 2423
rect -11568 2321 -11534 2355
rect -11568 2253 -11534 2287
rect -11568 2185 -11534 2219
rect -11568 2117 -11534 2151
rect -11568 2049 -11534 2083
rect -11568 1981 -11534 2015
rect -11568 1913 -11534 1947
rect -11472 2797 -11438 2831
rect -11472 2729 -11438 2763
rect -11472 2661 -11438 2695
rect -11472 2593 -11438 2627
rect -11472 2525 -11438 2559
rect -11472 2457 -11438 2491
rect -11472 2389 -11438 2423
rect -11472 2321 -11438 2355
rect -11472 2253 -11438 2287
rect -11472 2185 -11438 2219
rect -11472 2117 -11438 2151
rect -11472 2049 -11438 2083
rect -11472 1981 -11438 2015
rect -11472 1913 -11438 1947
rect -11376 2797 -11342 2831
rect -11376 2729 -11342 2763
rect -11376 2661 -11342 2695
rect -11376 2593 -11342 2627
rect -11376 2525 -11342 2559
rect -11376 2457 -11342 2491
rect -11376 2389 -11342 2423
rect -11376 2321 -11342 2355
rect -11376 2253 -11342 2287
rect -11376 2185 -11342 2219
rect -11376 2117 -11342 2151
rect -11376 2049 -11342 2083
rect -11376 1981 -11342 2015
rect -11376 1913 -11342 1947
rect -11280 2797 -11246 2831
rect -11280 2729 -11246 2763
rect -11280 2661 -11246 2695
rect -11280 2593 -11246 2627
rect -11280 2525 -11246 2559
rect -11280 2457 -11246 2491
rect -11280 2389 -11246 2423
rect -11280 2321 -11246 2355
rect -11280 2253 -11246 2287
rect -11280 2185 -11246 2219
rect -11280 2117 -11246 2151
rect -11280 2049 -11246 2083
rect -11280 1981 -11246 2015
rect -11280 1913 -11246 1947
rect -11184 2797 -11150 2831
rect -11184 2729 -11150 2763
rect -11184 2661 -11150 2695
rect -11184 2593 -11150 2627
rect -11184 2525 -11150 2559
rect -11184 2457 -11150 2491
rect -11184 2389 -11150 2423
rect -11184 2321 -11150 2355
rect -11184 2253 -11150 2287
rect -11184 2185 -11150 2219
rect -11184 2117 -11150 2151
rect -11184 2049 -11150 2083
rect -11184 1981 -11150 2015
rect -11184 1913 -11150 1947
rect -10196 2789 -10162 2823
rect -10196 2721 -10162 2755
rect -10196 2653 -10162 2687
rect -10196 2585 -10162 2619
rect -10196 2517 -10162 2551
rect -10196 2449 -10162 2483
rect -10196 2381 -10162 2415
rect -10196 2313 -10162 2347
rect -10196 2245 -10162 2279
rect -10196 2177 -10162 2211
rect -10196 2109 -10162 2143
rect -10196 2041 -10162 2075
rect -10196 1973 -10162 2007
rect -10196 1905 -10162 1939
rect -10100 2789 -10066 2823
rect -10100 2721 -10066 2755
rect -10100 2653 -10066 2687
rect -10100 2585 -10066 2619
rect -10100 2517 -10066 2551
rect -10100 2449 -10066 2483
rect -10100 2381 -10066 2415
rect -10100 2313 -10066 2347
rect -10100 2245 -10066 2279
rect -10100 2177 -10066 2211
rect -10100 2109 -10066 2143
rect -10100 2041 -10066 2075
rect -10100 1973 -10066 2007
rect -10100 1905 -10066 1939
rect -10004 2789 -9970 2823
rect -10004 2721 -9970 2755
rect -10004 2653 -9970 2687
rect -10004 2585 -9970 2619
rect -10004 2517 -9970 2551
rect -10004 2449 -9970 2483
rect -10004 2381 -9970 2415
rect -10004 2313 -9970 2347
rect -10004 2245 -9970 2279
rect -10004 2177 -9970 2211
rect -10004 2109 -9970 2143
rect -10004 2041 -9970 2075
rect -10004 1973 -9970 2007
rect -10004 1905 -9970 1939
rect -9908 2789 -9874 2823
rect -9908 2721 -9874 2755
rect -9908 2653 -9874 2687
rect -9908 2585 -9874 2619
rect -9908 2517 -9874 2551
rect -9908 2449 -9874 2483
rect -9908 2381 -9874 2415
rect -9908 2313 -9874 2347
rect -9908 2245 -9874 2279
rect -9908 2177 -9874 2211
rect -9908 2109 -9874 2143
rect -9908 2041 -9874 2075
rect -9908 1973 -9874 2007
rect -9908 1905 -9874 1939
rect -9812 2789 -9778 2823
rect -9812 2721 -9778 2755
rect -9812 2653 -9778 2687
rect -9812 2585 -9778 2619
rect -9812 2517 -9778 2551
rect -9812 2449 -9778 2483
rect -9812 2381 -9778 2415
rect -9812 2313 -9778 2347
rect -9812 2245 -9778 2279
rect -9812 2177 -9778 2211
rect -9812 2109 -9778 2143
rect -9812 2041 -9778 2075
rect -9812 1973 -9778 2007
rect -9812 1905 -9778 1939
rect -9716 2789 -9682 2823
rect -9716 2721 -9682 2755
rect -9716 2653 -9682 2687
rect -9716 2585 -9682 2619
rect -9716 2517 -9682 2551
rect -9716 2449 -9682 2483
rect -9716 2381 -9682 2415
rect -9716 2313 -9682 2347
rect -9716 2245 -9682 2279
rect -9716 2177 -9682 2211
rect -9716 2109 -9682 2143
rect -9716 2041 -9682 2075
rect -9716 1973 -9682 2007
rect -9716 1905 -9682 1939
rect -9620 2789 -9586 2823
rect -9620 2721 -9586 2755
rect -9620 2653 -9586 2687
rect -9620 2585 -9586 2619
rect -9620 2517 -9586 2551
rect -9620 2449 -9586 2483
rect -9620 2381 -9586 2415
rect -9620 2313 -9586 2347
rect -9620 2245 -9586 2279
rect -9620 2177 -9586 2211
rect -9620 2109 -9586 2143
rect -9620 2041 -9586 2075
rect -9620 1973 -9586 2007
rect -9620 1905 -9586 1939
rect -9524 2789 -9490 2823
rect -9524 2721 -9490 2755
rect -9524 2653 -9490 2687
rect -9524 2585 -9490 2619
rect -9524 2517 -9490 2551
rect -9524 2449 -9490 2483
rect -9524 2381 -9490 2415
rect -9524 2313 -9490 2347
rect -9524 2245 -9490 2279
rect -9524 2177 -9490 2211
rect -9524 2109 -9490 2143
rect -9524 2041 -9490 2075
rect -9524 1973 -9490 2007
rect -9524 1905 -9490 1939
rect -9428 2789 -9394 2823
rect -9428 2721 -9394 2755
rect -9428 2653 -9394 2687
rect -9428 2585 -9394 2619
rect -9428 2517 -9394 2551
rect -9428 2449 -9394 2483
rect -9428 2381 -9394 2415
rect -9428 2313 -9394 2347
rect -9428 2245 -9394 2279
rect -9428 2177 -9394 2211
rect -9428 2109 -9394 2143
rect -9428 2041 -9394 2075
rect -9428 1973 -9394 2007
rect -9428 1905 -9394 1939
rect -9332 2789 -9298 2823
rect -9332 2721 -9298 2755
rect -9332 2653 -9298 2687
rect -9332 2585 -9298 2619
rect -9332 2517 -9298 2551
rect -9332 2449 -9298 2483
rect -9332 2381 -9298 2415
rect -9332 2313 -9298 2347
rect -9332 2245 -9298 2279
rect -9332 2177 -9298 2211
rect -9332 2109 -9298 2143
rect -9332 2041 -9298 2075
rect -9332 1973 -9298 2007
rect -9332 1905 -9298 1939
rect -9236 2789 -9202 2823
rect -9236 2721 -9202 2755
rect -9236 2653 -9202 2687
rect -9236 2585 -9202 2619
rect -9236 2517 -9202 2551
rect -9236 2449 -9202 2483
rect -9236 2381 -9202 2415
rect -9236 2313 -9202 2347
rect -9236 2245 -9202 2279
rect -9236 2177 -9202 2211
rect -9236 2109 -9202 2143
rect -9236 2041 -9202 2075
rect -9236 1973 -9202 2007
rect -9236 1905 -9202 1939
rect -9140 2789 -9106 2823
rect -9140 2721 -9106 2755
rect -9140 2653 -9106 2687
rect -9140 2585 -9106 2619
rect -9140 2517 -9106 2551
rect -9140 2449 -9106 2483
rect -9140 2381 -9106 2415
rect -9140 2313 -9106 2347
rect -9140 2245 -9106 2279
rect -9140 2177 -9106 2211
rect -9140 2109 -9106 2143
rect -9140 2041 -9106 2075
rect -9140 1973 -9106 2007
rect -9140 1905 -9106 1939
rect -9044 2789 -9010 2823
rect -9044 2721 -9010 2755
rect -9044 2653 -9010 2687
rect -9044 2585 -9010 2619
rect -9044 2517 -9010 2551
rect -9044 2449 -9010 2483
rect -9044 2381 -9010 2415
rect -9044 2313 -9010 2347
rect -9044 2245 -9010 2279
rect -9044 2177 -9010 2211
rect -9044 2109 -9010 2143
rect -9044 2041 -9010 2075
rect -9044 1973 -9010 2007
rect -9044 1905 -9010 1939
rect -8948 2789 -8914 2823
rect -8948 2721 -8914 2755
rect -8948 2653 -8914 2687
rect -8948 2585 -8914 2619
rect -8948 2517 -8914 2551
rect -8948 2449 -8914 2483
rect -8948 2381 -8914 2415
rect -8948 2313 -8914 2347
rect -8948 2245 -8914 2279
rect -8948 2177 -8914 2211
rect -8948 2109 -8914 2143
rect -8948 2041 -8914 2075
rect -8948 1973 -8914 2007
rect -8948 1905 -8914 1939
rect -8852 2789 -8818 2823
rect -8852 2721 -8818 2755
rect -8852 2653 -8818 2687
rect -8852 2585 -8818 2619
rect -8852 2517 -8818 2551
rect -8852 2449 -8818 2483
rect -8852 2381 -8818 2415
rect -8852 2313 -8818 2347
rect -8852 2245 -8818 2279
rect -8852 2177 -8818 2211
rect -8852 2109 -8818 2143
rect -8852 2041 -8818 2075
rect -8852 1973 -8818 2007
rect -8852 1905 -8818 1939
rect -8756 2789 -8722 2823
rect -8756 2721 -8722 2755
rect -8756 2653 -8722 2687
rect -8756 2585 -8722 2619
rect -8756 2517 -8722 2551
rect -8756 2449 -8722 2483
rect -8756 2381 -8722 2415
rect -8756 2313 -8722 2347
rect -8756 2245 -8722 2279
rect -8756 2177 -8722 2211
rect -8756 2109 -8722 2143
rect -8756 2041 -8722 2075
rect -8756 1973 -8722 2007
rect -8756 1905 -8722 1939
rect -8660 2789 -8626 2823
rect -8660 2721 -8626 2755
rect -8660 2653 -8626 2687
rect -8660 2585 -8626 2619
rect -8660 2517 -8626 2551
rect -8660 2449 -8626 2483
rect -8660 2381 -8626 2415
rect -8660 2313 -8626 2347
rect -8660 2245 -8626 2279
rect -8660 2177 -8626 2211
rect -8660 2109 -8626 2143
rect -8660 2041 -8626 2075
rect -8660 1973 -8626 2007
rect -8660 1905 -8626 1939
rect -8564 2789 -8530 2823
rect -8564 2721 -8530 2755
rect -8564 2653 -8530 2687
rect -8564 2585 -8530 2619
rect -8564 2517 -8530 2551
rect -8564 2449 -8530 2483
rect -8564 2381 -8530 2415
rect -8564 2313 -8530 2347
rect -8564 2245 -8530 2279
rect -8564 2177 -8530 2211
rect -8564 2109 -8530 2143
rect -8564 2041 -8530 2075
rect -8564 1973 -8530 2007
rect -8564 1905 -8530 1939
rect -8468 2789 -8434 2823
rect -8468 2721 -8434 2755
rect -8468 2653 -8434 2687
rect -8468 2585 -8434 2619
rect -8468 2517 -8434 2551
rect -8468 2449 -8434 2483
rect -8468 2381 -8434 2415
rect -8468 2313 -8434 2347
rect -8468 2245 -8434 2279
rect -8468 2177 -8434 2211
rect -8468 2109 -8434 2143
rect -8468 2041 -8434 2075
rect -8468 1973 -8434 2007
rect -8468 1905 -8434 1939
rect -8372 2789 -8338 2823
rect -8372 2721 -8338 2755
rect -8372 2653 -8338 2687
rect -8372 2585 -8338 2619
rect -8372 2517 -8338 2551
rect -8372 2449 -8338 2483
rect -8372 2381 -8338 2415
rect -8372 2313 -8338 2347
rect -8372 2245 -8338 2279
rect -8372 2177 -8338 2211
rect -8372 2109 -8338 2143
rect -8372 2041 -8338 2075
rect -8372 1973 -8338 2007
rect -8372 1905 -8338 1939
rect -1686 2889 -1652 2923
rect -8276 2789 -8242 2823
rect -8276 2721 -8242 2755
rect -8276 2653 -8242 2687
rect -8276 2585 -8242 2619
rect -8276 2517 -8242 2551
rect -8276 2449 -8242 2483
rect -8276 2381 -8242 2415
rect -8276 2313 -8242 2347
rect -8276 2245 -8242 2279
rect -8276 2177 -8242 2211
rect -8276 2109 -8242 2143
rect -8276 2041 -8242 2075
rect -8276 1973 -8242 2007
rect -8276 1905 -8242 1939
rect -8048 2781 -8014 2815
rect -8048 2713 -8014 2747
rect -8048 2645 -8014 2679
rect -8048 2577 -8014 2611
rect -8048 2509 -8014 2543
rect -8048 2441 -8014 2475
rect -8048 2373 -8014 2407
rect -8048 2305 -8014 2339
rect -8048 2237 -8014 2271
rect -8048 2169 -8014 2203
rect -8048 2101 -8014 2135
rect -8048 2033 -8014 2067
rect -8048 1965 -8014 1999
rect -8048 1897 -8014 1931
rect -7952 2781 -7918 2815
rect -7952 2713 -7918 2747
rect -7952 2645 -7918 2679
rect -7952 2577 -7918 2611
rect -7952 2509 -7918 2543
rect -7952 2441 -7918 2475
rect -7952 2373 -7918 2407
rect -7952 2305 -7918 2339
rect -7952 2237 -7918 2271
rect -7952 2169 -7918 2203
rect -7952 2101 -7918 2135
rect -7952 2033 -7918 2067
rect -7952 1965 -7918 1999
rect -7952 1897 -7918 1931
rect -7856 2781 -7822 2815
rect -7856 2713 -7822 2747
rect -7856 2645 -7822 2679
rect -7856 2577 -7822 2611
rect -7856 2509 -7822 2543
rect -7856 2441 -7822 2475
rect -7856 2373 -7822 2407
rect -7856 2305 -7822 2339
rect -7856 2237 -7822 2271
rect -7856 2169 -7822 2203
rect -7856 2101 -7822 2135
rect -7856 2033 -7822 2067
rect -7856 1965 -7822 1999
rect -7856 1897 -7822 1931
rect -7760 2781 -7726 2815
rect -7760 2713 -7726 2747
rect -7760 2645 -7726 2679
rect -7760 2577 -7726 2611
rect -7760 2509 -7726 2543
rect -7760 2441 -7726 2475
rect -7760 2373 -7726 2407
rect -7760 2305 -7726 2339
rect -7760 2237 -7726 2271
rect -7760 2169 -7726 2203
rect -7760 2101 -7726 2135
rect -7760 2033 -7726 2067
rect -7760 1965 -7726 1999
rect -7760 1897 -7726 1931
rect -7664 2781 -7630 2815
rect -7664 2713 -7630 2747
rect -7664 2645 -7630 2679
rect -7664 2577 -7630 2611
rect -7664 2509 -7630 2543
rect -7664 2441 -7630 2475
rect -7664 2373 -7630 2407
rect -7664 2305 -7630 2339
rect -7664 2237 -7630 2271
rect -7664 2169 -7630 2203
rect -7664 2101 -7630 2135
rect -7664 2033 -7630 2067
rect -7664 1965 -7630 1999
rect -7664 1897 -7630 1931
rect -7568 2781 -7534 2815
rect -7568 2713 -7534 2747
rect -7568 2645 -7534 2679
rect -7568 2577 -7534 2611
rect -7568 2509 -7534 2543
rect -7568 2441 -7534 2475
rect -7568 2373 -7534 2407
rect -7568 2305 -7534 2339
rect -7568 2237 -7534 2271
rect -7568 2169 -7534 2203
rect -7568 2101 -7534 2135
rect -7568 2033 -7534 2067
rect -7568 1965 -7534 1999
rect -7568 1897 -7534 1931
rect -7472 2781 -7438 2815
rect -7472 2713 -7438 2747
rect -7472 2645 -7438 2679
rect -7472 2577 -7438 2611
rect -7472 2509 -7438 2543
rect -7472 2441 -7438 2475
rect -7472 2373 -7438 2407
rect -7472 2305 -7438 2339
rect -7472 2237 -7438 2271
rect -7472 2169 -7438 2203
rect -7472 2101 -7438 2135
rect -7472 2033 -7438 2067
rect -7472 1965 -7438 1999
rect -7472 1897 -7438 1931
rect -7376 2781 -7342 2815
rect -7376 2713 -7342 2747
rect -7376 2645 -7342 2679
rect -7376 2577 -7342 2611
rect -7376 2509 -7342 2543
rect -7376 2441 -7342 2475
rect -7376 2373 -7342 2407
rect -7376 2305 -7342 2339
rect -7376 2237 -7342 2271
rect -7376 2169 -7342 2203
rect -7376 2101 -7342 2135
rect -7376 2033 -7342 2067
rect -7376 1965 -7342 1999
rect -7376 1897 -7342 1931
rect -7280 2781 -7246 2815
rect -7280 2713 -7246 2747
rect -7280 2645 -7246 2679
rect -7280 2577 -7246 2611
rect -7280 2509 -7246 2543
rect -7280 2441 -7246 2475
rect -7280 2373 -7246 2407
rect -7280 2305 -7246 2339
rect -7280 2237 -7246 2271
rect -7280 2169 -7246 2203
rect -7280 2101 -7246 2135
rect -7280 2033 -7246 2067
rect -7280 1965 -7246 1999
rect -7280 1897 -7246 1931
rect -7184 2781 -7150 2815
rect -7184 2713 -7150 2747
rect -7184 2645 -7150 2679
rect -7184 2577 -7150 2611
rect -7184 2509 -7150 2543
rect -7184 2441 -7150 2475
rect -7184 2373 -7150 2407
rect -7184 2305 -7150 2339
rect -7184 2237 -7150 2271
rect -7184 2169 -7150 2203
rect -7184 2101 -7150 2135
rect -7184 2033 -7150 2067
rect -7184 1965 -7150 1999
rect -7184 1897 -7150 1931
rect -7088 2781 -7054 2815
rect -7088 2713 -7054 2747
rect -7088 2645 -7054 2679
rect -7088 2577 -7054 2611
rect -7088 2509 -7054 2543
rect -7088 2441 -7054 2475
rect -7088 2373 -7054 2407
rect -7088 2305 -7054 2339
rect -7088 2237 -7054 2271
rect -7088 2169 -7054 2203
rect -7088 2101 -7054 2135
rect -7088 2033 -7054 2067
rect -7088 1965 -7054 1999
rect -7088 1897 -7054 1931
rect -6992 2781 -6958 2815
rect -6992 2713 -6958 2747
rect -6992 2645 -6958 2679
rect -6992 2577 -6958 2611
rect -6992 2509 -6958 2543
rect -6992 2441 -6958 2475
rect -6992 2373 -6958 2407
rect -6992 2305 -6958 2339
rect -6992 2237 -6958 2271
rect -6992 2169 -6958 2203
rect -6992 2101 -6958 2135
rect -6992 2033 -6958 2067
rect -6992 1965 -6958 1999
rect -6992 1897 -6958 1931
rect -6896 2781 -6862 2815
rect -6896 2713 -6862 2747
rect -6896 2645 -6862 2679
rect -6896 2577 -6862 2611
rect -6896 2509 -6862 2543
rect -6896 2441 -6862 2475
rect -6896 2373 -6862 2407
rect -6896 2305 -6862 2339
rect -6896 2237 -6862 2271
rect -6896 2169 -6862 2203
rect -6896 2101 -6862 2135
rect -6896 2033 -6862 2067
rect -6896 1965 -6862 1999
rect -6896 1897 -6862 1931
rect -6800 2781 -6766 2815
rect -6800 2713 -6766 2747
rect -6800 2645 -6766 2679
rect -6800 2577 -6766 2611
rect -6800 2509 -6766 2543
rect -6800 2441 -6766 2475
rect -6800 2373 -6766 2407
rect -6800 2305 -6766 2339
rect -6800 2237 -6766 2271
rect -6800 2169 -6766 2203
rect -6800 2101 -6766 2135
rect -6800 2033 -6766 2067
rect -6800 1965 -6766 1999
rect -6800 1897 -6766 1931
rect -6704 2781 -6670 2815
rect -6704 2713 -6670 2747
rect -6704 2645 -6670 2679
rect -6704 2577 -6670 2611
rect -6704 2509 -6670 2543
rect -6704 2441 -6670 2475
rect -6704 2373 -6670 2407
rect -6704 2305 -6670 2339
rect -6704 2237 -6670 2271
rect -6704 2169 -6670 2203
rect -6704 2101 -6670 2135
rect -6704 2033 -6670 2067
rect -6704 1965 -6670 1999
rect -6704 1897 -6670 1931
rect -6608 2781 -6574 2815
rect -6608 2713 -6574 2747
rect -6608 2645 -6574 2679
rect -6608 2577 -6574 2611
rect -6608 2509 -6574 2543
rect -6608 2441 -6574 2475
rect -6608 2373 -6574 2407
rect -6608 2305 -6574 2339
rect -6608 2237 -6574 2271
rect -6608 2169 -6574 2203
rect -6608 2101 -6574 2135
rect -6608 2033 -6574 2067
rect -6608 1965 -6574 1999
rect -6608 1897 -6574 1931
rect -6370 2785 -6336 2819
rect -6370 2717 -6336 2751
rect -6370 2649 -6336 2683
rect -6370 2581 -6336 2615
rect -6370 2513 -6336 2547
rect -6370 2445 -6336 2479
rect -6370 2377 -6336 2411
rect -6370 2309 -6336 2343
rect -6370 2241 -6336 2275
rect -6370 2173 -6336 2207
rect -6370 2105 -6336 2139
rect -6370 2037 -6336 2071
rect -6370 1969 -6336 2003
rect -6370 1901 -6336 1935
rect -6274 2785 -6240 2819
rect -6274 2717 -6240 2751
rect -6274 2649 -6240 2683
rect -6274 2581 -6240 2615
rect -6274 2513 -6240 2547
rect -6274 2445 -6240 2479
rect -6274 2377 -6240 2411
rect -6274 2309 -6240 2343
rect -6274 2241 -6240 2275
rect -6274 2173 -6240 2207
rect -6274 2105 -6240 2139
rect -6274 2037 -6240 2071
rect -6274 1969 -6240 2003
rect -6274 1901 -6240 1935
rect -6178 2785 -6144 2819
rect -6178 2717 -6144 2751
rect -6178 2649 -6144 2683
rect -6178 2581 -6144 2615
rect -6178 2513 -6144 2547
rect -6178 2445 -6144 2479
rect -6178 2377 -6144 2411
rect -6178 2309 -6144 2343
rect -6178 2241 -6144 2275
rect -6178 2173 -6144 2207
rect -6178 2105 -6144 2139
rect -6178 2037 -6144 2071
rect -6178 1969 -6144 2003
rect -6178 1901 -6144 1935
rect -6082 2785 -6048 2819
rect -6082 2717 -6048 2751
rect -6082 2649 -6048 2683
rect -6082 2581 -6048 2615
rect -6082 2513 -6048 2547
rect -6082 2445 -6048 2479
rect -6082 2377 -6048 2411
rect -6082 2309 -6048 2343
rect -6082 2241 -6048 2275
rect -6082 2173 -6048 2207
rect -6082 2105 -6048 2139
rect -6082 2037 -6048 2071
rect -6082 1969 -6048 2003
rect -6082 1901 -6048 1935
rect -5986 2785 -5952 2819
rect -5986 2717 -5952 2751
rect -5986 2649 -5952 2683
rect -5986 2581 -5952 2615
rect -5986 2513 -5952 2547
rect -5986 2445 -5952 2479
rect -5986 2377 -5952 2411
rect -5986 2309 -5952 2343
rect -5986 2241 -5952 2275
rect -5986 2173 -5952 2207
rect -5986 2105 -5952 2139
rect -5986 2037 -5952 2071
rect -5986 1969 -5952 2003
rect -5986 1901 -5952 1935
rect -5890 2785 -5856 2819
rect -5890 2717 -5856 2751
rect -5890 2649 -5856 2683
rect -5890 2581 -5856 2615
rect -5890 2513 -5856 2547
rect -5890 2445 -5856 2479
rect -5890 2377 -5856 2411
rect -5890 2309 -5856 2343
rect -5890 2241 -5856 2275
rect -5890 2173 -5856 2207
rect -5890 2105 -5856 2139
rect -5890 2037 -5856 2071
rect -5890 1969 -5856 2003
rect -5890 1901 -5856 1935
rect -5794 2785 -5760 2819
rect -5794 2717 -5760 2751
rect -5794 2649 -5760 2683
rect -5794 2581 -5760 2615
rect -5794 2513 -5760 2547
rect -5794 2445 -5760 2479
rect -5794 2377 -5760 2411
rect -5794 2309 -5760 2343
rect -5794 2241 -5760 2275
rect -5794 2173 -5760 2207
rect -5794 2105 -5760 2139
rect -5794 2037 -5760 2071
rect -5794 1969 -5760 2003
rect -5794 1901 -5760 1935
rect -5698 2785 -5664 2819
rect -5698 2717 -5664 2751
rect -5698 2649 -5664 2683
rect -5698 2581 -5664 2615
rect -5698 2513 -5664 2547
rect -5698 2445 -5664 2479
rect -5698 2377 -5664 2411
rect -5698 2309 -5664 2343
rect -5698 2241 -5664 2275
rect -5698 2173 -5664 2207
rect -5698 2105 -5664 2139
rect -5698 2037 -5664 2071
rect -5698 1969 -5664 2003
rect -5698 1901 -5664 1935
rect -5602 2785 -5568 2819
rect -5602 2717 -5568 2751
rect -5602 2649 -5568 2683
rect -5602 2581 -5568 2615
rect -5602 2513 -5568 2547
rect -5602 2445 -5568 2479
rect -5602 2377 -5568 2411
rect -5602 2309 -5568 2343
rect -5602 2241 -5568 2275
rect -5602 2173 -5568 2207
rect -5602 2105 -5568 2139
rect -5602 2037 -5568 2071
rect -5602 1969 -5568 2003
rect -5602 1901 -5568 1935
rect -5506 2785 -5472 2819
rect -5506 2717 -5472 2751
rect -5506 2649 -5472 2683
rect -5506 2581 -5472 2615
rect -5506 2513 -5472 2547
rect -5506 2445 -5472 2479
rect -5506 2377 -5472 2411
rect -5506 2309 -5472 2343
rect -5506 2241 -5472 2275
rect -5506 2173 -5472 2207
rect -5506 2105 -5472 2139
rect -5506 2037 -5472 2071
rect -5506 1969 -5472 2003
rect -5506 1901 -5472 1935
rect -5410 2785 -5376 2819
rect -5410 2717 -5376 2751
rect -5410 2649 -5376 2683
rect -5410 2581 -5376 2615
rect -5410 2513 -5376 2547
rect -5410 2445 -5376 2479
rect -5410 2377 -5376 2411
rect -5410 2309 -5376 2343
rect -5410 2241 -5376 2275
rect -5410 2173 -5376 2207
rect -5410 2105 -5376 2139
rect -5410 2037 -5376 2071
rect -5410 1969 -5376 2003
rect -5410 1901 -5376 1935
rect -5198 2795 -5164 2829
rect -5198 2727 -5164 2761
rect -5198 2659 -5164 2693
rect -5198 2591 -5164 2625
rect -5198 2523 -5164 2557
rect -5198 2455 -5164 2489
rect -5198 2387 -5164 2421
rect -5198 2319 -5164 2353
rect -5198 2251 -5164 2285
rect -5198 2183 -5164 2217
rect -5198 2115 -5164 2149
rect -5198 2047 -5164 2081
rect -5198 1979 -5164 2013
rect -5198 1911 -5164 1945
rect -5102 2795 -5068 2829
rect -5102 2727 -5068 2761
rect -5102 2659 -5068 2693
rect -5102 2591 -5068 2625
rect -5102 2523 -5068 2557
rect -5102 2455 -5068 2489
rect -5102 2387 -5068 2421
rect -5102 2319 -5068 2353
rect -5102 2251 -5068 2285
rect -5102 2183 -5068 2217
rect -5102 2115 -5068 2149
rect -5102 2047 -5068 2081
rect -5102 1979 -5068 2013
rect -5102 1911 -5068 1945
rect -5006 2795 -4972 2829
rect -5006 2727 -4972 2761
rect -5006 2659 -4972 2693
rect -5006 2591 -4972 2625
rect -5006 2523 -4972 2557
rect -5006 2455 -4972 2489
rect -5006 2387 -4972 2421
rect -5006 2319 -4972 2353
rect -5006 2251 -4972 2285
rect -5006 2183 -4972 2217
rect -5006 2115 -4972 2149
rect -5006 2047 -4972 2081
rect -5006 1979 -4972 2013
rect -5006 1911 -4972 1945
rect -4910 2795 -4876 2829
rect -4910 2727 -4876 2761
rect -4910 2659 -4876 2693
rect -4910 2591 -4876 2625
rect -4910 2523 -4876 2557
rect -4910 2455 -4876 2489
rect -4910 2387 -4876 2421
rect -4910 2319 -4876 2353
rect -4910 2251 -4876 2285
rect -4910 2183 -4876 2217
rect -4910 2115 -4876 2149
rect -4910 2047 -4876 2081
rect -4910 1979 -4876 2013
rect -4910 1911 -4876 1945
rect -4814 2795 -4780 2829
rect -4814 2727 -4780 2761
rect -4814 2659 -4780 2693
rect -4814 2591 -4780 2625
rect -4814 2523 -4780 2557
rect -4814 2455 -4780 2489
rect -4814 2387 -4780 2421
rect -4814 2319 -4780 2353
rect -4814 2251 -4780 2285
rect -4814 2183 -4780 2217
rect -4814 2115 -4780 2149
rect -4814 2047 -4780 2081
rect -4814 1979 -4780 2013
rect -4814 1911 -4780 1945
rect -4718 2795 -4684 2829
rect -4718 2727 -4684 2761
rect -4718 2659 -4684 2693
rect -4718 2591 -4684 2625
rect -4718 2523 -4684 2557
rect -4718 2455 -4684 2489
rect -4718 2387 -4684 2421
rect -4718 2319 -4684 2353
rect -4718 2251 -4684 2285
rect -1686 2821 -1652 2855
rect -1686 2753 -1652 2787
rect -1686 2685 -1652 2719
rect -1686 2617 -1652 2651
rect -1686 2549 -1652 2583
rect -1686 2481 -1652 2515
rect -1686 2413 -1652 2447
rect -1686 2345 -1652 2379
rect -1686 2277 -1652 2311
rect -1590 3161 -1556 3195
rect -1590 3093 -1556 3127
rect -1590 3025 -1556 3059
rect -1590 2957 -1556 2991
rect -1590 2889 -1556 2923
rect -1590 2821 -1556 2855
rect -1590 2753 -1556 2787
rect -1590 2685 -1556 2719
rect -1590 2617 -1556 2651
rect -1590 2549 -1556 2583
rect -1590 2481 -1556 2515
rect -1590 2413 -1556 2447
rect -1590 2345 -1556 2379
rect -1590 2277 -1556 2311
rect -1494 3161 -1460 3195
rect -1494 3093 -1460 3127
rect -1494 3025 -1460 3059
rect -1494 2957 -1460 2991
rect -1494 2889 -1460 2923
rect -1494 2821 -1460 2855
rect -1494 2753 -1460 2787
rect -1494 2685 -1460 2719
rect -1494 2617 -1460 2651
rect -1494 2549 -1460 2583
rect -1494 2481 -1460 2515
rect -1494 2413 -1460 2447
rect -1494 2345 -1460 2379
rect -1494 2277 -1460 2311
rect -1398 3161 -1364 3195
rect -1398 3093 -1364 3127
rect -1398 3025 -1364 3059
rect -1398 2957 -1364 2991
rect -1398 2889 -1364 2923
rect -1398 2821 -1364 2855
rect -1398 2753 -1364 2787
rect -1398 2685 -1364 2719
rect -1398 2617 -1364 2651
rect -1398 2549 -1364 2583
rect -1398 2481 -1364 2515
rect -1398 2413 -1364 2447
rect -1398 2345 -1364 2379
rect -1398 2277 -1364 2311
rect -1302 3161 -1268 3195
rect -1302 3093 -1268 3127
rect -1302 3025 -1268 3059
rect -1302 2957 -1268 2991
rect -1302 2889 -1268 2923
rect -1302 2821 -1268 2855
rect -1302 2753 -1268 2787
rect -1302 2685 -1268 2719
rect -1302 2617 -1268 2651
rect -1302 2549 -1268 2583
rect -1302 2481 -1268 2515
rect -1302 2413 -1268 2447
rect -1302 2345 -1268 2379
rect -1302 2277 -1268 2311
rect -1206 3161 -1172 3195
rect -1206 3093 -1172 3127
rect -1206 3025 -1172 3059
rect -1206 2957 -1172 2991
rect -1206 2889 -1172 2923
rect -1206 2821 -1172 2855
rect -1206 2753 -1172 2787
rect -1206 2685 -1172 2719
rect -1206 2617 -1172 2651
rect -1206 2549 -1172 2583
rect -1206 2481 -1172 2515
rect -1206 2413 -1172 2447
rect -1206 2345 -1172 2379
rect -1206 2277 -1172 2311
rect -1110 3161 -1076 3195
rect -1110 3093 -1076 3127
rect -1110 3025 -1076 3059
rect -1110 2957 -1076 2991
rect -1110 2889 -1076 2923
rect -1110 2821 -1076 2855
rect -1110 2753 -1076 2787
rect -1110 2685 -1076 2719
rect -1110 2617 -1076 2651
rect -1110 2549 -1076 2583
rect -1110 2481 -1076 2515
rect -1110 2413 -1076 2447
rect -1110 2345 -1076 2379
rect -1110 2277 -1076 2311
rect -1014 3161 -980 3195
rect -1014 3093 -980 3127
rect -1014 3025 -980 3059
rect -1014 2957 -980 2991
rect -1014 2889 -980 2923
rect -1014 2821 -980 2855
rect -1014 2753 -980 2787
rect -1014 2685 -980 2719
rect -1014 2617 -980 2651
rect -1014 2549 -980 2583
rect -1014 2481 -980 2515
rect -1014 2413 -980 2447
rect -1014 2345 -980 2379
rect -1014 2277 -980 2311
rect -918 3161 -884 3195
rect -918 3093 -884 3127
rect -918 3025 -884 3059
rect 16686 3187 16720 3221
rect 16686 3119 16720 3153
rect 16686 3051 16720 3085
rect -918 2957 -884 2991
rect -918 2889 -884 2923
rect 16686 2983 16720 3017
rect -918 2821 -884 2855
rect -918 2753 -884 2787
rect -918 2685 -884 2719
rect -918 2617 -884 2651
rect -918 2549 -884 2583
rect -918 2481 -884 2515
rect -918 2413 -884 2447
rect -918 2345 -884 2379
rect -918 2277 -884 2311
rect 1482 2755 1516 2789
rect 1482 2687 1516 2721
rect 1482 2619 1516 2653
rect 1482 2551 1516 2585
rect 1482 2483 1516 2517
rect 1482 2415 1516 2449
rect 1482 2347 1516 2381
rect 1482 2279 1516 2313
rect -4718 2183 -4684 2217
rect 1482 2211 1516 2245
rect -4718 2115 -4684 2149
rect -4718 2047 -4684 2081
rect -4718 1979 -4684 2013
rect -4718 1911 -4684 1945
rect 1482 2143 1516 2177
rect 1482 2075 1516 2109
rect 1482 2007 1516 2041
rect 1482 1939 1516 1973
rect 1482 1871 1516 1905
rect 1578 2755 1612 2789
rect 1578 2687 1612 2721
rect 1578 2619 1612 2653
rect 1578 2551 1612 2585
rect 1578 2483 1612 2517
rect 1578 2415 1612 2449
rect 1578 2347 1612 2381
rect 1578 2279 1612 2313
rect 1578 2211 1612 2245
rect 1578 2143 1612 2177
rect 1578 2075 1612 2109
rect 1578 2007 1612 2041
rect 1578 1939 1612 1973
rect 1578 1871 1612 1905
rect 1674 2755 1708 2789
rect 1674 2687 1708 2721
rect 1674 2619 1708 2653
rect 1674 2551 1708 2585
rect 1674 2483 1708 2517
rect 1674 2415 1708 2449
rect 1674 2347 1708 2381
rect 1674 2279 1708 2313
rect 1674 2211 1708 2245
rect 1674 2143 1708 2177
rect 1674 2075 1708 2109
rect 1674 2007 1708 2041
rect 1674 1939 1708 1973
rect 1674 1871 1708 1905
rect 1770 2755 1804 2789
rect 1770 2687 1804 2721
rect 1770 2619 1804 2653
rect 1770 2551 1804 2585
rect 1770 2483 1804 2517
rect 1770 2415 1804 2449
rect 1770 2347 1804 2381
rect 1770 2279 1804 2313
rect 1770 2211 1804 2245
rect 1770 2143 1804 2177
rect 1770 2075 1804 2109
rect 1770 2007 1804 2041
rect 1770 1939 1804 1973
rect 1770 1871 1804 1905
rect 16686 2915 16720 2949
rect 1866 2755 1900 2789
rect 1866 2687 1900 2721
rect 1866 2619 1900 2653
rect 1866 2551 1900 2585
rect 1866 2483 1900 2517
rect 1866 2415 1900 2449
rect 4438 2739 4472 2773
rect 4438 2671 4472 2705
rect 4438 2603 4472 2637
rect 4438 2535 4472 2569
rect 4438 2467 4472 2501
rect 1866 2347 1900 2381
rect 1866 2279 1900 2313
rect 4438 2399 4472 2433
rect 4438 2331 4472 2365
rect 1866 2211 1900 2245
rect 1866 2143 1900 2177
rect 1866 2075 1900 2109
rect 2500 2227 2534 2261
rect 2500 2159 2534 2193
rect 2500 2091 2534 2125
rect 2658 2227 2692 2261
rect 2658 2159 2692 2193
rect 2658 2091 2692 2125
rect 4438 2263 4472 2297
rect 4438 2195 4472 2229
rect 4438 2127 4472 2161
rect 4438 2059 4472 2093
rect 1866 2007 1900 2041
rect 1866 1939 1900 1973
rect 1866 1871 1900 1905
rect 4438 1991 4472 2025
rect 4438 1923 4472 1957
rect 4438 1855 4472 1889
rect 4534 2739 4568 2773
rect 4534 2671 4568 2705
rect 4534 2603 4568 2637
rect 4534 2535 4568 2569
rect 4534 2467 4568 2501
rect 4534 2399 4568 2433
rect 4534 2331 4568 2365
rect 4534 2263 4568 2297
rect 4534 2195 4568 2229
rect 4534 2127 4568 2161
rect 4534 2059 4568 2093
rect 4534 1991 4568 2025
rect 4534 1923 4568 1957
rect 4534 1855 4568 1889
rect 4630 2739 4664 2773
rect 4630 2671 4664 2705
rect 4630 2603 4664 2637
rect 4630 2535 4664 2569
rect 4630 2467 4664 2501
rect 4630 2399 4664 2433
rect 4630 2331 4664 2365
rect 4630 2263 4664 2297
rect 4630 2195 4664 2229
rect 4630 2127 4664 2161
rect 4630 2059 4664 2093
rect 4630 1991 4664 2025
rect 4630 1923 4664 1957
rect 4630 1855 4664 1889
rect 4726 2739 4760 2773
rect 4726 2671 4760 2705
rect 4726 2603 4760 2637
rect 4726 2535 4760 2569
rect 4726 2467 4760 2501
rect 4726 2399 4760 2433
rect 4726 2331 4760 2365
rect 4726 2263 4760 2297
rect 4726 2195 4760 2229
rect 4726 2127 4760 2161
rect 4726 2059 4760 2093
rect 4726 1991 4760 2025
rect 4726 1923 4760 1957
rect 4726 1855 4760 1889
rect 4822 2739 4856 2773
rect 4822 2671 4856 2705
rect 4822 2603 4856 2637
rect 4822 2535 4856 2569
rect 4822 2467 4856 2501
rect 7468 2739 7502 2773
rect 7468 2671 7502 2705
rect 7468 2603 7502 2637
rect 7468 2535 7502 2569
rect 7468 2467 7502 2501
rect 4822 2399 4856 2433
rect 4822 2331 4856 2365
rect 4822 2263 4856 2297
rect 7468 2399 7502 2433
rect 7468 2331 7502 2365
rect 4822 2195 4856 2229
rect 4822 2127 4856 2161
rect 4822 2059 4856 2093
rect 5500 2227 5534 2261
rect 5500 2159 5534 2193
rect 5500 2091 5534 2125
rect 5658 2227 5692 2261
rect 5658 2159 5692 2193
rect 5658 2091 5692 2125
rect 7468 2263 7502 2297
rect 7468 2195 7502 2229
rect 7468 2127 7502 2161
rect 7468 2059 7502 2093
rect 4822 1991 4856 2025
rect 4822 1923 4856 1957
rect 4822 1855 4856 1889
rect 7468 1991 7502 2025
rect 7468 1923 7502 1957
rect 7468 1855 7502 1889
rect 7564 2739 7598 2773
rect 7564 2671 7598 2705
rect 7564 2603 7598 2637
rect 7564 2535 7598 2569
rect 7564 2467 7598 2501
rect 7564 2399 7598 2433
rect 7564 2331 7598 2365
rect 7564 2263 7598 2297
rect 7564 2195 7598 2229
rect 7564 2127 7598 2161
rect 7564 2059 7598 2093
rect 7564 1991 7598 2025
rect 7564 1923 7598 1957
rect 7564 1855 7598 1889
rect 7660 2739 7694 2773
rect 7660 2671 7694 2705
rect 7660 2603 7694 2637
rect 7660 2535 7694 2569
rect 7660 2467 7694 2501
rect 7660 2399 7694 2433
rect 7660 2331 7694 2365
rect 7660 2263 7694 2297
rect 7660 2195 7694 2229
rect 7660 2127 7694 2161
rect 7660 2059 7694 2093
rect 7660 1991 7694 2025
rect 7660 1923 7694 1957
rect 7660 1855 7694 1889
rect 7756 2739 7790 2773
rect 7756 2671 7790 2705
rect 7756 2603 7790 2637
rect 7756 2535 7790 2569
rect 7756 2467 7790 2501
rect 7756 2399 7790 2433
rect 7756 2331 7790 2365
rect 7756 2263 7790 2297
rect 7756 2195 7790 2229
rect 7756 2127 7790 2161
rect 7756 2059 7790 2093
rect 7756 1991 7790 2025
rect 7756 1923 7790 1957
rect 7756 1855 7790 1889
rect 7852 2739 7886 2773
rect 7852 2671 7886 2705
rect 7852 2603 7886 2637
rect 7852 2535 7886 2569
rect 7852 2467 7886 2501
rect 10556 2737 10590 2771
rect 10556 2669 10590 2703
rect 10556 2601 10590 2635
rect 10556 2533 10590 2567
rect 10556 2465 10590 2499
rect 7852 2399 7886 2433
rect 7852 2331 7886 2365
rect 7852 2263 7886 2297
rect 10556 2397 10590 2431
rect 10556 2329 10590 2363
rect 7852 2195 7886 2229
rect 7852 2127 7886 2161
rect 7852 2059 7886 2093
rect 8500 2227 8534 2261
rect 8500 2159 8534 2193
rect 8500 2091 8534 2125
rect 8658 2227 8692 2261
rect 8658 2159 8692 2193
rect 8658 2091 8692 2125
rect 10556 2261 10590 2295
rect 10556 2193 10590 2227
rect 10556 2125 10590 2159
rect 10556 2057 10590 2091
rect 7852 1991 7886 2025
rect 7852 1923 7886 1957
rect 7852 1855 7886 1889
rect 10556 1989 10590 2023
rect 10556 1921 10590 1955
rect 10556 1853 10590 1887
rect 10652 2737 10686 2771
rect 10652 2669 10686 2703
rect 10652 2601 10686 2635
rect 10652 2533 10686 2567
rect 10652 2465 10686 2499
rect 10652 2397 10686 2431
rect 10652 2329 10686 2363
rect 10652 2261 10686 2295
rect 10652 2193 10686 2227
rect 10652 2125 10686 2159
rect 10652 2057 10686 2091
rect 10652 1989 10686 2023
rect 10652 1921 10686 1955
rect 10652 1853 10686 1887
rect 10748 2737 10782 2771
rect 10748 2669 10782 2703
rect 10748 2601 10782 2635
rect 10748 2533 10782 2567
rect 10748 2465 10782 2499
rect 10748 2397 10782 2431
rect 10748 2329 10782 2363
rect 10748 2261 10782 2295
rect 10748 2193 10782 2227
rect 10748 2125 10782 2159
rect 10748 2057 10782 2091
rect 10748 1989 10782 2023
rect 10748 1921 10782 1955
rect 10748 1853 10782 1887
rect 10844 2737 10878 2771
rect 10844 2669 10878 2703
rect 10844 2601 10878 2635
rect 10844 2533 10878 2567
rect 10844 2465 10878 2499
rect 10844 2397 10878 2431
rect 10844 2329 10878 2363
rect 10844 2261 10878 2295
rect 10844 2193 10878 2227
rect 10844 2125 10878 2159
rect 10844 2057 10878 2091
rect 10844 1989 10878 2023
rect 10844 1921 10878 1955
rect 10844 1853 10878 1887
rect 16686 2847 16720 2881
rect 10940 2737 10974 2771
rect 10940 2669 10974 2703
rect 10940 2601 10974 2635
rect 10940 2533 10974 2567
rect 10940 2465 10974 2499
rect 13712 2711 13746 2745
rect 13712 2643 13746 2677
rect 13712 2575 13746 2609
rect 13712 2507 13746 2541
rect 10940 2397 10974 2431
rect 10940 2329 10974 2363
rect 10940 2261 10974 2295
rect 13712 2439 13746 2473
rect 13712 2371 13746 2405
rect 13712 2303 13746 2337
rect 10940 2193 10974 2227
rect 10940 2125 10974 2159
rect 10940 2057 10974 2091
rect 11500 2227 11534 2261
rect 11500 2159 11534 2193
rect 11500 2091 11534 2125
rect 11658 2227 11692 2261
rect 11658 2159 11692 2193
rect 11658 2091 11692 2125
rect 13712 2235 13746 2269
rect 13712 2167 13746 2201
rect 13712 2099 13746 2133
rect 10940 1989 10974 2023
rect 10940 1921 10974 1955
rect 10940 1853 10974 1887
rect 13712 2031 13746 2065
rect 13712 1963 13746 1997
rect 13712 1895 13746 1929
rect 13712 1827 13746 1861
rect 13808 2711 13842 2745
rect 13808 2643 13842 2677
rect 13808 2575 13842 2609
rect 13808 2507 13842 2541
rect 13808 2439 13842 2473
rect 13808 2371 13842 2405
rect 13808 2303 13842 2337
rect 13808 2235 13842 2269
rect 13808 2167 13842 2201
rect 13808 2099 13842 2133
rect 13808 2031 13842 2065
rect 13808 1963 13842 1997
rect 13808 1895 13842 1929
rect 13808 1827 13842 1861
rect 13904 2711 13938 2745
rect 13904 2643 13938 2677
rect 13904 2575 13938 2609
rect 13904 2507 13938 2541
rect 13904 2439 13938 2473
rect 13904 2371 13938 2405
rect 13904 2303 13938 2337
rect 13904 2235 13938 2269
rect 13904 2167 13938 2201
rect 13904 2099 13938 2133
rect 13904 2031 13938 2065
rect 13904 1963 13938 1997
rect 13904 1895 13938 1929
rect 13904 1827 13938 1861
rect 14000 2711 14034 2745
rect 14000 2643 14034 2677
rect 14000 2575 14034 2609
rect 14000 2507 14034 2541
rect 14000 2439 14034 2473
rect 14000 2371 14034 2405
rect 14000 2303 14034 2337
rect 14000 2235 14034 2269
rect 14000 2167 14034 2201
rect 14000 2099 14034 2133
rect 14000 2031 14034 2065
rect 14000 1963 14034 1997
rect 14000 1895 14034 1929
rect 14000 1827 14034 1861
rect 14096 2711 14130 2745
rect 14096 2643 14130 2677
rect 14096 2575 14130 2609
rect 14096 2507 14130 2541
rect 16686 2779 16720 2813
rect 16686 2711 16720 2745
rect 16686 2643 16720 2677
rect 16686 2575 16720 2609
rect 16782 3459 16816 3493
rect 16782 3391 16816 3425
rect 16782 3323 16816 3357
rect 16782 3255 16816 3289
rect 16782 3187 16816 3221
rect 16782 3119 16816 3153
rect 16782 3051 16816 3085
rect 16782 2983 16816 3017
rect 16782 2915 16816 2949
rect 16782 2847 16816 2881
rect 16782 2779 16816 2813
rect 16782 2711 16816 2745
rect 16782 2643 16816 2677
rect 16782 2575 16816 2609
rect 16878 3459 16912 3493
rect 16878 3391 16912 3425
rect 16878 3323 16912 3357
rect 16878 3255 16912 3289
rect 16878 3187 16912 3221
rect 16878 3119 16912 3153
rect 16878 3051 16912 3085
rect 16878 2983 16912 3017
rect 16878 2915 16912 2949
rect 16878 2847 16912 2881
rect 16878 2779 16912 2813
rect 16878 2711 16912 2745
rect 16878 2643 16912 2677
rect 16878 2575 16912 2609
rect 16974 3459 17008 3493
rect 16974 3391 17008 3425
rect 16974 3323 17008 3357
rect 16974 3255 17008 3289
rect 16974 3187 17008 3221
rect 16974 3119 17008 3153
rect 16974 3051 17008 3085
rect 16974 2983 17008 3017
rect 16974 2915 17008 2949
rect 16974 2847 17008 2881
rect 16974 2779 17008 2813
rect 16974 2711 17008 2745
rect 16974 2643 17008 2677
rect 16974 2575 17008 2609
rect 17070 3459 17104 3493
rect 17070 3391 17104 3425
rect 17070 3323 17104 3357
rect 17070 3255 17104 3289
rect 17070 3187 17104 3221
rect 17070 3119 17104 3153
rect 17070 3051 17104 3085
rect 17070 2983 17104 3017
rect 17070 2915 17104 2949
rect 17070 2847 17104 2881
rect 17070 2779 17104 2813
rect 17070 2711 17104 2745
rect 17070 2643 17104 2677
rect 17070 2575 17104 2609
rect 17166 3459 17200 3493
rect 17166 3391 17200 3425
rect 17166 3323 17200 3357
rect 17166 3255 17200 3289
rect 17166 3187 17200 3221
rect 17166 3119 17200 3153
rect 17166 3051 17200 3085
rect 17166 2983 17200 3017
rect 17166 2915 17200 2949
rect 17166 2847 17200 2881
rect 17166 2779 17200 2813
rect 17166 2711 17200 2745
rect 17166 2643 17200 2677
rect 17166 2575 17200 2609
rect 17378 3449 17412 3483
rect 17378 3381 17412 3415
rect 17378 3313 17412 3347
rect 17378 3245 17412 3279
rect 17378 3177 17412 3211
rect 17378 3109 17412 3143
rect 17378 3041 17412 3075
rect 17378 2973 17412 3007
rect 17378 2905 17412 2939
rect 17378 2837 17412 2871
rect 17378 2769 17412 2803
rect 17378 2701 17412 2735
rect 17378 2633 17412 2667
rect 17378 2565 17412 2599
rect 17474 3449 17508 3483
rect 17474 3381 17508 3415
rect 17474 3313 17508 3347
rect 17474 3245 17508 3279
rect 17474 3177 17508 3211
rect 17474 3109 17508 3143
rect 17474 3041 17508 3075
rect 17474 2973 17508 3007
rect 17474 2905 17508 2939
rect 17474 2837 17508 2871
rect 17474 2769 17508 2803
rect 17474 2701 17508 2735
rect 17474 2633 17508 2667
rect 17474 2565 17508 2599
rect 17570 3449 17604 3483
rect 17570 3381 17604 3415
rect 17570 3313 17604 3347
rect 17570 3245 17604 3279
rect 17570 3177 17604 3211
rect 17570 3109 17604 3143
rect 17570 3041 17604 3075
rect 17570 2973 17604 3007
rect 17570 2905 17604 2939
rect 17570 2837 17604 2871
rect 17570 2769 17604 2803
rect 17570 2701 17604 2735
rect 17570 2633 17604 2667
rect 17570 2565 17604 2599
rect 17666 3449 17700 3483
rect 17666 3381 17700 3415
rect 17666 3313 17700 3347
rect 17666 3245 17700 3279
rect 17666 3177 17700 3211
rect 17666 3109 17700 3143
rect 17666 3041 17700 3075
rect 17666 2973 17700 3007
rect 17666 2905 17700 2939
rect 17666 2837 17700 2871
rect 17666 2769 17700 2803
rect 17666 2701 17700 2735
rect 17666 2633 17700 2667
rect 17666 2565 17700 2599
rect 17762 3449 17796 3483
rect 17762 3381 17796 3415
rect 17762 3313 17796 3347
rect 17762 3245 17796 3279
rect 17762 3177 17796 3211
rect 17762 3109 17796 3143
rect 17762 3041 17796 3075
rect 17762 2973 17796 3007
rect 17762 2905 17796 2939
rect 17762 2837 17796 2871
rect 17762 2769 17796 2803
rect 17762 2701 17796 2735
rect 17762 2633 17796 2667
rect 17762 2565 17796 2599
rect 17858 3449 17892 3483
rect 17858 3381 17892 3415
rect 17858 3313 17892 3347
rect 17858 3245 17892 3279
rect 17858 3177 17892 3211
rect 17858 3109 17892 3143
rect 17858 3041 17892 3075
rect 17858 2973 17892 3007
rect 17858 2905 17892 2939
rect 17858 2837 17892 2871
rect 17858 2769 17892 2803
rect 17858 2701 17892 2735
rect 17858 2633 17892 2667
rect 17858 2565 17892 2599
rect 17954 3449 17988 3483
rect 17954 3381 17988 3415
rect 17954 3313 17988 3347
rect 17954 3245 17988 3279
rect 17954 3177 17988 3211
rect 17954 3109 17988 3143
rect 17954 3041 17988 3075
rect 17954 2973 17988 3007
rect 17954 2905 17988 2939
rect 17954 2837 17988 2871
rect 17954 2769 17988 2803
rect 17954 2701 17988 2735
rect 17954 2633 17988 2667
rect 17954 2565 17988 2599
rect 18050 3449 18084 3483
rect 18050 3381 18084 3415
rect 18050 3313 18084 3347
rect 18050 3245 18084 3279
rect 18050 3177 18084 3211
rect 18050 3109 18084 3143
rect 18050 3041 18084 3075
rect 18050 2973 18084 3007
rect 18050 2905 18084 2939
rect 18050 2837 18084 2871
rect 18050 2769 18084 2803
rect 18050 2701 18084 2735
rect 18050 2633 18084 2667
rect 18050 2565 18084 2599
rect 18146 3449 18180 3483
rect 18146 3381 18180 3415
rect 18146 3313 18180 3347
rect 18146 3245 18180 3279
rect 18146 3177 18180 3211
rect 18146 3109 18180 3143
rect 18146 3041 18180 3075
rect 18146 2973 18180 3007
rect 18146 2905 18180 2939
rect 18146 2837 18180 2871
rect 18146 2769 18180 2803
rect 18146 2701 18180 2735
rect 18146 2633 18180 2667
rect 18146 2565 18180 2599
rect 18242 3449 18276 3483
rect 18242 3381 18276 3415
rect 18242 3313 18276 3347
rect 18242 3245 18276 3279
rect 18242 3177 18276 3211
rect 18242 3109 18276 3143
rect 18242 3041 18276 3075
rect 18242 2973 18276 3007
rect 18242 2905 18276 2939
rect 18242 2837 18276 2871
rect 18242 2769 18276 2803
rect 18242 2701 18276 2735
rect 18242 2633 18276 2667
rect 18242 2565 18276 2599
rect 18338 3449 18372 3483
rect 18338 3381 18372 3415
rect 18338 3313 18372 3347
rect 18338 3245 18372 3279
rect 18338 3177 18372 3211
rect 18338 3109 18372 3143
rect 18338 3041 18372 3075
rect 18338 2973 18372 3007
rect 18338 2905 18372 2939
rect 18338 2837 18372 2871
rect 18338 2769 18372 2803
rect 18338 2701 18372 2735
rect 18338 2633 18372 2667
rect 18338 2565 18372 2599
rect 18576 3445 18610 3479
rect 18576 3377 18610 3411
rect 18576 3309 18610 3343
rect 18576 3241 18610 3275
rect 18576 3173 18610 3207
rect 18576 3105 18610 3139
rect 18576 3037 18610 3071
rect 18576 2969 18610 3003
rect 18576 2901 18610 2935
rect 18576 2833 18610 2867
rect 18576 2765 18610 2799
rect 18576 2697 18610 2731
rect 18576 2629 18610 2663
rect 18576 2561 18610 2595
rect 18672 3445 18706 3479
rect 18672 3377 18706 3411
rect 18672 3309 18706 3343
rect 18672 3241 18706 3275
rect 18672 3173 18706 3207
rect 18672 3105 18706 3139
rect 18672 3037 18706 3071
rect 18672 2969 18706 3003
rect 18672 2901 18706 2935
rect 18672 2833 18706 2867
rect 18672 2765 18706 2799
rect 18672 2697 18706 2731
rect 18672 2629 18706 2663
rect 18672 2561 18706 2595
rect 18768 3445 18802 3479
rect 18768 3377 18802 3411
rect 18768 3309 18802 3343
rect 18768 3241 18802 3275
rect 18768 3173 18802 3207
rect 18768 3105 18802 3139
rect 18768 3037 18802 3071
rect 18768 2969 18802 3003
rect 18768 2901 18802 2935
rect 18768 2833 18802 2867
rect 18768 2765 18802 2799
rect 18768 2697 18802 2731
rect 18768 2629 18802 2663
rect 18768 2561 18802 2595
rect 18864 3445 18898 3479
rect 18864 3377 18898 3411
rect 18864 3309 18898 3343
rect 18864 3241 18898 3275
rect 18864 3173 18898 3207
rect 18864 3105 18898 3139
rect 18864 3037 18898 3071
rect 18864 2969 18898 3003
rect 18864 2901 18898 2935
rect 18864 2833 18898 2867
rect 18864 2765 18898 2799
rect 18864 2697 18898 2731
rect 18864 2629 18898 2663
rect 18864 2561 18898 2595
rect 18960 3445 18994 3479
rect 18960 3377 18994 3411
rect 18960 3309 18994 3343
rect 18960 3241 18994 3275
rect 18960 3173 18994 3207
rect 18960 3105 18994 3139
rect 18960 3037 18994 3071
rect 18960 2969 18994 3003
rect 18960 2901 18994 2935
rect 18960 2833 18994 2867
rect 18960 2765 18994 2799
rect 18960 2697 18994 2731
rect 18960 2629 18994 2663
rect 18960 2561 18994 2595
rect 19056 3445 19090 3479
rect 19056 3377 19090 3411
rect 19056 3309 19090 3343
rect 19056 3241 19090 3275
rect 19056 3173 19090 3207
rect 19056 3105 19090 3139
rect 19056 3037 19090 3071
rect 19056 2969 19090 3003
rect 19056 2901 19090 2935
rect 19056 2833 19090 2867
rect 19056 2765 19090 2799
rect 19056 2697 19090 2731
rect 19056 2629 19090 2663
rect 19056 2561 19090 2595
rect 19152 3445 19186 3479
rect 19152 3377 19186 3411
rect 19152 3309 19186 3343
rect 19152 3241 19186 3275
rect 19152 3173 19186 3207
rect 19152 3105 19186 3139
rect 19152 3037 19186 3071
rect 19152 2969 19186 3003
rect 19152 2901 19186 2935
rect 19152 2833 19186 2867
rect 19152 2765 19186 2799
rect 19152 2697 19186 2731
rect 19152 2629 19186 2663
rect 19152 2561 19186 2595
rect 19248 3445 19282 3479
rect 19248 3377 19282 3411
rect 19248 3309 19282 3343
rect 19248 3241 19282 3275
rect 19248 3173 19282 3207
rect 19248 3105 19282 3139
rect 19248 3037 19282 3071
rect 19248 2969 19282 3003
rect 19248 2901 19282 2935
rect 19248 2833 19282 2867
rect 19248 2765 19282 2799
rect 19248 2697 19282 2731
rect 19248 2629 19282 2663
rect 19248 2561 19282 2595
rect 19344 3445 19378 3479
rect 19344 3377 19378 3411
rect 19344 3309 19378 3343
rect 19344 3241 19378 3275
rect 19344 3173 19378 3207
rect 19344 3105 19378 3139
rect 19344 3037 19378 3071
rect 19344 2969 19378 3003
rect 19344 2901 19378 2935
rect 19344 2833 19378 2867
rect 19344 2765 19378 2799
rect 19344 2697 19378 2731
rect 19344 2629 19378 2663
rect 19344 2561 19378 2595
rect 19440 3445 19474 3479
rect 19440 3377 19474 3411
rect 19440 3309 19474 3343
rect 19440 3241 19474 3275
rect 19440 3173 19474 3207
rect 19440 3105 19474 3139
rect 19440 3037 19474 3071
rect 19440 2969 19474 3003
rect 19440 2901 19474 2935
rect 19440 2833 19474 2867
rect 19440 2765 19474 2799
rect 19440 2697 19474 2731
rect 19440 2629 19474 2663
rect 19440 2561 19474 2595
rect 19536 3445 19570 3479
rect 19536 3377 19570 3411
rect 19536 3309 19570 3343
rect 19536 3241 19570 3275
rect 19536 3173 19570 3207
rect 19536 3105 19570 3139
rect 19536 3037 19570 3071
rect 19536 2969 19570 3003
rect 19536 2901 19570 2935
rect 19536 2833 19570 2867
rect 19536 2765 19570 2799
rect 19536 2697 19570 2731
rect 19536 2629 19570 2663
rect 19536 2561 19570 2595
rect 19632 3445 19666 3479
rect 19632 3377 19666 3411
rect 19632 3309 19666 3343
rect 19632 3241 19666 3275
rect 19632 3173 19666 3207
rect 19632 3105 19666 3139
rect 19632 3037 19666 3071
rect 19632 2969 19666 3003
rect 19632 2901 19666 2935
rect 19632 2833 19666 2867
rect 19632 2765 19666 2799
rect 19632 2697 19666 2731
rect 19632 2629 19666 2663
rect 19632 2561 19666 2595
rect 19728 3445 19762 3479
rect 19728 3377 19762 3411
rect 19728 3309 19762 3343
rect 19728 3241 19762 3275
rect 19728 3173 19762 3207
rect 19728 3105 19762 3139
rect 19728 3037 19762 3071
rect 19728 2969 19762 3003
rect 19728 2901 19762 2935
rect 19728 2833 19762 2867
rect 19728 2765 19762 2799
rect 19728 2697 19762 2731
rect 19728 2629 19762 2663
rect 19728 2561 19762 2595
rect 19824 3445 19858 3479
rect 19824 3377 19858 3411
rect 19824 3309 19858 3343
rect 19824 3241 19858 3275
rect 19824 3173 19858 3207
rect 19824 3105 19858 3139
rect 19824 3037 19858 3071
rect 19824 2969 19858 3003
rect 19824 2901 19858 2935
rect 19824 2833 19858 2867
rect 19824 2765 19858 2799
rect 19824 2697 19858 2731
rect 19824 2629 19858 2663
rect 19824 2561 19858 2595
rect 19920 3445 19954 3479
rect 19920 3377 19954 3411
rect 19920 3309 19954 3343
rect 19920 3241 19954 3275
rect 19920 3173 19954 3207
rect 19920 3105 19954 3139
rect 19920 3037 19954 3071
rect 19920 2969 19954 3003
rect 19920 2901 19954 2935
rect 19920 2833 19954 2867
rect 19920 2765 19954 2799
rect 19920 2697 19954 2731
rect 19920 2629 19954 2663
rect 19920 2561 19954 2595
rect 20016 3445 20050 3479
rect 20016 3377 20050 3411
rect 20016 3309 20050 3343
rect 20016 3241 20050 3275
rect 20016 3173 20050 3207
rect 20016 3105 20050 3139
rect 20016 3037 20050 3071
rect 20016 2969 20050 3003
rect 20016 2901 20050 2935
rect 20016 2833 20050 2867
rect 20016 2765 20050 2799
rect 20016 2697 20050 2731
rect 20016 2629 20050 2663
rect 20016 2561 20050 2595
rect 20244 3453 20278 3487
rect 20244 3385 20278 3419
rect 20244 3317 20278 3351
rect 20244 3249 20278 3283
rect 20244 3181 20278 3215
rect 20244 3113 20278 3147
rect 20244 3045 20278 3079
rect 20244 2977 20278 3011
rect 20244 2909 20278 2943
rect 20244 2841 20278 2875
rect 20244 2773 20278 2807
rect 20244 2705 20278 2739
rect 20244 2637 20278 2671
rect 20244 2569 20278 2603
rect 20340 3453 20374 3487
rect 20340 3385 20374 3419
rect 20340 3317 20374 3351
rect 20340 3249 20374 3283
rect 20340 3181 20374 3215
rect 20340 3113 20374 3147
rect 20340 3045 20374 3079
rect 20340 2977 20374 3011
rect 20340 2909 20374 2943
rect 20340 2841 20374 2875
rect 20340 2773 20374 2807
rect 20340 2705 20374 2739
rect 20340 2637 20374 2671
rect 20340 2569 20374 2603
rect 20436 3453 20470 3487
rect 20436 3385 20470 3419
rect 20436 3317 20470 3351
rect 20436 3249 20470 3283
rect 20436 3181 20470 3215
rect 20436 3113 20470 3147
rect 20436 3045 20470 3079
rect 20436 2977 20470 3011
rect 20436 2909 20470 2943
rect 20436 2841 20470 2875
rect 20436 2773 20470 2807
rect 20436 2705 20470 2739
rect 20436 2637 20470 2671
rect 20436 2569 20470 2603
rect 20532 3453 20566 3487
rect 20532 3385 20566 3419
rect 20532 3317 20566 3351
rect 20532 3249 20566 3283
rect 20532 3181 20566 3215
rect 20532 3113 20566 3147
rect 20532 3045 20566 3079
rect 20532 2977 20566 3011
rect 20532 2909 20566 2943
rect 20532 2841 20566 2875
rect 20532 2773 20566 2807
rect 20532 2705 20566 2739
rect 20532 2637 20566 2671
rect 20532 2569 20566 2603
rect 20628 3453 20662 3487
rect 20628 3385 20662 3419
rect 20628 3317 20662 3351
rect 20628 3249 20662 3283
rect 20628 3181 20662 3215
rect 20628 3113 20662 3147
rect 20628 3045 20662 3079
rect 20628 2977 20662 3011
rect 20628 2909 20662 2943
rect 20628 2841 20662 2875
rect 20628 2773 20662 2807
rect 20628 2705 20662 2739
rect 20628 2637 20662 2671
rect 20628 2569 20662 2603
rect 20724 3453 20758 3487
rect 20724 3385 20758 3419
rect 20724 3317 20758 3351
rect 20724 3249 20758 3283
rect 20724 3181 20758 3215
rect 20724 3113 20758 3147
rect 20724 3045 20758 3079
rect 20724 2977 20758 3011
rect 20724 2909 20758 2943
rect 20724 2841 20758 2875
rect 20724 2773 20758 2807
rect 20724 2705 20758 2739
rect 20724 2637 20758 2671
rect 20724 2569 20758 2603
rect 20820 3453 20854 3487
rect 20820 3385 20854 3419
rect 20820 3317 20854 3351
rect 20820 3249 20854 3283
rect 20820 3181 20854 3215
rect 20820 3113 20854 3147
rect 20820 3045 20854 3079
rect 20820 2977 20854 3011
rect 20820 2909 20854 2943
rect 20820 2841 20854 2875
rect 20820 2773 20854 2807
rect 20820 2705 20854 2739
rect 20820 2637 20854 2671
rect 20820 2569 20854 2603
rect 20916 3453 20950 3487
rect 20916 3385 20950 3419
rect 20916 3317 20950 3351
rect 20916 3249 20950 3283
rect 20916 3181 20950 3215
rect 20916 3113 20950 3147
rect 20916 3045 20950 3079
rect 20916 2977 20950 3011
rect 20916 2909 20950 2943
rect 20916 2841 20950 2875
rect 20916 2773 20950 2807
rect 20916 2705 20950 2739
rect 20916 2637 20950 2671
rect 20916 2569 20950 2603
rect 21012 3453 21046 3487
rect 21012 3385 21046 3419
rect 21012 3317 21046 3351
rect 21012 3249 21046 3283
rect 21012 3181 21046 3215
rect 21012 3113 21046 3147
rect 21012 3045 21046 3079
rect 21012 2977 21046 3011
rect 21012 2909 21046 2943
rect 21012 2841 21046 2875
rect 21012 2773 21046 2807
rect 21012 2705 21046 2739
rect 21012 2637 21046 2671
rect 21012 2569 21046 2603
rect 21108 3453 21142 3487
rect 21108 3385 21142 3419
rect 21108 3317 21142 3351
rect 21108 3249 21142 3283
rect 21108 3181 21142 3215
rect 21108 3113 21142 3147
rect 21108 3045 21142 3079
rect 21108 2977 21142 3011
rect 21108 2909 21142 2943
rect 21108 2841 21142 2875
rect 21108 2773 21142 2807
rect 21108 2705 21142 2739
rect 21108 2637 21142 2671
rect 21108 2569 21142 2603
rect 21204 3453 21238 3487
rect 21204 3385 21238 3419
rect 21204 3317 21238 3351
rect 21204 3249 21238 3283
rect 21204 3181 21238 3215
rect 21204 3113 21238 3147
rect 21204 3045 21238 3079
rect 21204 2977 21238 3011
rect 21204 2909 21238 2943
rect 21204 2841 21238 2875
rect 21204 2773 21238 2807
rect 21204 2705 21238 2739
rect 21204 2637 21238 2671
rect 21204 2569 21238 2603
rect 21300 3453 21334 3487
rect 21300 3385 21334 3419
rect 21300 3317 21334 3351
rect 21300 3249 21334 3283
rect 21300 3181 21334 3215
rect 21300 3113 21334 3147
rect 21300 3045 21334 3079
rect 21300 2977 21334 3011
rect 21300 2909 21334 2943
rect 21300 2841 21334 2875
rect 21300 2773 21334 2807
rect 21300 2705 21334 2739
rect 21300 2637 21334 2671
rect 21300 2569 21334 2603
rect 21396 3453 21430 3487
rect 21396 3385 21430 3419
rect 21396 3317 21430 3351
rect 21396 3249 21430 3283
rect 21396 3181 21430 3215
rect 21396 3113 21430 3147
rect 21396 3045 21430 3079
rect 21396 2977 21430 3011
rect 21396 2909 21430 2943
rect 21396 2841 21430 2875
rect 21396 2773 21430 2807
rect 21396 2705 21430 2739
rect 21396 2637 21430 2671
rect 21396 2569 21430 2603
rect 21492 3453 21526 3487
rect 21492 3385 21526 3419
rect 21492 3317 21526 3351
rect 21492 3249 21526 3283
rect 21492 3181 21526 3215
rect 21492 3113 21526 3147
rect 21492 3045 21526 3079
rect 21492 2977 21526 3011
rect 21492 2909 21526 2943
rect 21492 2841 21526 2875
rect 21492 2773 21526 2807
rect 21492 2705 21526 2739
rect 21492 2637 21526 2671
rect 21492 2569 21526 2603
rect 21588 3453 21622 3487
rect 21588 3385 21622 3419
rect 21588 3317 21622 3351
rect 21588 3249 21622 3283
rect 21588 3181 21622 3215
rect 21588 3113 21622 3147
rect 21588 3045 21622 3079
rect 21588 2977 21622 3011
rect 21588 2909 21622 2943
rect 21588 2841 21622 2875
rect 21588 2773 21622 2807
rect 21588 2705 21622 2739
rect 21588 2637 21622 2671
rect 21588 2569 21622 2603
rect 21684 3453 21718 3487
rect 21684 3385 21718 3419
rect 21684 3317 21718 3351
rect 21684 3249 21718 3283
rect 21684 3181 21718 3215
rect 21684 3113 21718 3147
rect 21684 3045 21718 3079
rect 21684 2977 21718 3011
rect 21684 2909 21718 2943
rect 21684 2841 21718 2875
rect 21684 2773 21718 2807
rect 21684 2705 21718 2739
rect 21684 2637 21718 2671
rect 21684 2569 21718 2603
rect 21780 3453 21814 3487
rect 21780 3385 21814 3419
rect 21780 3317 21814 3351
rect 21780 3249 21814 3283
rect 21780 3181 21814 3215
rect 21780 3113 21814 3147
rect 21780 3045 21814 3079
rect 21780 2977 21814 3011
rect 21780 2909 21814 2943
rect 21780 2841 21814 2875
rect 21780 2773 21814 2807
rect 21780 2705 21814 2739
rect 21780 2637 21814 2671
rect 21780 2569 21814 2603
rect 21876 3453 21910 3487
rect 21876 3385 21910 3419
rect 21876 3317 21910 3351
rect 21876 3249 21910 3283
rect 21876 3181 21910 3215
rect 21876 3113 21910 3147
rect 21876 3045 21910 3079
rect 21876 2977 21910 3011
rect 21876 2909 21910 2943
rect 21876 2841 21910 2875
rect 21876 2773 21910 2807
rect 21876 2705 21910 2739
rect 21876 2637 21910 2671
rect 21876 2569 21910 2603
rect 21972 3453 22006 3487
rect 21972 3385 22006 3419
rect 21972 3317 22006 3351
rect 21972 3249 22006 3283
rect 21972 3181 22006 3215
rect 21972 3113 22006 3147
rect 21972 3045 22006 3079
rect 21972 2977 22006 3011
rect 21972 2909 22006 2943
rect 21972 2841 22006 2875
rect 21972 2773 22006 2807
rect 21972 2705 22006 2739
rect 21972 2637 22006 2671
rect 21972 2569 22006 2603
rect 22068 3453 22102 3487
rect 22068 3385 22102 3419
rect 22068 3317 22102 3351
rect 22068 3249 22102 3283
rect 22068 3181 22102 3215
rect 22068 3113 22102 3147
rect 22068 3045 22102 3079
rect 22068 2977 22102 3011
rect 22068 2909 22102 2943
rect 22068 2841 22102 2875
rect 22068 2773 22102 2807
rect 22068 2705 22102 2739
rect 22068 2637 22102 2671
rect 22068 2569 22102 2603
rect 22164 3453 22198 3487
rect 22164 3385 22198 3419
rect 22164 3317 22198 3351
rect 22164 3249 22198 3283
rect 22164 3181 22198 3215
rect 22164 3113 22198 3147
rect 22164 3045 22198 3079
rect 22164 2977 22198 3011
rect 22164 2909 22198 2943
rect 22164 2841 22198 2875
rect 22164 2773 22198 2807
rect 22164 2705 22198 2739
rect 22164 2637 22198 2671
rect 22164 2569 22198 2603
rect 23174 3457 23208 3491
rect 23174 3389 23208 3423
rect 23174 3321 23208 3355
rect 23174 3253 23208 3287
rect 23174 3185 23208 3219
rect 23174 3117 23208 3151
rect 23174 3049 23208 3083
rect 23174 2981 23208 3015
rect 23174 2913 23208 2947
rect 23174 2845 23208 2879
rect 23174 2777 23208 2811
rect 23174 2709 23208 2743
rect 23174 2641 23208 2675
rect 23174 2573 23208 2607
rect 23270 3457 23304 3491
rect 23270 3389 23304 3423
rect 23270 3321 23304 3355
rect 23270 3253 23304 3287
rect 23270 3185 23304 3219
rect 23270 3117 23304 3151
rect 23270 3049 23304 3083
rect 23270 2981 23304 3015
rect 23270 2913 23304 2947
rect 23270 2845 23304 2879
rect 23270 2777 23304 2811
rect 23270 2709 23304 2743
rect 23270 2641 23304 2675
rect 23270 2573 23304 2607
rect 23366 3457 23400 3491
rect 23366 3389 23400 3423
rect 23366 3321 23400 3355
rect 23366 3253 23400 3287
rect 23366 3185 23400 3219
rect 23366 3117 23400 3151
rect 23366 3049 23400 3083
rect 23366 2981 23400 3015
rect 23366 2913 23400 2947
rect 23366 2845 23400 2879
rect 23366 2777 23400 2811
rect 23366 2709 23400 2743
rect 23366 2641 23400 2675
rect 23366 2573 23400 2607
rect 23462 3457 23496 3491
rect 23462 3389 23496 3423
rect 23462 3321 23496 3355
rect 23462 3253 23496 3287
rect 23462 3185 23496 3219
rect 23462 3117 23496 3151
rect 23462 3049 23496 3083
rect 23462 2981 23496 3015
rect 23462 2913 23496 2947
rect 23462 2845 23496 2879
rect 23462 2777 23496 2811
rect 23462 2709 23496 2743
rect 23462 2641 23496 2675
rect 23462 2573 23496 2607
rect 23558 3457 23592 3491
rect 23558 3389 23592 3423
rect 23558 3321 23592 3355
rect 23558 3253 23592 3287
rect 23558 3185 23592 3219
rect 23558 3117 23592 3151
rect 23558 3049 23592 3083
rect 23558 2981 23592 3015
rect 23558 2913 23592 2947
rect 23558 2845 23592 2879
rect 23558 2777 23592 2811
rect 23558 2709 23592 2743
rect 23558 2641 23592 2675
rect 23558 2573 23592 2607
rect 23654 3457 23688 3491
rect 23654 3389 23688 3423
rect 23654 3321 23688 3355
rect 23654 3253 23688 3287
rect 23654 3185 23688 3219
rect 23654 3117 23688 3151
rect 23654 3049 23688 3083
rect 23654 2981 23688 3015
rect 23654 2913 23688 2947
rect 23654 2845 23688 2879
rect 23654 2777 23688 2811
rect 23654 2709 23688 2743
rect 23654 2641 23688 2675
rect 23654 2573 23688 2607
rect 23866 3447 23900 3481
rect 23866 3379 23900 3413
rect 23866 3311 23900 3345
rect 23866 3243 23900 3277
rect 23866 3175 23900 3209
rect 23866 3107 23900 3141
rect 23866 3039 23900 3073
rect 23866 2971 23900 3005
rect 23866 2903 23900 2937
rect 23866 2835 23900 2869
rect 23866 2767 23900 2801
rect 23866 2699 23900 2733
rect 23866 2631 23900 2665
rect 23866 2563 23900 2597
rect 23962 3447 23996 3481
rect 23962 3379 23996 3413
rect 23962 3311 23996 3345
rect 23962 3243 23996 3277
rect 23962 3175 23996 3209
rect 23962 3107 23996 3141
rect 23962 3039 23996 3073
rect 23962 2971 23996 3005
rect 23962 2903 23996 2937
rect 23962 2835 23996 2869
rect 23962 2767 23996 2801
rect 23962 2699 23996 2733
rect 23962 2631 23996 2665
rect 23962 2563 23996 2597
rect 24058 3447 24092 3481
rect 24058 3379 24092 3413
rect 24058 3311 24092 3345
rect 24058 3243 24092 3277
rect 24058 3175 24092 3209
rect 24058 3107 24092 3141
rect 24058 3039 24092 3073
rect 24058 2971 24092 3005
rect 24058 2903 24092 2937
rect 24058 2835 24092 2869
rect 24058 2767 24092 2801
rect 24058 2699 24092 2733
rect 24058 2631 24092 2665
rect 24058 2563 24092 2597
rect 24154 3447 24188 3481
rect 24154 3379 24188 3413
rect 24154 3311 24188 3345
rect 24154 3243 24188 3277
rect 24154 3175 24188 3209
rect 24154 3107 24188 3141
rect 24154 3039 24188 3073
rect 24154 2971 24188 3005
rect 24154 2903 24188 2937
rect 24154 2835 24188 2869
rect 24154 2767 24188 2801
rect 24154 2699 24188 2733
rect 24154 2631 24188 2665
rect 24154 2563 24188 2597
rect 24250 3447 24284 3481
rect 24250 3379 24284 3413
rect 24250 3311 24284 3345
rect 24250 3243 24284 3277
rect 24250 3175 24284 3209
rect 24250 3107 24284 3141
rect 24250 3039 24284 3073
rect 24250 2971 24284 3005
rect 24250 2903 24284 2937
rect 24250 2835 24284 2869
rect 24250 2767 24284 2801
rect 24250 2699 24284 2733
rect 24250 2631 24284 2665
rect 24250 2563 24284 2597
rect 24346 3447 24380 3481
rect 24346 3379 24380 3413
rect 24346 3311 24380 3345
rect 24346 3243 24380 3277
rect 24346 3175 24380 3209
rect 24346 3107 24380 3141
rect 24346 3039 24380 3073
rect 24346 2971 24380 3005
rect 24346 2903 24380 2937
rect 24346 2835 24380 2869
rect 24346 2767 24380 2801
rect 24346 2699 24380 2733
rect 24346 2631 24380 2665
rect 24346 2563 24380 2597
rect 24442 3447 24476 3481
rect 24442 3379 24476 3413
rect 24442 3311 24476 3345
rect 24442 3243 24476 3277
rect 24442 3175 24476 3209
rect 24442 3107 24476 3141
rect 24442 3039 24476 3073
rect 24442 2971 24476 3005
rect 24442 2903 24476 2937
rect 24442 2835 24476 2869
rect 24442 2767 24476 2801
rect 24442 2699 24476 2733
rect 24442 2631 24476 2665
rect 24442 2563 24476 2597
rect 24538 3447 24572 3481
rect 24538 3379 24572 3413
rect 24538 3311 24572 3345
rect 24538 3243 24572 3277
rect 24538 3175 24572 3209
rect 24538 3107 24572 3141
rect 24538 3039 24572 3073
rect 24538 2971 24572 3005
rect 24538 2903 24572 2937
rect 24538 2835 24572 2869
rect 24538 2767 24572 2801
rect 24538 2699 24572 2733
rect 24538 2631 24572 2665
rect 24538 2563 24572 2597
rect 24634 3447 24668 3481
rect 24634 3379 24668 3413
rect 24634 3311 24668 3345
rect 24634 3243 24668 3277
rect 24634 3175 24668 3209
rect 24634 3107 24668 3141
rect 24634 3039 24668 3073
rect 24634 2971 24668 3005
rect 24634 2903 24668 2937
rect 24634 2835 24668 2869
rect 24634 2767 24668 2801
rect 24634 2699 24668 2733
rect 24634 2631 24668 2665
rect 24634 2563 24668 2597
rect 24730 3447 24764 3481
rect 24730 3379 24764 3413
rect 24730 3311 24764 3345
rect 24730 3243 24764 3277
rect 24730 3175 24764 3209
rect 24730 3107 24764 3141
rect 24730 3039 24764 3073
rect 24730 2971 24764 3005
rect 24730 2903 24764 2937
rect 24730 2835 24764 2869
rect 24730 2767 24764 2801
rect 24730 2699 24764 2733
rect 24730 2631 24764 2665
rect 24730 2563 24764 2597
rect 24826 3447 24860 3481
rect 24826 3379 24860 3413
rect 24826 3311 24860 3345
rect 24826 3243 24860 3277
rect 24826 3175 24860 3209
rect 24826 3107 24860 3141
rect 24826 3039 24860 3073
rect 24826 2971 24860 3005
rect 24826 2903 24860 2937
rect 24826 2835 24860 2869
rect 24826 2767 24860 2801
rect 24826 2699 24860 2733
rect 24826 2631 24860 2665
rect 24826 2563 24860 2597
rect 25064 3443 25098 3477
rect 25064 3375 25098 3409
rect 25064 3307 25098 3341
rect 25064 3239 25098 3273
rect 25064 3171 25098 3205
rect 25064 3103 25098 3137
rect 25064 3035 25098 3069
rect 25064 2967 25098 3001
rect 25064 2899 25098 2933
rect 25064 2831 25098 2865
rect 25064 2763 25098 2797
rect 25064 2695 25098 2729
rect 25064 2627 25098 2661
rect 25064 2559 25098 2593
rect 25160 3443 25194 3477
rect 25160 3375 25194 3409
rect 25160 3307 25194 3341
rect 25160 3239 25194 3273
rect 25160 3171 25194 3205
rect 25160 3103 25194 3137
rect 25160 3035 25194 3069
rect 25160 2967 25194 3001
rect 25160 2899 25194 2933
rect 25160 2831 25194 2865
rect 25160 2763 25194 2797
rect 25160 2695 25194 2729
rect 25160 2627 25194 2661
rect 25160 2559 25194 2593
rect 25256 3443 25290 3477
rect 25256 3375 25290 3409
rect 25256 3307 25290 3341
rect 25256 3239 25290 3273
rect 25256 3171 25290 3205
rect 25256 3103 25290 3137
rect 25256 3035 25290 3069
rect 25256 2967 25290 3001
rect 25256 2899 25290 2933
rect 25256 2831 25290 2865
rect 25256 2763 25290 2797
rect 25256 2695 25290 2729
rect 25256 2627 25290 2661
rect 25256 2559 25290 2593
rect 25352 3443 25386 3477
rect 25352 3375 25386 3409
rect 25352 3307 25386 3341
rect 25352 3239 25386 3273
rect 25352 3171 25386 3205
rect 25352 3103 25386 3137
rect 25352 3035 25386 3069
rect 25352 2967 25386 3001
rect 25352 2899 25386 2933
rect 25352 2831 25386 2865
rect 25352 2763 25386 2797
rect 25352 2695 25386 2729
rect 25352 2627 25386 2661
rect 25352 2559 25386 2593
rect 25448 3443 25482 3477
rect 25448 3375 25482 3409
rect 25448 3307 25482 3341
rect 25448 3239 25482 3273
rect 25448 3171 25482 3205
rect 25448 3103 25482 3137
rect 25448 3035 25482 3069
rect 25448 2967 25482 3001
rect 25448 2899 25482 2933
rect 25448 2831 25482 2865
rect 25448 2763 25482 2797
rect 25448 2695 25482 2729
rect 25448 2627 25482 2661
rect 25448 2559 25482 2593
rect 25544 3443 25578 3477
rect 25544 3375 25578 3409
rect 25544 3307 25578 3341
rect 25544 3239 25578 3273
rect 25544 3171 25578 3205
rect 25544 3103 25578 3137
rect 25544 3035 25578 3069
rect 25544 2967 25578 3001
rect 25544 2899 25578 2933
rect 25544 2831 25578 2865
rect 25544 2763 25578 2797
rect 25544 2695 25578 2729
rect 25544 2627 25578 2661
rect 25544 2559 25578 2593
rect 25640 3443 25674 3477
rect 25640 3375 25674 3409
rect 25640 3307 25674 3341
rect 25640 3239 25674 3273
rect 25640 3171 25674 3205
rect 25640 3103 25674 3137
rect 25640 3035 25674 3069
rect 25640 2967 25674 3001
rect 25640 2899 25674 2933
rect 25640 2831 25674 2865
rect 25640 2763 25674 2797
rect 25640 2695 25674 2729
rect 25640 2627 25674 2661
rect 25640 2559 25674 2593
rect 25736 3443 25770 3477
rect 25736 3375 25770 3409
rect 25736 3307 25770 3341
rect 25736 3239 25770 3273
rect 25736 3171 25770 3205
rect 25736 3103 25770 3137
rect 25736 3035 25770 3069
rect 25736 2967 25770 3001
rect 25736 2899 25770 2933
rect 25736 2831 25770 2865
rect 25736 2763 25770 2797
rect 25736 2695 25770 2729
rect 25736 2627 25770 2661
rect 25736 2559 25770 2593
rect 25832 3443 25866 3477
rect 25832 3375 25866 3409
rect 25832 3307 25866 3341
rect 25832 3239 25866 3273
rect 25832 3171 25866 3205
rect 25832 3103 25866 3137
rect 25832 3035 25866 3069
rect 25832 2967 25866 3001
rect 25832 2899 25866 2933
rect 25832 2831 25866 2865
rect 25832 2763 25866 2797
rect 25832 2695 25866 2729
rect 25832 2627 25866 2661
rect 25832 2559 25866 2593
rect 25928 3443 25962 3477
rect 25928 3375 25962 3409
rect 25928 3307 25962 3341
rect 25928 3239 25962 3273
rect 25928 3171 25962 3205
rect 25928 3103 25962 3137
rect 25928 3035 25962 3069
rect 25928 2967 25962 3001
rect 25928 2899 25962 2933
rect 25928 2831 25962 2865
rect 25928 2763 25962 2797
rect 25928 2695 25962 2729
rect 25928 2627 25962 2661
rect 25928 2559 25962 2593
rect 26024 3443 26058 3477
rect 26024 3375 26058 3409
rect 26024 3307 26058 3341
rect 26024 3239 26058 3273
rect 26024 3171 26058 3205
rect 26024 3103 26058 3137
rect 26024 3035 26058 3069
rect 26024 2967 26058 3001
rect 26024 2899 26058 2933
rect 26024 2831 26058 2865
rect 26024 2763 26058 2797
rect 26024 2695 26058 2729
rect 26024 2627 26058 2661
rect 26024 2559 26058 2593
rect 26120 3443 26154 3477
rect 26120 3375 26154 3409
rect 26120 3307 26154 3341
rect 26120 3239 26154 3273
rect 26120 3171 26154 3205
rect 26120 3103 26154 3137
rect 26120 3035 26154 3069
rect 26120 2967 26154 3001
rect 26120 2899 26154 2933
rect 26120 2831 26154 2865
rect 26120 2763 26154 2797
rect 26120 2695 26154 2729
rect 26120 2627 26154 2661
rect 26120 2559 26154 2593
rect 26216 3443 26250 3477
rect 26216 3375 26250 3409
rect 26216 3307 26250 3341
rect 26216 3239 26250 3273
rect 26216 3171 26250 3205
rect 26216 3103 26250 3137
rect 26216 3035 26250 3069
rect 26216 2967 26250 3001
rect 26216 2899 26250 2933
rect 26216 2831 26250 2865
rect 26216 2763 26250 2797
rect 26216 2695 26250 2729
rect 26216 2627 26250 2661
rect 26216 2559 26250 2593
rect 26312 3443 26346 3477
rect 26312 3375 26346 3409
rect 26312 3307 26346 3341
rect 26312 3239 26346 3273
rect 26312 3171 26346 3205
rect 26312 3103 26346 3137
rect 26312 3035 26346 3069
rect 26312 2967 26346 3001
rect 26312 2899 26346 2933
rect 26312 2831 26346 2865
rect 26312 2763 26346 2797
rect 26312 2695 26346 2729
rect 26312 2627 26346 2661
rect 26312 2559 26346 2593
rect 26408 3443 26442 3477
rect 26408 3375 26442 3409
rect 26408 3307 26442 3341
rect 26408 3239 26442 3273
rect 26408 3171 26442 3205
rect 26408 3103 26442 3137
rect 26408 3035 26442 3069
rect 26408 2967 26442 3001
rect 26408 2899 26442 2933
rect 26408 2831 26442 2865
rect 26408 2763 26442 2797
rect 26408 2695 26442 2729
rect 26408 2627 26442 2661
rect 26408 2559 26442 2593
rect 26504 3443 26538 3477
rect 26504 3375 26538 3409
rect 26504 3307 26538 3341
rect 26504 3239 26538 3273
rect 26504 3171 26538 3205
rect 26504 3103 26538 3137
rect 26504 3035 26538 3069
rect 26504 2967 26538 3001
rect 26504 2899 26538 2933
rect 26504 2831 26538 2865
rect 26504 2763 26538 2797
rect 26504 2695 26538 2729
rect 26504 2627 26538 2661
rect 26504 2559 26538 2593
rect 26732 3451 26766 3485
rect 26732 3383 26766 3417
rect 26732 3315 26766 3349
rect 26732 3247 26766 3281
rect 26732 3179 26766 3213
rect 26732 3111 26766 3145
rect 26732 3043 26766 3077
rect 26732 2975 26766 3009
rect 26732 2907 26766 2941
rect 26732 2839 26766 2873
rect 26732 2771 26766 2805
rect 26732 2703 26766 2737
rect 26732 2635 26766 2669
rect 26732 2567 26766 2601
rect 26828 3451 26862 3485
rect 26828 3383 26862 3417
rect 26828 3315 26862 3349
rect 26828 3247 26862 3281
rect 26828 3179 26862 3213
rect 26828 3111 26862 3145
rect 26828 3043 26862 3077
rect 26828 2975 26862 3009
rect 26828 2907 26862 2941
rect 26828 2839 26862 2873
rect 26828 2771 26862 2805
rect 26828 2703 26862 2737
rect 26828 2635 26862 2669
rect 26828 2567 26862 2601
rect 26924 3451 26958 3485
rect 26924 3383 26958 3417
rect 26924 3315 26958 3349
rect 26924 3247 26958 3281
rect 26924 3179 26958 3213
rect 26924 3111 26958 3145
rect 26924 3043 26958 3077
rect 26924 2975 26958 3009
rect 26924 2907 26958 2941
rect 26924 2839 26958 2873
rect 26924 2771 26958 2805
rect 26924 2703 26958 2737
rect 26924 2635 26958 2669
rect 26924 2567 26958 2601
rect 27020 3451 27054 3485
rect 27020 3383 27054 3417
rect 27020 3315 27054 3349
rect 27020 3247 27054 3281
rect 27020 3179 27054 3213
rect 27020 3111 27054 3145
rect 27020 3043 27054 3077
rect 27020 2975 27054 3009
rect 27020 2907 27054 2941
rect 27020 2839 27054 2873
rect 27020 2771 27054 2805
rect 27020 2703 27054 2737
rect 27020 2635 27054 2669
rect 27020 2567 27054 2601
rect 27116 3451 27150 3485
rect 27116 3383 27150 3417
rect 27116 3315 27150 3349
rect 27116 3247 27150 3281
rect 27116 3179 27150 3213
rect 27116 3111 27150 3145
rect 27116 3043 27150 3077
rect 27116 2975 27150 3009
rect 27116 2907 27150 2941
rect 27116 2839 27150 2873
rect 27116 2771 27150 2805
rect 27116 2703 27150 2737
rect 27116 2635 27150 2669
rect 27116 2567 27150 2601
rect 27212 3451 27246 3485
rect 27212 3383 27246 3417
rect 27212 3315 27246 3349
rect 27212 3247 27246 3281
rect 27212 3179 27246 3213
rect 27212 3111 27246 3145
rect 27212 3043 27246 3077
rect 27212 2975 27246 3009
rect 27212 2907 27246 2941
rect 27212 2839 27246 2873
rect 27212 2771 27246 2805
rect 27212 2703 27246 2737
rect 27212 2635 27246 2669
rect 27212 2567 27246 2601
rect 27308 3451 27342 3485
rect 27308 3383 27342 3417
rect 27308 3315 27342 3349
rect 27308 3247 27342 3281
rect 27308 3179 27342 3213
rect 27308 3111 27342 3145
rect 27308 3043 27342 3077
rect 27308 2975 27342 3009
rect 27308 2907 27342 2941
rect 27308 2839 27342 2873
rect 27308 2771 27342 2805
rect 27308 2703 27342 2737
rect 27308 2635 27342 2669
rect 27308 2567 27342 2601
rect 27404 3451 27438 3485
rect 27404 3383 27438 3417
rect 27404 3315 27438 3349
rect 27404 3247 27438 3281
rect 27404 3179 27438 3213
rect 27404 3111 27438 3145
rect 27404 3043 27438 3077
rect 27404 2975 27438 3009
rect 27404 2907 27438 2941
rect 27404 2839 27438 2873
rect 27404 2771 27438 2805
rect 27404 2703 27438 2737
rect 27404 2635 27438 2669
rect 27404 2567 27438 2601
rect 27500 3451 27534 3485
rect 27500 3383 27534 3417
rect 27500 3315 27534 3349
rect 27500 3247 27534 3281
rect 27500 3179 27534 3213
rect 27500 3111 27534 3145
rect 27500 3043 27534 3077
rect 27500 2975 27534 3009
rect 27500 2907 27534 2941
rect 27500 2839 27534 2873
rect 27500 2771 27534 2805
rect 27500 2703 27534 2737
rect 27500 2635 27534 2669
rect 27500 2567 27534 2601
rect 27596 3451 27630 3485
rect 27596 3383 27630 3417
rect 27596 3315 27630 3349
rect 27596 3247 27630 3281
rect 27596 3179 27630 3213
rect 27596 3111 27630 3145
rect 27596 3043 27630 3077
rect 27596 2975 27630 3009
rect 27596 2907 27630 2941
rect 27596 2839 27630 2873
rect 27596 2771 27630 2805
rect 27596 2703 27630 2737
rect 27596 2635 27630 2669
rect 27596 2567 27630 2601
rect 27692 3451 27726 3485
rect 27692 3383 27726 3417
rect 27692 3315 27726 3349
rect 27692 3247 27726 3281
rect 27692 3179 27726 3213
rect 27692 3111 27726 3145
rect 27692 3043 27726 3077
rect 27692 2975 27726 3009
rect 27692 2907 27726 2941
rect 27692 2839 27726 2873
rect 27692 2771 27726 2805
rect 27692 2703 27726 2737
rect 27692 2635 27726 2669
rect 27692 2567 27726 2601
rect 27788 3451 27822 3485
rect 27788 3383 27822 3417
rect 27788 3315 27822 3349
rect 27788 3247 27822 3281
rect 27788 3179 27822 3213
rect 27788 3111 27822 3145
rect 27788 3043 27822 3077
rect 27788 2975 27822 3009
rect 27788 2907 27822 2941
rect 27788 2839 27822 2873
rect 27788 2771 27822 2805
rect 27788 2703 27822 2737
rect 27788 2635 27822 2669
rect 27788 2567 27822 2601
rect 27884 3451 27918 3485
rect 27884 3383 27918 3417
rect 27884 3315 27918 3349
rect 27884 3247 27918 3281
rect 27884 3179 27918 3213
rect 27884 3111 27918 3145
rect 27884 3043 27918 3077
rect 27884 2975 27918 3009
rect 27884 2907 27918 2941
rect 27884 2839 27918 2873
rect 27884 2771 27918 2805
rect 27884 2703 27918 2737
rect 27884 2635 27918 2669
rect 27884 2567 27918 2601
rect 27980 3451 28014 3485
rect 27980 3383 28014 3417
rect 27980 3315 28014 3349
rect 27980 3247 28014 3281
rect 27980 3179 28014 3213
rect 27980 3111 28014 3145
rect 27980 3043 28014 3077
rect 27980 2975 28014 3009
rect 27980 2907 28014 2941
rect 27980 2839 28014 2873
rect 27980 2771 28014 2805
rect 27980 2703 28014 2737
rect 27980 2635 28014 2669
rect 27980 2567 28014 2601
rect 28076 3451 28110 3485
rect 28076 3383 28110 3417
rect 28076 3315 28110 3349
rect 28076 3247 28110 3281
rect 28076 3179 28110 3213
rect 28076 3111 28110 3145
rect 28076 3043 28110 3077
rect 28076 2975 28110 3009
rect 28076 2907 28110 2941
rect 28076 2839 28110 2873
rect 28076 2771 28110 2805
rect 28076 2703 28110 2737
rect 28076 2635 28110 2669
rect 28076 2567 28110 2601
rect 28172 3451 28206 3485
rect 28172 3383 28206 3417
rect 28172 3315 28206 3349
rect 28172 3247 28206 3281
rect 28172 3179 28206 3213
rect 28172 3111 28206 3145
rect 28172 3043 28206 3077
rect 28172 2975 28206 3009
rect 28172 2907 28206 2941
rect 28172 2839 28206 2873
rect 28172 2771 28206 2805
rect 28172 2703 28206 2737
rect 28172 2635 28206 2669
rect 28172 2567 28206 2601
rect 28268 3451 28302 3485
rect 28268 3383 28302 3417
rect 28268 3315 28302 3349
rect 28268 3247 28302 3281
rect 28268 3179 28302 3213
rect 28268 3111 28302 3145
rect 28268 3043 28302 3077
rect 28268 2975 28302 3009
rect 28268 2907 28302 2941
rect 28268 2839 28302 2873
rect 28268 2771 28302 2805
rect 28268 2703 28302 2737
rect 28268 2635 28302 2669
rect 28268 2567 28302 2601
rect 28364 3451 28398 3485
rect 28364 3383 28398 3417
rect 28364 3315 28398 3349
rect 28364 3247 28398 3281
rect 28364 3179 28398 3213
rect 28364 3111 28398 3145
rect 28364 3043 28398 3077
rect 28364 2975 28398 3009
rect 28364 2907 28398 2941
rect 28364 2839 28398 2873
rect 28364 2771 28398 2805
rect 28364 2703 28398 2737
rect 28364 2635 28398 2669
rect 28364 2567 28398 2601
rect 28460 3451 28494 3485
rect 28460 3383 28494 3417
rect 28460 3315 28494 3349
rect 28460 3247 28494 3281
rect 28460 3179 28494 3213
rect 28460 3111 28494 3145
rect 28460 3043 28494 3077
rect 28460 2975 28494 3009
rect 28460 2907 28494 2941
rect 28460 2839 28494 2873
rect 28460 2771 28494 2805
rect 28460 2703 28494 2737
rect 28460 2635 28494 2669
rect 28460 2567 28494 2601
rect 28556 3451 28590 3485
rect 28556 3383 28590 3417
rect 28556 3315 28590 3349
rect 28556 3247 28590 3281
rect 28556 3179 28590 3213
rect 28556 3111 28590 3145
rect 28556 3043 28590 3077
rect 28556 2975 28590 3009
rect 28556 2907 28590 2941
rect 28556 2839 28590 2873
rect 28556 2771 28590 2805
rect 28556 2703 28590 2737
rect 28556 2635 28590 2669
rect 28556 2567 28590 2601
rect 28652 3451 28686 3485
rect 28652 3383 28686 3417
rect 28652 3315 28686 3349
rect 28652 3247 28686 3281
rect 28652 3179 28686 3213
rect 28652 3111 28686 3145
rect 28652 3043 28686 3077
rect 28652 2975 28686 3009
rect 28652 2907 28686 2941
rect 28652 2839 28686 2873
rect 28652 2771 28686 2805
rect 28652 2703 28686 2737
rect 28652 2635 28686 2669
rect 28652 2567 28686 2601
rect 14096 2439 14130 2473
rect 14096 2371 14130 2405
rect 14096 2303 14130 2337
rect 14096 2235 14130 2269
rect 14096 2167 14130 2201
rect 14096 2099 14130 2133
rect 14500 2227 14534 2261
rect 14500 2159 14534 2193
rect 14500 2091 14534 2125
rect 14658 2227 14692 2261
rect 14658 2159 14692 2193
rect 14658 2091 14692 2125
rect 14096 2031 14130 2065
rect 14096 1963 14130 1997
rect 14096 1895 14130 1929
rect 14096 1827 14130 1861
rect 158 1193 192 1227
rect 158 1125 192 1159
rect -1686 991 -1652 1025
rect -1686 923 -1652 957
rect -1686 855 -1652 889
rect -1686 787 -1652 821
rect -1686 719 -1652 753
rect -1686 651 -1652 685
rect -1686 583 -1652 617
rect -1686 515 -1652 549
rect -1686 447 -1652 481
rect -1686 379 -1652 413
rect -1686 311 -1652 345
rect -1686 243 -1652 277
rect -1686 175 -1652 209
rect -1686 107 -1652 141
rect -1588 991 -1554 1025
rect -1588 923 -1554 957
rect -1588 855 -1554 889
rect -1588 787 -1554 821
rect -1588 719 -1554 753
rect -1588 651 -1554 685
rect -1588 583 -1554 617
rect -1588 515 -1554 549
rect -1588 447 -1554 481
rect -1588 379 -1554 413
rect -1588 311 -1554 345
rect -1588 243 -1554 277
rect -1588 175 -1554 209
rect -1588 107 -1554 141
rect -1490 991 -1456 1025
rect -1490 923 -1456 957
rect -1490 855 -1456 889
rect -1490 787 -1456 821
rect -1490 719 -1456 753
rect -1490 651 -1456 685
rect -1490 583 -1456 617
rect -1490 515 -1456 549
rect -1490 447 -1456 481
rect -1490 379 -1456 413
rect -1490 311 -1456 345
rect -1490 243 -1456 277
rect -1490 175 -1456 209
rect -1490 107 -1456 141
rect -1392 991 -1358 1025
rect -1392 923 -1358 957
rect -1392 855 -1358 889
rect -1392 787 -1358 821
rect -1392 719 -1358 753
rect -1392 651 -1358 685
rect -1392 583 -1358 617
rect -1392 515 -1358 549
rect -1392 447 -1358 481
rect -1392 379 -1358 413
rect -1392 311 -1358 345
rect -1392 243 -1358 277
rect -1392 175 -1358 209
rect -1392 107 -1358 141
rect -1294 991 -1260 1025
rect -1294 923 -1260 957
rect -1294 855 -1260 889
rect -1294 787 -1260 821
rect -1294 719 -1260 753
rect -1294 651 -1260 685
rect -1294 583 -1260 617
rect -1294 515 -1260 549
rect -1294 447 -1260 481
rect -1294 379 -1260 413
rect -1294 311 -1260 345
rect -1294 243 -1260 277
rect -1294 175 -1260 209
rect -1294 107 -1260 141
rect -1196 991 -1162 1025
rect -1196 923 -1162 957
rect -1196 855 -1162 889
rect -1196 787 -1162 821
rect -1196 719 -1162 753
rect -1196 651 -1162 685
rect -1196 583 -1162 617
rect -1196 515 -1162 549
rect -1196 447 -1162 481
rect -1196 379 -1162 413
rect -1196 311 -1162 345
rect -1196 243 -1162 277
rect -1196 175 -1162 209
rect -1196 107 -1162 141
rect -1098 991 -1064 1025
rect -1098 923 -1064 957
rect -1098 855 -1064 889
rect -1098 787 -1064 821
rect -1098 719 -1064 753
rect -1098 651 -1064 685
rect -1098 583 -1064 617
rect -1098 515 -1064 549
rect -1098 447 -1064 481
rect -1098 379 -1064 413
rect -1098 311 -1064 345
rect -1098 243 -1064 277
rect -1098 175 -1064 209
rect -1098 107 -1064 141
rect -1000 991 -966 1025
rect -1000 923 -966 957
rect -1000 855 -966 889
rect -1000 787 -966 821
rect -1000 719 -966 753
rect -1000 651 -966 685
rect -1000 583 -966 617
rect -1000 515 -966 549
rect -1000 447 -966 481
rect -1000 379 -966 413
rect -1000 311 -966 345
rect -1000 243 -966 277
rect -1000 175 -966 209
rect -1000 107 -966 141
rect -902 991 -868 1025
rect -902 923 -868 957
rect -902 855 -868 889
rect -902 787 -868 821
rect -902 719 -868 753
rect -902 651 -868 685
rect -902 583 -868 617
rect -902 515 -868 549
rect -902 447 -868 481
rect -902 379 -868 413
rect -902 311 -868 345
rect -902 243 -868 277
rect 158 1057 192 1091
rect 158 989 192 1023
rect 158 921 192 955
rect 158 853 192 887
rect 158 785 192 819
rect 158 717 192 751
rect 158 649 192 683
rect 158 581 192 615
rect 158 513 192 547
rect 158 445 192 479
rect 158 377 192 411
rect 158 309 192 343
rect 254 1193 288 1227
rect 254 1125 288 1159
rect 254 1057 288 1091
rect 254 989 288 1023
rect 254 921 288 955
rect 254 853 288 887
rect 254 785 288 819
rect 254 717 288 751
rect 254 649 288 683
rect 254 581 288 615
rect 254 513 288 547
rect 254 445 288 479
rect 254 377 288 411
rect 254 309 288 343
rect 350 1193 384 1227
rect 350 1125 384 1159
rect 350 1057 384 1091
rect 350 989 384 1023
rect 350 921 384 955
rect 350 853 384 887
rect 350 785 384 819
rect 350 717 384 751
rect 350 649 384 683
rect 350 581 384 615
rect 350 513 384 547
rect 350 445 384 479
rect 350 377 384 411
rect 350 309 384 343
rect 446 1193 480 1227
rect 446 1125 480 1159
rect 446 1057 480 1091
rect 446 989 480 1023
rect 446 921 480 955
rect 446 853 480 887
rect 446 785 480 819
rect 446 717 480 751
rect 446 649 480 683
rect 446 581 480 615
rect 446 513 480 547
rect 446 445 480 479
rect 446 377 480 411
rect 446 309 480 343
rect 542 1193 576 1227
rect 542 1125 576 1159
rect 542 1057 576 1091
rect 542 989 576 1023
rect 542 921 576 955
rect 542 853 576 887
rect 542 785 576 819
rect 542 717 576 751
rect 542 649 576 683
rect 542 581 576 615
rect 542 513 576 547
rect 542 445 576 479
rect 542 377 576 411
rect 542 309 576 343
rect 638 1193 672 1227
rect 638 1125 672 1159
rect 638 1057 672 1091
rect 638 989 672 1023
rect 638 921 672 955
rect 638 853 672 887
rect 638 785 672 819
rect 638 717 672 751
rect 638 649 672 683
rect 638 581 672 615
rect 638 513 672 547
rect 638 445 672 479
rect 638 377 672 411
rect 638 309 672 343
rect 734 1193 768 1227
rect 734 1125 768 1159
rect 734 1057 768 1091
rect 734 989 768 1023
rect 734 921 768 955
rect 734 853 768 887
rect 734 785 768 819
rect 734 717 768 751
rect 734 649 768 683
rect 734 581 768 615
rect 734 513 768 547
rect 734 445 768 479
rect 734 377 768 411
rect 734 309 768 343
rect 830 1193 864 1227
rect 830 1125 864 1159
rect 830 1057 864 1091
rect 830 989 864 1023
rect 830 921 864 955
rect 830 853 864 887
rect 830 785 864 819
rect 830 717 864 751
rect 830 649 864 683
rect 830 581 864 615
rect 830 513 864 547
rect 830 445 864 479
rect 830 377 864 411
rect 830 309 864 343
rect 926 1193 960 1227
rect 926 1125 960 1159
rect 926 1057 960 1091
rect 926 989 960 1023
rect 926 921 960 955
rect 926 853 960 887
rect 926 785 960 819
rect 926 717 960 751
rect 926 649 960 683
rect 926 581 960 615
rect 926 513 960 547
rect 926 445 960 479
rect 926 377 960 411
rect 926 309 960 343
rect 1022 1193 1056 1227
rect 1022 1125 1056 1159
rect 1022 1057 1056 1091
rect 1022 989 1056 1023
rect 1022 921 1056 955
rect 1022 853 1056 887
rect 1022 785 1056 819
rect 1022 717 1056 751
rect 1022 649 1056 683
rect 1022 581 1056 615
rect 1022 513 1056 547
rect 1022 445 1056 479
rect 1022 377 1056 411
rect 1022 309 1056 343
rect 1118 1193 1152 1227
rect 1118 1125 1152 1159
rect 1118 1057 1152 1091
rect 1118 989 1152 1023
rect 1118 921 1152 955
rect 1118 853 1152 887
rect 1118 785 1152 819
rect 1118 717 1152 751
rect 1118 649 1152 683
rect 1118 581 1152 615
rect 1118 513 1152 547
rect 1118 445 1152 479
rect 1118 377 1152 411
rect 1118 309 1152 343
rect 1214 1193 1248 1227
rect 1214 1125 1248 1159
rect 1214 1057 1248 1091
rect 1214 989 1248 1023
rect 1214 921 1248 955
rect 1214 853 1248 887
rect 1214 785 1248 819
rect 1214 717 1248 751
rect 1214 649 1248 683
rect 1214 581 1248 615
rect 1214 513 1248 547
rect 1214 445 1248 479
rect 1214 377 1248 411
rect 1214 309 1248 343
rect 1310 1193 1344 1227
rect 1310 1125 1344 1159
rect 1310 1057 1344 1091
rect 1310 989 1344 1023
rect 1310 921 1344 955
rect 1310 853 1344 887
rect 1310 785 1344 819
rect 1310 717 1344 751
rect 1310 649 1344 683
rect 1310 581 1344 615
rect 1310 513 1344 547
rect 1310 445 1344 479
rect 1310 377 1344 411
rect 1310 309 1344 343
rect 1926 1193 1960 1227
rect 1926 1125 1960 1159
rect 1926 1057 1960 1091
rect 1926 989 1960 1023
rect 1926 921 1960 955
rect 1926 853 1960 887
rect 1926 785 1960 819
rect 1926 717 1960 751
rect 1926 649 1960 683
rect 1926 581 1960 615
rect 1926 513 1960 547
rect 1926 445 1960 479
rect 1926 377 1960 411
rect 1926 309 1960 343
rect 2022 1193 2056 1227
rect 2022 1125 2056 1159
rect 2022 1057 2056 1091
rect 2022 989 2056 1023
rect 2022 921 2056 955
rect 2022 853 2056 887
rect 2022 785 2056 819
rect 2022 717 2056 751
rect 2022 649 2056 683
rect 2022 581 2056 615
rect 2022 513 2056 547
rect 2022 445 2056 479
rect 2022 377 2056 411
rect 2022 309 2056 343
rect 2118 1193 2152 1227
rect 2118 1125 2152 1159
rect 2118 1057 2152 1091
rect 2118 989 2152 1023
rect 2118 921 2152 955
rect 2118 853 2152 887
rect 2118 785 2152 819
rect 2118 717 2152 751
rect 2118 649 2152 683
rect 2118 581 2152 615
rect 2118 513 2152 547
rect 2118 445 2152 479
rect 2118 377 2152 411
rect 2118 309 2152 343
rect 2214 1193 2248 1227
rect 2214 1125 2248 1159
rect 2214 1057 2248 1091
rect 2214 989 2248 1023
rect 2214 921 2248 955
rect 2214 853 2248 887
rect 2214 785 2248 819
rect 2214 717 2248 751
rect 2214 649 2248 683
rect 2214 581 2248 615
rect 2214 513 2248 547
rect 2214 445 2248 479
rect 2214 377 2248 411
rect 2214 309 2248 343
rect 2310 1193 2344 1227
rect 2310 1125 2344 1159
rect 2310 1057 2344 1091
rect 2310 989 2344 1023
rect 2310 921 2344 955
rect 2310 853 2344 887
rect 2310 785 2344 819
rect 2310 717 2344 751
rect 2310 649 2344 683
rect 2310 581 2344 615
rect 2310 513 2344 547
rect 2310 445 2344 479
rect 2310 377 2344 411
rect 2310 309 2344 343
rect 2406 1193 2440 1227
rect 2406 1125 2440 1159
rect 2406 1057 2440 1091
rect 2406 989 2440 1023
rect 2406 921 2440 955
rect 2406 853 2440 887
rect 2406 785 2440 819
rect 2406 717 2440 751
rect 2406 649 2440 683
rect 2406 581 2440 615
rect 2406 513 2440 547
rect 2406 445 2440 479
rect 2406 377 2440 411
rect 2406 309 2440 343
rect 2502 1193 2536 1227
rect 2502 1125 2536 1159
rect 2502 1057 2536 1091
rect 2502 989 2536 1023
rect 2502 921 2536 955
rect 2502 853 2536 887
rect 2502 785 2536 819
rect 2502 717 2536 751
rect 2502 649 2536 683
rect 2502 581 2536 615
rect 2502 513 2536 547
rect 2502 445 2536 479
rect 2502 377 2536 411
rect 2502 309 2536 343
rect 2598 1193 2632 1227
rect 2598 1125 2632 1159
rect 2598 1057 2632 1091
rect 2598 989 2632 1023
rect 2598 921 2632 955
rect 2598 853 2632 887
rect 2598 785 2632 819
rect 2598 717 2632 751
rect 2598 649 2632 683
rect 2598 581 2632 615
rect 2598 513 2632 547
rect 2598 445 2632 479
rect 2598 377 2632 411
rect 2598 309 2632 343
rect 2694 1193 2728 1227
rect 2694 1125 2728 1159
rect 2694 1057 2728 1091
rect 2694 989 2728 1023
rect 2694 921 2728 955
rect 2694 853 2728 887
rect 2694 785 2728 819
rect 2694 717 2728 751
rect 2694 649 2728 683
rect 2694 581 2728 615
rect 2694 513 2728 547
rect 2694 445 2728 479
rect 2694 377 2728 411
rect 2694 309 2728 343
rect 2790 1193 2824 1227
rect 2790 1125 2824 1159
rect 2790 1057 2824 1091
rect 2790 989 2824 1023
rect 2790 921 2824 955
rect 2790 853 2824 887
rect 2790 785 2824 819
rect 2790 717 2824 751
rect 2790 649 2824 683
rect 2790 581 2824 615
rect 2790 513 2824 547
rect 2790 445 2824 479
rect 2790 377 2824 411
rect 2790 309 2824 343
rect 2886 1193 2920 1227
rect 2886 1125 2920 1159
rect 2886 1057 2920 1091
rect 2886 989 2920 1023
rect 2886 921 2920 955
rect 2886 853 2920 887
rect 2886 785 2920 819
rect 2886 717 2920 751
rect 2886 649 2920 683
rect 2886 581 2920 615
rect 2886 513 2920 547
rect 2886 445 2920 479
rect 2886 377 2920 411
rect 2886 309 2920 343
rect 2982 1193 3016 1227
rect 2982 1125 3016 1159
rect 2982 1057 3016 1091
rect 2982 989 3016 1023
rect 2982 921 3016 955
rect 2982 853 3016 887
rect 2982 785 3016 819
rect 2982 717 3016 751
rect 2982 649 3016 683
rect 2982 581 3016 615
rect 2982 513 3016 547
rect 2982 445 3016 479
rect 2982 377 3016 411
rect 2982 309 3016 343
rect 3114 1177 3148 1211
rect 3114 1109 3148 1143
rect 3114 1041 3148 1075
rect 3114 973 3148 1007
rect 3114 905 3148 939
rect 3114 837 3148 871
rect 3114 769 3148 803
rect 3114 701 3148 735
rect 3114 633 3148 667
rect 3114 565 3148 599
rect 3114 497 3148 531
rect 3114 429 3148 463
rect 3114 361 3148 395
rect 3114 293 3148 327
rect -902 175 -868 209
rect 3210 1177 3244 1211
rect 3210 1109 3244 1143
rect 3210 1041 3244 1075
rect 3210 973 3244 1007
rect 3210 905 3244 939
rect 3210 837 3244 871
rect 3210 769 3244 803
rect 3210 701 3244 735
rect 3210 633 3244 667
rect 3210 565 3244 599
rect 3210 497 3244 531
rect 3210 429 3244 463
rect 3210 361 3244 395
rect 3210 293 3244 327
rect 3306 1177 3340 1211
rect 3306 1109 3340 1143
rect 3306 1041 3340 1075
rect 3306 973 3340 1007
rect 3306 905 3340 939
rect 3306 837 3340 871
rect 3306 769 3340 803
rect 3306 701 3340 735
rect 3306 633 3340 667
rect 3306 565 3340 599
rect 3306 497 3340 531
rect 3306 429 3340 463
rect 3306 361 3340 395
rect 3306 293 3340 327
rect 3402 1177 3436 1211
rect 3402 1109 3436 1143
rect 3402 1041 3436 1075
rect 3402 973 3436 1007
rect 3402 905 3436 939
rect 3402 837 3436 871
rect 3402 769 3436 803
rect 3402 701 3436 735
rect 3402 633 3436 667
rect 3402 565 3436 599
rect 3402 497 3436 531
rect 3402 429 3436 463
rect 3402 361 3436 395
rect 3402 293 3436 327
rect 3498 1177 3532 1211
rect 3498 1109 3532 1143
rect 3498 1041 3532 1075
rect 3498 973 3532 1007
rect 3498 905 3532 939
rect 3498 837 3532 871
rect 3498 769 3532 803
rect 3498 701 3532 735
rect 3498 633 3532 667
rect 3498 565 3532 599
rect 3498 497 3532 531
rect 3498 429 3532 463
rect 3498 361 3532 395
rect 3498 293 3532 327
rect 3594 1177 3628 1211
rect 3594 1109 3628 1143
rect 3594 1041 3628 1075
rect 3594 973 3628 1007
rect 3594 905 3628 939
rect 3594 837 3628 871
rect 3594 769 3628 803
rect 3594 701 3628 735
rect 3594 633 3628 667
rect 3594 565 3628 599
rect 3594 497 3628 531
rect 3594 429 3628 463
rect 3594 361 3628 395
rect 3594 293 3628 327
rect 3690 1177 3724 1211
rect 3690 1109 3724 1143
rect 3690 1041 3724 1075
rect 3690 973 3724 1007
rect 3690 905 3724 939
rect 3690 837 3724 871
rect 3690 769 3724 803
rect 3690 701 3724 735
rect 3690 633 3724 667
rect 3690 565 3724 599
rect 3690 497 3724 531
rect 3690 429 3724 463
rect 3690 361 3724 395
rect 3690 293 3724 327
rect 3786 1177 3820 1211
rect 3786 1109 3820 1143
rect 3786 1041 3820 1075
rect 3786 973 3820 1007
rect 3786 905 3820 939
rect 3786 837 3820 871
rect 3786 769 3820 803
rect 3786 701 3820 735
rect 3786 633 3820 667
rect 3786 565 3820 599
rect 3786 497 3820 531
rect 3786 429 3820 463
rect 3786 361 3820 395
rect 3786 293 3820 327
rect 3882 1177 3916 1211
rect 3882 1109 3916 1143
rect 3882 1041 3916 1075
rect 3882 973 3916 1007
rect 3882 905 3916 939
rect 3882 837 3916 871
rect 3882 769 3916 803
rect 3882 701 3916 735
rect 3882 633 3916 667
rect 3882 565 3916 599
rect 3882 497 3916 531
rect 3882 429 3916 463
rect 3882 361 3916 395
rect 3882 293 3916 327
rect 3978 1177 4012 1211
rect 3978 1109 4012 1143
rect 3978 1041 4012 1075
rect 3978 973 4012 1007
rect 3978 905 4012 939
rect 3978 837 4012 871
rect 3978 769 4012 803
rect 3978 701 4012 735
rect 3978 633 4012 667
rect 3978 565 4012 599
rect 3978 497 4012 531
rect 3978 429 4012 463
rect 3978 361 4012 395
rect 3978 293 4012 327
rect 4074 1177 4108 1211
rect 4074 1109 4108 1143
rect 4074 1041 4108 1075
rect 4074 973 4108 1007
rect 4074 905 4108 939
rect 4074 837 4108 871
rect 4074 769 4108 803
rect 4074 701 4108 735
rect 4074 633 4108 667
rect 4074 565 4108 599
rect 4074 497 4108 531
rect 4074 429 4108 463
rect 4074 361 4108 395
rect 4074 293 4108 327
rect 4170 1177 4204 1211
rect 4170 1109 4204 1143
rect 4170 1041 4204 1075
rect 4170 973 4204 1007
rect 4170 905 4204 939
rect 4170 837 4204 871
rect 4170 769 4204 803
rect 4170 701 4204 735
rect 4170 633 4204 667
rect 4170 565 4204 599
rect 4170 497 4204 531
rect 4170 429 4204 463
rect 4170 361 4204 395
rect 4170 293 4204 327
rect 4266 1177 4300 1211
rect 4266 1109 4300 1143
rect 4266 1041 4300 1075
rect 4266 973 4300 1007
rect 4266 905 4300 939
rect 4266 837 4300 871
rect 4266 769 4300 803
rect 4266 701 4300 735
rect 4266 633 4300 667
rect 4266 565 4300 599
rect 4266 497 4300 531
rect 4266 429 4300 463
rect 4266 361 4300 395
rect 4266 293 4300 327
rect 4882 1177 4916 1211
rect 4882 1109 4916 1143
rect 4882 1041 4916 1075
rect 4882 973 4916 1007
rect 4882 905 4916 939
rect 4882 837 4916 871
rect 4882 769 4916 803
rect 4882 701 4916 735
rect 4882 633 4916 667
rect 4882 565 4916 599
rect 4882 497 4916 531
rect 4882 429 4916 463
rect 4882 361 4916 395
rect 4882 293 4916 327
rect 4978 1177 5012 1211
rect 4978 1109 5012 1143
rect 4978 1041 5012 1075
rect 4978 973 5012 1007
rect 4978 905 5012 939
rect 4978 837 5012 871
rect 4978 769 5012 803
rect 4978 701 5012 735
rect 4978 633 5012 667
rect 4978 565 5012 599
rect 4978 497 5012 531
rect 4978 429 5012 463
rect 4978 361 5012 395
rect 4978 293 5012 327
rect 5074 1177 5108 1211
rect 5074 1109 5108 1143
rect 5074 1041 5108 1075
rect 5074 973 5108 1007
rect 5074 905 5108 939
rect 5074 837 5108 871
rect 5074 769 5108 803
rect 5074 701 5108 735
rect 5074 633 5108 667
rect 5074 565 5108 599
rect 5074 497 5108 531
rect 5074 429 5108 463
rect 5074 361 5108 395
rect 5074 293 5108 327
rect 5170 1177 5204 1211
rect 5170 1109 5204 1143
rect 5170 1041 5204 1075
rect 5170 973 5204 1007
rect 5170 905 5204 939
rect 5170 837 5204 871
rect 5170 769 5204 803
rect 5170 701 5204 735
rect 5170 633 5204 667
rect 5170 565 5204 599
rect 5170 497 5204 531
rect 5170 429 5204 463
rect 5170 361 5204 395
rect 5170 293 5204 327
rect 5266 1177 5300 1211
rect 5266 1109 5300 1143
rect 5266 1041 5300 1075
rect 5266 973 5300 1007
rect 5266 905 5300 939
rect 5266 837 5300 871
rect 5266 769 5300 803
rect 5266 701 5300 735
rect 5266 633 5300 667
rect 5266 565 5300 599
rect 5266 497 5300 531
rect 5266 429 5300 463
rect 5266 361 5300 395
rect 5266 293 5300 327
rect 5362 1177 5396 1211
rect 5362 1109 5396 1143
rect 5362 1041 5396 1075
rect 5362 973 5396 1007
rect 5362 905 5396 939
rect 5362 837 5396 871
rect 5362 769 5396 803
rect 5362 701 5396 735
rect 5362 633 5396 667
rect 5362 565 5396 599
rect 5362 497 5396 531
rect 5362 429 5396 463
rect 5362 361 5396 395
rect 5362 293 5396 327
rect 5458 1177 5492 1211
rect 5458 1109 5492 1143
rect 5458 1041 5492 1075
rect 5458 973 5492 1007
rect 5458 905 5492 939
rect 5458 837 5492 871
rect 5458 769 5492 803
rect 5458 701 5492 735
rect 5458 633 5492 667
rect 5458 565 5492 599
rect 5458 497 5492 531
rect 5458 429 5492 463
rect 5458 361 5492 395
rect 5458 293 5492 327
rect 5554 1177 5588 1211
rect 5554 1109 5588 1143
rect 5554 1041 5588 1075
rect 5554 973 5588 1007
rect 5554 905 5588 939
rect 5554 837 5588 871
rect 5554 769 5588 803
rect 5554 701 5588 735
rect 5554 633 5588 667
rect 5554 565 5588 599
rect 5554 497 5588 531
rect 5554 429 5588 463
rect 5554 361 5588 395
rect 5554 293 5588 327
rect 5650 1177 5684 1211
rect 5650 1109 5684 1143
rect 5650 1041 5684 1075
rect 5650 973 5684 1007
rect 5650 905 5684 939
rect 5650 837 5684 871
rect 5650 769 5684 803
rect 5650 701 5684 735
rect 5650 633 5684 667
rect 5650 565 5684 599
rect 5650 497 5684 531
rect 5650 429 5684 463
rect 5650 361 5684 395
rect 5650 293 5684 327
rect 5746 1177 5780 1211
rect 5746 1109 5780 1143
rect 5746 1041 5780 1075
rect 5746 973 5780 1007
rect 5746 905 5780 939
rect 5746 837 5780 871
rect 5746 769 5780 803
rect 5746 701 5780 735
rect 5746 633 5780 667
rect 5746 565 5780 599
rect 5746 497 5780 531
rect 5746 429 5780 463
rect 5746 361 5780 395
rect 5746 293 5780 327
rect 5842 1177 5876 1211
rect 5842 1109 5876 1143
rect 5842 1041 5876 1075
rect 5842 973 5876 1007
rect 5842 905 5876 939
rect 5842 837 5876 871
rect 5842 769 5876 803
rect 5842 701 5876 735
rect 5842 633 5876 667
rect 5842 565 5876 599
rect 5842 497 5876 531
rect 5842 429 5876 463
rect 5842 361 5876 395
rect 5842 293 5876 327
rect 5938 1177 5972 1211
rect 5938 1109 5972 1143
rect 5938 1041 5972 1075
rect 5938 973 5972 1007
rect 5938 905 5972 939
rect 5938 837 5972 871
rect 5938 769 5972 803
rect 5938 701 5972 735
rect 5938 633 5972 667
rect 5938 565 5972 599
rect 5938 497 5972 531
rect 5938 429 5972 463
rect 5938 361 5972 395
rect 5938 293 5972 327
rect 6144 1177 6178 1211
rect 6144 1109 6178 1143
rect 6144 1041 6178 1075
rect 6144 973 6178 1007
rect 6144 905 6178 939
rect 6144 837 6178 871
rect 6144 769 6178 803
rect 6144 701 6178 735
rect 6144 633 6178 667
rect 6144 565 6178 599
rect 6144 497 6178 531
rect 6144 429 6178 463
rect 6144 361 6178 395
rect 6144 293 6178 327
rect 6240 1177 6274 1211
rect 6240 1109 6274 1143
rect 6240 1041 6274 1075
rect 6240 973 6274 1007
rect 6240 905 6274 939
rect 6240 837 6274 871
rect 6240 769 6274 803
rect 6240 701 6274 735
rect 6240 633 6274 667
rect 6240 565 6274 599
rect 6240 497 6274 531
rect 6240 429 6274 463
rect 6240 361 6274 395
rect 6240 293 6274 327
rect 6336 1177 6370 1211
rect 6336 1109 6370 1143
rect 6336 1041 6370 1075
rect 6336 973 6370 1007
rect 6336 905 6370 939
rect 6336 837 6370 871
rect 6336 769 6370 803
rect 6336 701 6370 735
rect 6336 633 6370 667
rect 6336 565 6370 599
rect 6336 497 6370 531
rect 6336 429 6370 463
rect 6336 361 6370 395
rect 6336 293 6370 327
rect 6432 1177 6466 1211
rect 6432 1109 6466 1143
rect 6432 1041 6466 1075
rect 6432 973 6466 1007
rect 6432 905 6466 939
rect 6432 837 6466 871
rect 6432 769 6466 803
rect 6432 701 6466 735
rect 6432 633 6466 667
rect 6432 565 6466 599
rect 6432 497 6466 531
rect 6432 429 6466 463
rect 6432 361 6466 395
rect 6432 293 6466 327
rect 6528 1177 6562 1211
rect 6528 1109 6562 1143
rect 6528 1041 6562 1075
rect 6528 973 6562 1007
rect 6528 905 6562 939
rect 6528 837 6562 871
rect 6528 769 6562 803
rect 6528 701 6562 735
rect 6528 633 6562 667
rect 6528 565 6562 599
rect 6528 497 6562 531
rect 6528 429 6562 463
rect 6528 361 6562 395
rect 6528 293 6562 327
rect 6624 1177 6658 1211
rect 6624 1109 6658 1143
rect 6624 1041 6658 1075
rect 6624 973 6658 1007
rect 6624 905 6658 939
rect 6624 837 6658 871
rect 6624 769 6658 803
rect 6624 701 6658 735
rect 6624 633 6658 667
rect 6624 565 6658 599
rect 6624 497 6658 531
rect 6624 429 6658 463
rect 6624 361 6658 395
rect 6624 293 6658 327
rect 6720 1177 6754 1211
rect 6720 1109 6754 1143
rect 6720 1041 6754 1075
rect 6720 973 6754 1007
rect 6720 905 6754 939
rect 6720 837 6754 871
rect 6720 769 6754 803
rect 6720 701 6754 735
rect 6720 633 6754 667
rect 6720 565 6754 599
rect 6720 497 6754 531
rect 6720 429 6754 463
rect 6720 361 6754 395
rect 6720 293 6754 327
rect 6816 1177 6850 1211
rect 6816 1109 6850 1143
rect 6816 1041 6850 1075
rect 6816 973 6850 1007
rect 6816 905 6850 939
rect 6816 837 6850 871
rect 6816 769 6850 803
rect 6816 701 6850 735
rect 6816 633 6850 667
rect 6816 565 6850 599
rect 6816 497 6850 531
rect 6816 429 6850 463
rect 6816 361 6850 395
rect 6816 293 6850 327
rect 6912 1177 6946 1211
rect 6912 1109 6946 1143
rect 6912 1041 6946 1075
rect 6912 973 6946 1007
rect 6912 905 6946 939
rect 6912 837 6946 871
rect 6912 769 6946 803
rect 6912 701 6946 735
rect 6912 633 6946 667
rect 6912 565 6946 599
rect 6912 497 6946 531
rect 6912 429 6946 463
rect 6912 361 6946 395
rect 6912 293 6946 327
rect 7008 1177 7042 1211
rect 7008 1109 7042 1143
rect 7008 1041 7042 1075
rect 7008 973 7042 1007
rect 7008 905 7042 939
rect 7008 837 7042 871
rect 7008 769 7042 803
rect 7008 701 7042 735
rect 7008 633 7042 667
rect 7008 565 7042 599
rect 7008 497 7042 531
rect 7008 429 7042 463
rect 7008 361 7042 395
rect 7008 293 7042 327
rect 7104 1177 7138 1211
rect 7104 1109 7138 1143
rect 7104 1041 7138 1075
rect 7104 973 7138 1007
rect 7104 905 7138 939
rect 7104 837 7138 871
rect 7104 769 7138 803
rect 7104 701 7138 735
rect 7104 633 7138 667
rect 7104 565 7138 599
rect 7104 497 7138 531
rect 7104 429 7138 463
rect 7104 361 7138 395
rect 7104 293 7138 327
rect 7200 1177 7234 1211
rect 7200 1109 7234 1143
rect 7200 1041 7234 1075
rect 7200 973 7234 1007
rect 7200 905 7234 939
rect 7200 837 7234 871
rect 7200 769 7234 803
rect 7200 701 7234 735
rect 7200 633 7234 667
rect 7200 565 7234 599
rect 7200 497 7234 531
rect 7200 429 7234 463
rect 7200 361 7234 395
rect 7200 293 7234 327
rect 7296 1177 7330 1211
rect 7296 1109 7330 1143
rect 7296 1041 7330 1075
rect 7296 973 7330 1007
rect 7296 905 7330 939
rect 7296 837 7330 871
rect 7296 769 7330 803
rect 7296 701 7330 735
rect 7296 633 7330 667
rect 7296 565 7330 599
rect 7296 497 7330 531
rect 7296 429 7330 463
rect 7296 361 7330 395
rect 7296 293 7330 327
rect 7912 1177 7946 1211
rect 7912 1109 7946 1143
rect 7912 1041 7946 1075
rect 7912 973 7946 1007
rect 7912 905 7946 939
rect 7912 837 7946 871
rect 7912 769 7946 803
rect 7912 701 7946 735
rect 7912 633 7946 667
rect 7912 565 7946 599
rect 7912 497 7946 531
rect 7912 429 7946 463
rect 7912 361 7946 395
rect 7912 293 7946 327
rect 8008 1177 8042 1211
rect 8008 1109 8042 1143
rect 8008 1041 8042 1075
rect 8008 973 8042 1007
rect 8008 905 8042 939
rect 8008 837 8042 871
rect 8008 769 8042 803
rect 8008 701 8042 735
rect 8008 633 8042 667
rect 8008 565 8042 599
rect 8008 497 8042 531
rect 8008 429 8042 463
rect 8008 361 8042 395
rect 8008 293 8042 327
rect 8104 1177 8138 1211
rect 8104 1109 8138 1143
rect 8104 1041 8138 1075
rect 8104 973 8138 1007
rect 8104 905 8138 939
rect 8104 837 8138 871
rect 8104 769 8138 803
rect 8104 701 8138 735
rect 8104 633 8138 667
rect 8104 565 8138 599
rect 8104 497 8138 531
rect 8104 429 8138 463
rect 8104 361 8138 395
rect 8104 293 8138 327
rect 8200 1177 8234 1211
rect 8200 1109 8234 1143
rect 8200 1041 8234 1075
rect 8200 973 8234 1007
rect 8200 905 8234 939
rect 8200 837 8234 871
rect 8200 769 8234 803
rect 8200 701 8234 735
rect 8200 633 8234 667
rect 8200 565 8234 599
rect 8200 497 8234 531
rect 8200 429 8234 463
rect 8200 361 8234 395
rect 8200 293 8234 327
rect 8296 1177 8330 1211
rect 8296 1109 8330 1143
rect 8296 1041 8330 1075
rect 8296 973 8330 1007
rect 8296 905 8330 939
rect 8296 837 8330 871
rect 8296 769 8330 803
rect 8296 701 8330 735
rect 8296 633 8330 667
rect 8296 565 8330 599
rect 8296 497 8330 531
rect 8296 429 8330 463
rect 8296 361 8330 395
rect 8296 293 8330 327
rect 8392 1177 8426 1211
rect 8392 1109 8426 1143
rect 8392 1041 8426 1075
rect 8392 973 8426 1007
rect 8392 905 8426 939
rect 8392 837 8426 871
rect 8392 769 8426 803
rect 8392 701 8426 735
rect 8392 633 8426 667
rect 8392 565 8426 599
rect 8392 497 8426 531
rect 8392 429 8426 463
rect 8392 361 8426 395
rect 8392 293 8426 327
rect 8488 1177 8522 1211
rect 8488 1109 8522 1143
rect 8488 1041 8522 1075
rect 8488 973 8522 1007
rect 8488 905 8522 939
rect 8488 837 8522 871
rect 8488 769 8522 803
rect 8488 701 8522 735
rect 8488 633 8522 667
rect 8488 565 8522 599
rect 8488 497 8522 531
rect 8488 429 8522 463
rect 8488 361 8522 395
rect 8488 293 8522 327
rect 8584 1177 8618 1211
rect 8584 1109 8618 1143
rect 8584 1041 8618 1075
rect 8584 973 8618 1007
rect 8584 905 8618 939
rect 8584 837 8618 871
rect 8584 769 8618 803
rect 8584 701 8618 735
rect 8584 633 8618 667
rect 8584 565 8618 599
rect 8584 497 8618 531
rect 8584 429 8618 463
rect 8584 361 8618 395
rect 8584 293 8618 327
rect 8680 1177 8714 1211
rect 8680 1109 8714 1143
rect 8680 1041 8714 1075
rect 8680 973 8714 1007
rect 8680 905 8714 939
rect 8680 837 8714 871
rect 8680 769 8714 803
rect 8680 701 8714 735
rect 8680 633 8714 667
rect 8680 565 8714 599
rect 8680 497 8714 531
rect 8680 429 8714 463
rect 8680 361 8714 395
rect 8680 293 8714 327
rect 8776 1177 8810 1211
rect 8776 1109 8810 1143
rect 8776 1041 8810 1075
rect 8776 973 8810 1007
rect 8776 905 8810 939
rect 8776 837 8810 871
rect 8776 769 8810 803
rect 8776 701 8810 735
rect 8776 633 8810 667
rect 8776 565 8810 599
rect 8776 497 8810 531
rect 8776 429 8810 463
rect 8776 361 8810 395
rect 8776 293 8810 327
rect 8872 1177 8906 1211
rect 8872 1109 8906 1143
rect 8872 1041 8906 1075
rect 8872 973 8906 1007
rect 8872 905 8906 939
rect 8872 837 8906 871
rect 8872 769 8906 803
rect 8872 701 8906 735
rect 8872 633 8906 667
rect 8872 565 8906 599
rect 8872 497 8906 531
rect 8872 429 8906 463
rect 8872 361 8906 395
rect 8872 293 8906 327
rect 8968 1177 9002 1211
rect 8968 1109 9002 1143
rect 8968 1041 9002 1075
rect 8968 973 9002 1007
rect 8968 905 9002 939
rect 8968 837 9002 871
rect 8968 769 9002 803
rect 8968 701 9002 735
rect 8968 633 9002 667
rect 8968 565 9002 599
rect 8968 497 9002 531
rect 8968 429 9002 463
rect 8968 361 9002 395
rect 8968 293 9002 327
rect 9232 1175 9266 1209
rect 9232 1107 9266 1141
rect 9232 1039 9266 1073
rect 9232 971 9266 1005
rect 9232 903 9266 937
rect 9232 835 9266 869
rect 9232 767 9266 801
rect 9232 699 9266 733
rect 9232 631 9266 665
rect 9232 563 9266 597
rect 9232 495 9266 529
rect 9232 427 9266 461
rect 9232 359 9266 393
rect 9232 291 9266 325
rect -902 107 -868 141
rect 9328 1175 9362 1209
rect 9328 1107 9362 1141
rect 9328 1039 9362 1073
rect 9328 971 9362 1005
rect 9328 903 9362 937
rect 9328 835 9362 869
rect 9328 767 9362 801
rect 9328 699 9362 733
rect 9328 631 9362 665
rect 9328 563 9362 597
rect 9328 495 9362 529
rect 9328 427 9362 461
rect 9328 359 9362 393
rect 9328 291 9362 325
rect 9424 1175 9458 1209
rect 9424 1107 9458 1141
rect 9424 1039 9458 1073
rect 9424 971 9458 1005
rect 9424 903 9458 937
rect 9424 835 9458 869
rect 9424 767 9458 801
rect 9424 699 9458 733
rect 9424 631 9458 665
rect 9424 563 9458 597
rect 9424 495 9458 529
rect 9424 427 9458 461
rect 9424 359 9458 393
rect 9424 291 9458 325
rect 9520 1175 9554 1209
rect 9520 1107 9554 1141
rect 9520 1039 9554 1073
rect 9520 971 9554 1005
rect 9520 903 9554 937
rect 9520 835 9554 869
rect 9520 767 9554 801
rect 9520 699 9554 733
rect 9520 631 9554 665
rect 9520 563 9554 597
rect 9520 495 9554 529
rect 9520 427 9554 461
rect 9520 359 9554 393
rect 9520 291 9554 325
rect 9616 1175 9650 1209
rect 9616 1107 9650 1141
rect 9616 1039 9650 1073
rect 9616 971 9650 1005
rect 9616 903 9650 937
rect 9616 835 9650 869
rect 9616 767 9650 801
rect 9616 699 9650 733
rect 9616 631 9650 665
rect 9616 563 9650 597
rect 9616 495 9650 529
rect 9616 427 9650 461
rect 9616 359 9650 393
rect 9616 291 9650 325
rect 9712 1175 9746 1209
rect 9712 1107 9746 1141
rect 9712 1039 9746 1073
rect 9712 971 9746 1005
rect 9712 903 9746 937
rect 9712 835 9746 869
rect 9712 767 9746 801
rect 9712 699 9746 733
rect 9712 631 9746 665
rect 9712 563 9746 597
rect 9712 495 9746 529
rect 9712 427 9746 461
rect 9712 359 9746 393
rect 9712 291 9746 325
rect 9808 1175 9842 1209
rect 9808 1107 9842 1141
rect 9808 1039 9842 1073
rect 9808 971 9842 1005
rect 9808 903 9842 937
rect 9808 835 9842 869
rect 9808 767 9842 801
rect 9808 699 9842 733
rect 9808 631 9842 665
rect 9808 563 9842 597
rect 9808 495 9842 529
rect 9808 427 9842 461
rect 9808 359 9842 393
rect 9808 291 9842 325
rect 9904 1175 9938 1209
rect 9904 1107 9938 1141
rect 9904 1039 9938 1073
rect 9904 971 9938 1005
rect 9904 903 9938 937
rect 9904 835 9938 869
rect 9904 767 9938 801
rect 9904 699 9938 733
rect 9904 631 9938 665
rect 9904 563 9938 597
rect 9904 495 9938 529
rect 9904 427 9938 461
rect 9904 359 9938 393
rect 9904 291 9938 325
rect 10000 1175 10034 1209
rect 10000 1107 10034 1141
rect 10000 1039 10034 1073
rect 10000 971 10034 1005
rect 10000 903 10034 937
rect 10000 835 10034 869
rect 10000 767 10034 801
rect 10000 699 10034 733
rect 10000 631 10034 665
rect 10000 563 10034 597
rect 10000 495 10034 529
rect 10000 427 10034 461
rect 10000 359 10034 393
rect 10000 291 10034 325
rect 10096 1175 10130 1209
rect 10096 1107 10130 1141
rect 10096 1039 10130 1073
rect 10096 971 10130 1005
rect 10096 903 10130 937
rect 10096 835 10130 869
rect 10096 767 10130 801
rect 10096 699 10130 733
rect 10096 631 10130 665
rect 10096 563 10130 597
rect 10096 495 10130 529
rect 10096 427 10130 461
rect 10096 359 10130 393
rect 10096 291 10130 325
rect 10192 1175 10226 1209
rect 10192 1107 10226 1141
rect 10192 1039 10226 1073
rect 10192 971 10226 1005
rect 10192 903 10226 937
rect 10192 835 10226 869
rect 10192 767 10226 801
rect 10192 699 10226 733
rect 10192 631 10226 665
rect 10192 563 10226 597
rect 10192 495 10226 529
rect 10192 427 10226 461
rect 10192 359 10226 393
rect 10192 291 10226 325
rect 10288 1175 10322 1209
rect 10288 1107 10322 1141
rect 10288 1039 10322 1073
rect 10288 971 10322 1005
rect 10288 903 10322 937
rect 10288 835 10322 869
rect 10288 767 10322 801
rect 10288 699 10322 733
rect 10288 631 10322 665
rect 10288 563 10322 597
rect 10288 495 10322 529
rect 10288 427 10322 461
rect 10288 359 10322 393
rect 10288 291 10322 325
rect 10384 1175 10418 1209
rect 10384 1107 10418 1141
rect 10384 1039 10418 1073
rect 10384 971 10418 1005
rect 10384 903 10418 937
rect 10384 835 10418 869
rect 10384 767 10418 801
rect 10384 699 10418 733
rect 10384 631 10418 665
rect 10384 563 10418 597
rect 10384 495 10418 529
rect 10384 427 10418 461
rect 10384 359 10418 393
rect 10384 291 10418 325
rect 11000 1175 11034 1209
rect 11000 1107 11034 1141
rect 11000 1039 11034 1073
rect 11000 971 11034 1005
rect 11000 903 11034 937
rect 11000 835 11034 869
rect 11000 767 11034 801
rect 11000 699 11034 733
rect 11000 631 11034 665
rect 11000 563 11034 597
rect 11000 495 11034 529
rect 11000 427 11034 461
rect 11000 359 11034 393
rect 11000 291 11034 325
rect 11096 1175 11130 1209
rect 11096 1107 11130 1141
rect 11096 1039 11130 1073
rect 11096 971 11130 1005
rect 11096 903 11130 937
rect 11096 835 11130 869
rect 11096 767 11130 801
rect 11096 699 11130 733
rect 11096 631 11130 665
rect 11096 563 11130 597
rect 11096 495 11130 529
rect 11096 427 11130 461
rect 11096 359 11130 393
rect 11096 291 11130 325
rect 11192 1175 11226 1209
rect 11192 1107 11226 1141
rect 11192 1039 11226 1073
rect 11192 971 11226 1005
rect 11192 903 11226 937
rect 11192 835 11226 869
rect 11192 767 11226 801
rect 11192 699 11226 733
rect 11192 631 11226 665
rect 11192 563 11226 597
rect 11192 495 11226 529
rect 11192 427 11226 461
rect 11192 359 11226 393
rect 11192 291 11226 325
rect 11288 1175 11322 1209
rect 11288 1107 11322 1141
rect 11288 1039 11322 1073
rect 11288 971 11322 1005
rect 11288 903 11322 937
rect 11288 835 11322 869
rect 11288 767 11322 801
rect 11288 699 11322 733
rect 11288 631 11322 665
rect 11288 563 11322 597
rect 11288 495 11322 529
rect 11288 427 11322 461
rect 11288 359 11322 393
rect 11288 291 11322 325
rect 11384 1175 11418 1209
rect 11384 1107 11418 1141
rect 11384 1039 11418 1073
rect 11384 971 11418 1005
rect 11384 903 11418 937
rect 11384 835 11418 869
rect 11384 767 11418 801
rect 11384 699 11418 733
rect 11384 631 11418 665
rect 11384 563 11418 597
rect 11384 495 11418 529
rect 11384 427 11418 461
rect 11384 359 11418 393
rect 11384 291 11418 325
rect 11480 1175 11514 1209
rect 11480 1107 11514 1141
rect 11480 1039 11514 1073
rect 11480 971 11514 1005
rect 11480 903 11514 937
rect 11480 835 11514 869
rect 11480 767 11514 801
rect 11480 699 11514 733
rect 11480 631 11514 665
rect 11480 563 11514 597
rect 11480 495 11514 529
rect 11480 427 11514 461
rect 11480 359 11514 393
rect 11480 291 11514 325
rect 11576 1175 11610 1209
rect 11576 1107 11610 1141
rect 11576 1039 11610 1073
rect 11576 971 11610 1005
rect 11576 903 11610 937
rect 11576 835 11610 869
rect 11576 767 11610 801
rect 11576 699 11610 733
rect 11576 631 11610 665
rect 11576 563 11610 597
rect 11576 495 11610 529
rect 11576 427 11610 461
rect 11576 359 11610 393
rect 11576 291 11610 325
rect 11672 1175 11706 1209
rect 11672 1107 11706 1141
rect 11672 1039 11706 1073
rect 11672 971 11706 1005
rect 11672 903 11706 937
rect 11672 835 11706 869
rect 11672 767 11706 801
rect 11672 699 11706 733
rect 11672 631 11706 665
rect 11672 563 11706 597
rect 11672 495 11706 529
rect 11672 427 11706 461
rect 11672 359 11706 393
rect 11672 291 11706 325
rect 11768 1175 11802 1209
rect 11768 1107 11802 1141
rect 11768 1039 11802 1073
rect 11768 971 11802 1005
rect 11768 903 11802 937
rect 11768 835 11802 869
rect 11768 767 11802 801
rect 11768 699 11802 733
rect 11768 631 11802 665
rect 11768 563 11802 597
rect 11768 495 11802 529
rect 11768 427 11802 461
rect 11768 359 11802 393
rect 11768 291 11802 325
rect 11864 1175 11898 1209
rect 11864 1107 11898 1141
rect 11864 1039 11898 1073
rect 11864 971 11898 1005
rect 11864 903 11898 937
rect 11864 835 11898 869
rect 11864 767 11898 801
rect 11864 699 11898 733
rect 11864 631 11898 665
rect 11864 563 11898 597
rect 11864 495 11898 529
rect 11864 427 11898 461
rect 11864 359 11898 393
rect 11864 291 11898 325
rect 11960 1175 11994 1209
rect 11960 1107 11994 1141
rect 11960 1039 11994 1073
rect 11960 971 11994 1005
rect 11960 903 11994 937
rect 11960 835 11994 869
rect 11960 767 11994 801
rect 11960 699 11994 733
rect 11960 631 11994 665
rect 11960 563 11994 597
rect 11960 495 11994 529
rect 11960 427 11994 461
rect 11960 359 11994 393
rect 11960 291 11994 325
rect 15422 1227 15456 1261
rect 12056 1175 12090 1209
rect 12056 1107 12090 1141
rect 12056 1039 12090 1073
rect 12056 971 12090 1005
rect 12056 903 12090 937
rect 12056 835 12090 869
rect 12056 767 12090 801
rect 12056 699 12090 733
rect 12056 631 12090 665
rect 12056 563 12090 597
rect 12056 495 12090 529
rect 12056 427 12090 461
rect 12056 359 12090 393
rect 12056 291 12090 325
rect 12388 1149 12422 1183
rect 12388 1081 12422 1115
rect 12388 1013 12422 1047
rect 12388 945 12422 979
rect 12388 877 12422 911
rect 12388 809 12422 843
rect 12388 741 12422 775
rect 12388 673 12422 707
rect 12388 605 12422 639
rect 12388 537 12422 571
rect 12388 469 12422 503
rect 12388 401 12422 435
rect 12388 333 12422 367
rect 12388 265 12422 299
rect 12484 1149 12518 1183
rect 12484 1081 12518 1115
rect 12484 1013 12518 1047
rect 12484 945 12518 979
rect 12484 877 12518 911
rect 12484 809 12518 843
rect 12484 741 12518 775
rect 12484 673 12518 707
rect 12484 605 12518 639
rect 12484 537 12518 571
rect 12484 469 12518 503
rect 12484 401 12518 435
rect 12484 333 12518 367
rect 12484 265 12518 299
rect 12580 1149 12614 1183
rect 12580 1081 12614 1115
rect 12580 1013 12614 1047
rect 12580 945 12614 979
rect 12580 877 12614 911
rect 12580 809 12614 843
rect 12580 741 12614 775
rect 12580 673 12614 707
rect 12580 605 12614 639
rect 12580 537 12614 571
rect 12580 469 12614 503
rect 12580 401 12614 435
rect 12580 333 12614 367
rect 12580 265 12614 299
rect 12676 1149 12710 1183
rect 12676 1081 12710 1115
rect 12676 1013 12710 1047
rect 12676 945 12710 979
rect 12676 877 12710 911
rect 12676 809 12710 843
rect 12676 741 12710 775
rect 12676 673 12710 707
rect 12676 605 12710 639
rect 12676 537 12710 571
rect 12676 469 12710 503
rect 12676 401 12710 435
rect 12676 333 12710 367
rect 12676 265 12710 299
rect 12772 1149 12806 1183
rect 12772 1081 12806 1115
rect 12772 1013 12806 1047
rect 12772 945 12806 979
rect 12772 877 12806 911
rect 12772 809 12806 843
rect 12772 741 12806 775
rect 12772 673 12806 707
rect 12772 605 12806 639
rect 12772 537 12806 571
rect 12772 469 12806 503
rect 12772 401 12806 435
rect 12772 333 12806 367
rect 12772 265 12806 299
rect 12868 1149 12902 1183
rect 12868 1081 12902 1115
rect 12868 1013 12902 1047
rect 12868 945 12902 979
rect 12868 877 12902 911
rect 12868 809 12902 843
rect 12868 741 12902 775
rect 12868 673 12902 707
rect 12868 605 12902 639
rect 12868 537 12902 571
rect 12868 469 12902 503
rect 12868 401 12902 435
rect 12868 333 12902 367
rect 12868 265 12902 299
rect 12964 1149 12998 1183
rect 12964 1081 12998 1115
rect 12964 1013 12998 1047
rect 12964 945 12998 979
rect 12964 877 12998 911
rect 12964 809 12998 843
rect 12964 741 12998 775
rect 12964 673 12998 707
rect 12964 605 12998 639
rect 12964 537 12998 571
rect 12964 469 12998 503
rect 12964 401 12998 435
rect 12964 333 12998 367
rect 12964 265 12998 299
rect 13060 1149 13094 1183
rect 13060 1081 13094 1115
rect 13060 1013 13094 1047
rect 13060 945 13094 979
rect 13060 877 13094 911
rect 13060 809 13094 843
rect 13060 741 13094 775
rect 13060 673 13094 707
rect 13060 605 13094 639
rect 13060 537 13094 571
rect 13060 469 13094 503
rect 13060 401 13094 435
rect 13060 333 13094 367
rect 13060 265 13094 299
rect 13156 1149 13190 1183
rect 13156 1081 13190 1115
rect 13156 1013 13190 1047
rect 13156 945 13190 979
rect 13156 877 13190 911
rect 13156 809 13190 843
rect 13156 741 13190 775
rect 13156 673 13190 707
rect 13156 605 13190 639
rect 13156 537 13190 571
rect 13156 469 13190 503
rect 13156 401 13190 435
rect 13156 333 13190 367
rect 13156 265 13190 299
rect 13252 1149 13286 1183
rect 13252 1081 13286 1115
rect 13252 1013 13286 1047
rect 13252 945 13286 979
rect 13252 877 13286 911
rect 13252 809 13286 843
rect 13252 741 13286 775
rect 13252 673 13286 707
rect 13252 605 13286 639
rect 13252 537 13286 571
rect 13252 469 13286 503
rect 13252 401 13286 435
rect 13252 333 13286 367
rect 13252 265 13286 299
rect 13348 1149 13382 1183
rect 13348 1081 13382 1115
rect 13348 1013 13382 1047
rect 13348 945 13382 979
rect 13348 877 13382 911
rect 13348 809 13382 843
rect 13348 741 13382 775
rect 13348 673 13382 707
rect 13348 605 13382 639
rect 13348 537 13382 571
rect 13348 469 13382 503
rect 13348 401 13382 435
rect 13348 333 13382 367
rect 13348 265 13382 299
rect 13444 1149 13478 1183
rect 13444 1081 13478 1115
rect 13444 1013 13478 1047
rect 13444 945 13478 979
rect 13444 877 13478 911
rect 13444 809 13478 843
rect 13444 741 13478 775
rect 13444 673 13478 707
rect 13444 605 13478 639
rect 13444 537 13478 571
rect 13444 469 13478 503
rect 13444 401 13478 435
rect 13444 333 13478 367
rect 13444 265 13478 299
rect 13540 1149 13574 1183
rect 13540 1081 13574 1115
rect 13540 1013 13574 1047
rect 13540 945 13574 979
rect 13540 877 13574 911
rect 13540 809 13574 843
rect 13540 741 13574 775
rect 13540 673 13574 707
rect 13540 605 13574 639
rect 13540 537 13574 571
rect 13540 469 13574 503
rect 13540 401 13574 435
rect 13540 333 13574 367
rect 13540 265 13574 299
rect 14156 1149 14190 1183
rect 14156 1081 14190 1115
rect 14156 1013 14190 1047
rect 14156 945 14190 979
rect 14156 877 14190 911
rect 14156 809 14190 843
rect 14156 741 14190 775
rect 14156 673 14190 707
rect 14156 605 14190 639
rect 14156 537 14190 571
rect 14156 469 14190 503
rect 14156 401 14190 435
rect 14156 333 14190 367
rect 14156 265 14190 299
rect 14252 1149 14286 1183
rect 14252 1081 14286 1115
rect 14252 1013 14286 1047
rect 14252 945 14286 979
rect 14252 877 14286 911
rect 14252 809 14286 843
rect 14252 741 14286 775
rect 14252 673 14286 707
rect 14252 605 14286 639
rect 14252 537 14286 571
rect 14252 469 14286 503
rect 14252 401 14286 435
rect 14252 333 14286 367
rect 14252 265 14286 299
rect 14348 1149 14382 1183
rect 14348 1081 14382 1115
rect 14348 1013 14382 1047
rect 14348 945 14382 979
rect 14348 877 14382 911
rect 14348 809 14382 843
rect 14348 741 14382 775
rect 14348 673 14382 707
rect 14348 605 14382 639
rect 14348 537 14382 571
rect 14348 469 14382 503
rect 14348 401 14382 435
rect 14348 333 14382 367
rect 14348 265 14382 299
rect 14444 1149 14478 1183
rect 14444 1081 14478 1115
rect 14444 1013 14478 1047
rect 14444 945 14478 979
rect 14444 877 14478 911
rect 14444 809 14478 843
rect 14444 741 14478 775
rect 14444 673 14478 707
rect 14444 605 14478 639
rect 14444 537 14478 571
rect 14444 469 14478 503
rect 14444 401 14478 435
rect 14444 333 14478 367
rect 14444 265 14478 299
rect 14540 1149 14574 1183
rect 14540 1081 14574 1115
rect 14540 1013 14574 1047
rect 14540 945 14574 979
rect 14540 877 14574 911
rect 14540 809 14574 843
rect 14540 741 14574 775
rect 14540 673 14574 707
rect 14540 605 14574 639
rect 14540 537 14574 571
rect 14540 469 14574 503
rect 14540 401 14574 435
rect 14540 333 14574 367
rect 14540 265 14574 299
rect 14636 1149 14670 1183
rect 14636 1081 14670 1115
rect 14636 1013 14670 1047
rect 14636 945 14670 979
rect 14636 877 14670 911
rect 14636 809 14670 843
rect 14636 741 14670 775
rect 14636 673 14670 707
rect 14636 605 14670 639
rect 14636 537 14670 571
rect 14636 469 14670 503
rect 14636 401 14670 435
rect 14636 333 14670 367
rect 14636 265 14670 299
rect 14732 1149 14766 1183
rect 14732 1081 14766 1115
rect 14732 1013 14766 1047
rect 14732 945 14766 979
rect 14732 877 14766 911
rect 14732 809 14766 843
rect 14732 741 14766 775
rect 14732 673 14766 707
rect 14732 605 14766 639
rect 14732 537 14766 571
rect 14732 469 14766 503
rect 14732 401 14766 435
rect 14732 333 14766 367
rect 14732 265 14766 299
rect 14828 1149 14862 1183
rect 14828 1081 14862 1115
rect 14828 1013 14862 1047
rect 14828 945 14862 979
rect 14828 877 14862 911
rect 14828 809 14862 843
rect 14828 741 14862 775
rect 14828 673 14862 707
rect 14828 605 14862 639
rect 14828 537 14862 571
rect 14828 469 14862 503
rect 14828 401 14862 435
rect 14828 333 14862 367
rect 14828 265 14862 299
rect 14924 1149 14958 1183
rect 14924 1081 14958 1115
rect 14924 1013 14958 1047
rect 14924 945 14958 979
rect 14924 877 14958 911
rect 14924 809 14958 843
rect 14924 741 14958 775
rect 14924 673 14958 707
rect 14924 605 14958 639
rect 14924 537 14958 571
rect 14924 469 14958 503
rect 14924 401 14958 435
rect 14924 333 14958 367
rect 14924 265 14958 299
rect 15020 1149 15054 1183
rect 15020 1081 15054 1115
rect 15020 1013 15054 1047
rect 15020 945 15054 979
rect 15020 877 15054 911
rect 15020 809 15054 843
rect 15020 741 15054 775
rect 15020 673 15054 707
rect 15020 605 15054 639
rect 15020 537 15054 571
rect 15020 469 15054 503
rect 15020 401 15054 435
rect 15020 333 15054 367
rect 15020 265 15054 299
rect 15116 1149 15150 1183
rect 15116 1081 15150 1115
rect 15116 1013 15150 1047
rect 15116 945 15150 979
rect 15116 877 15150 911
rect 15116 809 15150 843
rect 15116 741 15150 775
rect 15116 673 15150 707
rect 15116 605 15150 639
rect 15116 537 15150 571
rect 15116 469 15150 503
rect 15116 401 15150 435
rect 15116 333 15150 367
rect 15116 265 15150 299
rect 15212 1149 15246 1183
rect 15212 1081 15246 1115
rect 15212 1013 15246 1047
rect 15212 945 15246 979
rect 15212 877 15246 911
rect 15212 809 15246 843
rect 15212 741 15246 775
rect 15212 673 15246 707
rect 15212 605 15246 639
rect 15212 537 15246 571
rect 15212 469 15246 503
rect 15212 401 15246 435
rect 15212 333 15246 367
rect 15212 265 15246 299
rect 15422 1159 15456 1193
rect 15422 1091 15456 1125
rect 15422 1023 15456 1057
rect 15422 955 15456 989
rect 15422 887 15456 921
rect 15422 819 15456 853
rect 15422 751 15456 785
rect 15422 683 15456 717
rect 15422 615 15456 649
rect 15422 547 15456 581
rect 15422 479 15456 513
rect 15422 411 15456 445
rect 15422 343 15456 377
rect 15422 275 15456 309
rect 15422 207 15456 241
rect 15422 139 15456 173
rect 15510 1227 15544 1261
rect 15510 1159 15544 1193
rect 15510 1091 15544 1125
rect 15510 1023 15544 1057
rect 15510 955 15544 989
rect 15510 887 15544 921
rect 15510 819 15544 853
rect 15510 751 15544 785
rect 15510 683 15544 717
rect 15510 615 15544 649
rect 15510 547 15544 581
rect 15510 479 15544 513
rect 15510 411 15544 445
rect 15510 343 15544 377
rect 15510 275 15544 309
rect 15510 207 15544 241
rect 15510 139 15544 173
<< pdiffc >>
rect 194 6531 228 6565
rect 194 6463 228 6497
rect 194 6395 228 6429
rect 194 6327 228 6361
rect 194 6259 228 6293
rect 194 6191 228 6225
rect 194 6123 228 6157
rect 194 6055 228 6089
rect 194 5987 228 6021
rect -1652 5861 -1618 5895
rect -1652 5793 -1618 5827
rect -1652 5725 -1618 5759
rect -1652 5657 -1618 5691
rect -1652 5589 -1618 5623
rect -1652 5521 -1618 5555
rect -1652 5453 -1618 5487
rect -1652 5385 -1618 5419
rect -1652 5317 -1618 5351
rect -1652 5249 -1618 5283
rect -1652 5181 -1618 5215
rect -1652 5113 -1618 5147
rect -1652 5045 -1618 5079
rect -1652 4977 -1618 5011
rect -1554 5861 -1520 5895
rect -1554 5793 -1520 5827
rect -1554 5725 -1520 5759
rect -1554 5657 -1520 5691
rect -1554 5589 -1520 5623
rect -1554 5521 -1520 5555
rect -1554 5453 -1520 5487
rect -1554 5385 -1520 5419
rect -1554 5317 -1520 5351
rect -1554 5249 -1520 5283
rect -1554 5181 -1520 5215
rect -1554 5113 -1520 5147
rect -1554 5045 -1520 5079
rect -1554 4977 -1520 5011
rect -1456 5861 -1422 5895
rect -1456 5793 -1422 5827
rect -1456 5725 -1422 5759
rect -1456 5657 -1422 5691
rect -1456 5589 -1422 5623
rect -1456 5521 -1422 5555
rect -1456 5453 -1422 5487
rect -1456 5385 -1422 5419
rect -1456 5317 -1422 5351
rect -1456 5249 -1422 5283
rect -1456 5181 -1422 5215
rect -1456 5113 -1422 5147
rect -1456 5045 -1422 5079
rect -1456 4977 -1422 5011
rect -1358 5861 -1324 5895
rect -1358 5793 -1324 5827
rect -1358 5725 -1324 5759
rect -1358 5657 -1324 5691
rect -1358 5589 -1324 5623
rect -1358 5521 -1324 5555
rect -1358 5453 -1324 5487
rect -1358 5385 -1324 5419
rect -1358 5317 -1324 5351
rect -1358 5249 -1324 5283
rect -1358 5181 -1324 5215
rect -1358 5113 -1324 5147
rect -1358 5045 -1324 5079
rect -1358 4977 -1324 5011
rect -1260 5861 -1226 5895
rect -1260 5793 -1226 5827
rect -1260 5725 -1226 5759
rect -1260 5657 -1226 5691
rect -1260 5589 -1226 5623
rect -1260 5521 -1226 5555
rect -1260 5453 -1226 5487
rect -1260 5385 -1226 5419
rect -1260 5317 -1226 5351
rect -1260 5249 -1226 5283
rect -1260 5181 -1226 5215
rect -1260 5113 -1226 5147
rect -1260 5045 -1226 5079
rect -1260 4977 -1226 5011
rect -1162 5861 -1128 5895
rect -1162 5793 -1128 5827
rect -1162 5725 -1128 5759
rect -1162 5657 -1128 5691
rect -1162 5589 -1128 5623
rect -1162 5521 -1128 5555
rect -1162 5453 -1128 5487
rect -1162 5385 -1128 5419
rect -1162 5317 -1128 5351
rect -1162 5249 -1128 5283
rect -1162 5181 -1128 5215
rect -1162 5113 -1128 5147
rect -1162 5045 -1128 5079
rect -1162 4977 -1128 5011
rect -1064 5861 -1030 5895
rect -1064 5793 -1030 5827
rect -1064 5725 -1030 5759
rect -1064 5657 -1030 5691
rect -1064 5589 -1030 5623
rect -1064 5521 -1030 5555
rect -1064 5453 -1030 5487
rect -1064 5385 -1030 5419
rect -1064 5317 -1030 5351
rect -1064 5249 -1030 5283
rect -1064 5181 -1030 5215
rect -1064 5113 -1030 5147
rect -1064 5045 -1030 5079
rect -1064 4977 -1030 5011
rect -966 5861 -932 5895
rect -966 5793 -932 5827
rect -966 5725 -932 5759
rect -966 5657 -932 5691
rect -966 5589 -932 5623
rect -966 5521 -932 5555
rect -966 5453 -932 5487
rect -966 5385 -932 5419
rect -966 5317 -932 5351
rect -966 5249 -932 5283
rect -966 5181 -932 5215
rect -966 5113 -932 5147
rect -966 5045 -932 5079
rect -966 4977 -932 5011
rect -868 5861 -834 5895
rect -868 5793 -834 5827
rect -868 5725 -834 5759
rect -868 5657 -834 5691
rect -868 5589 -834 5623
rect 194 5919 228 5953
rect 194 5851 228 5885
rect 194 5783 228 5817
rect 194 5715 228 5749
rect 194 5647 228 5681
rect 290 6531 324 6565
rect 290 6463 324 6497
rect 290 6395 324 6429
rect 290 6327 324 6361
rect 290 6259 324 6293
rect 290 6191 324 6225
rect 290 6123 324 6157
rect 290 6055 324 6089
rect 290 5987 324 6021
rect 290 5919 324 5953
rect 290 5851 324 5885
rect 290 5783 324 5817
rect 290 5715 324 5749
rect 290 5647 324 5681
rect 386 6531 420 6565
rect 386 6463 420 6497
rect 386 6395 420 6429
rect 386 6327 420 6361
rect 386 6259 420 6293
rect 386 6191 420 6225
rect 386 6123 420 6157
rect 386 6055 420 6089
rect 386 5987 420 6021
rect 386 5919 420 5953
rect 386 5851 420 5885
rect 386 5783 420 5817
rect 386 5715 420 5749
rect 386 5647 420 5681
rect 482 6531 516 6565
rect 482 6463 516 6497
rect 482 6395 516 6429
rect 482 6327 516 6361
rect 482 6259 516 6293
rect 482 6191 516 6225
rect 482 6123 516 6157
rect 482 6055 516 6089
rect 482 5987 516 6021
rect 482 5919 516 5953
rect 482 5851 516 5885
rect 482 5783 516 5817
rect 482 5715 516 5749
rect 482 5647 516 5681
rect 578 6531 612 6565
rect 578 6463 612 6497
rect 578 6395 612 6429
rect 578 6327 612 6361
rect 578 6259 612 6293
rect 578 6191 612 6225
rect 578 6123 612 6157
rect 578 6055 612 6089
rect 578 5987 612 6021
rect 578 5919 612 5953
rect 578 5851 612 5885
rect 578 5783 612 5817
rect 578 5715 612 5749
rect 578 5647 612 5681
rect 674 6531 708 6565
rect 674 6463 708 6497
rect 674 6395 708 6429
rect 674 6327 708 6361
rect 674 6259 708 6293
rect 674 6191 708 6225
rect 674 6123 708 6157
rect 674 6055 708 6089
rect 674 5987 708 6021
rect 674 5919 708 5953
rect 674 5851 708 5885
rect 674 5783 708 5817
rect 674 5715 708 5749
rect 674 5647 708 5681
rect 770 6531 804 6565
rect 770 6463 804 6497
rect 770 6395 804 6429
rect 770 6327 804 6361
rect 770 6259 804 6293
rect 770 6191 804 6225
rect 770 6123 804 6157
rect 770 6055 804 6089
rect 770 5987 804 6021
rect 770 5919 804 5953
rect 770 5851 804 5885
rect 770 5783 804 5817
rect 770 5715 804 5749
rect 770 5647 804 5681
rect 866 6531 900 6565
rect 866 6463 900 6497
rect 866 6395 900 6429
rect 866 6327 900 6361
rect 866 6259 900 6293
rect 866 6191 900 6225
rect 866 6123 900 6157
rect 866 6055 900 6089
rect 866 5987 900 6021
rect 866 5919 900 5953
rect 866 5851 900 5885
rect 866 5783 900 5817
rect 866 5715 900 5749
rect 866 5647 900 5681
rect 962 6531 996 6565
rect 962 6463 996 6497
rect 962 6395 996 6429
rect 962 6327 996 6361
rect 962 6259 996 6293
rect 962 6191 996 6225
rect 962 6123 996 6157
rect 962 6055 996 6089
rect 962 5987 996 6021
rect 962 5919 996 5953
rect 962 5851 996 5885
rect 962 5783 996 5817
rect 962 5715 996 5749
rect 962 5647 996 5681
rect 1058 6531 1092 6565
rect 1058 6463 1092 6497
rect 1058 6395 1092 6429
rect 1058 6327 1092 6361
rect 1058 6259 1092 6293
rect 1058 6191 1092 6225
rect 1058 6123 1092 6157
rect 1058 6055 1092 6089
rect 1058 5987 1092 6021
rect 1058 5919 1092 5953
rect 1058 5851 1092 5885
rect 1058 5783 1092 5817
rect 1058 5715 1092 5749
rect 1058 5647 1092 5681
rect 1154 6531 1188 6565
rect 1154 6463 1188 6497
rect 1154 6395 1188 6429
rect 1154 6327 1188 6361
rect 1154 6259 1188 6293
rect 1154 6191 1188 6225
rect 1154 6123 1188 6157
rect 1154 6055 1188 6089
rect 1154 5987 1188 6021
rect 1154 5919 1188 5953
rect 1154 5851 1188 5885
rect 1154 5783 1188 5817
rect 1154 5715 1188 5749
rect 1154 5647 1188 5681
rect 1250 6531 1284 6565
rect 1250 6463 1284 6497
rect 1250 6395 1284 6429
rect 1250 6327 1284 6361
rect 1250 6259 1284 6293
rect 1250 6191 1284 6225
rect 1250 6123 1284 6157
rect 1250 6055 1284 6089
rect 1250 5987 1284 6021
rect 1250 5919 1284 5953
rect 1250 5851 1284 5885
rect 1250 5783 1284 5817
rect 1250 5715 1284 5749
rect 1250 5647 1284 5681
rect 1346 6531 1380 6565
rect 1346 6463 1380 6497
rect 1346 6395 1380 6429
rect 1346 6327 1380 6361
rect 1346 6259 1380 6293
rect 1346 6191 1380 6225
rect 1346 6123 1380 6157
rect 1346 6055 1380 6089
rect 1346 5987 1380 6021
rect 1346 5919 1380 5953
rect 1346 5851 1380 5885
rect 1346 5783 1380 5817
rect 1346 5715 1380 5749
rect 1346 5647 1380 5681
rect 1960 6527 1994 6561
rect 1960 6459 1994 6493
rect 1960 6391 1994 6425
rect 1960 6323 1994 6357
rect 1960 6255 1994 6289
rect 1960 6187 1994 6221
rect 1960 6119 1994 6153
rect 1960 6051 1994 6085
rect 1960 5983 1994 6017
rect 1960 5915 1994 5949
rect 1960 5847 1994 5881
rect 1960 5779 1994 5813
rect 1960 5711 1994 5745
rect 1960 5643 1994 5677
rect 2056 6527 2090 6561
rect 2056 6459 2090 6493
rect 2056 6391 2090 6425
rect 2056 6323 2090 6357
rect 2056 6255 2090 6289
rect 2056 6187 2090 6221
rect 2056 6119 2090 6153
rect 2056 6051 2090 6085
rect 2056 5983 2090 6017
rect 2056 5915 2090 5949
rect 2056 5847 2090 5881
rect 2056 5779 2090 5813
rect 2056 5711 2090 5745
rect 2056 5643 2090 5677
rect 2152 6527 2186 6561
rect 2152 6459 2186 6493
rect 2152 6391 2186 6425
rect 2152 6323 2186 6357
rect 2152 6255 2186 6289
rect 2152 6187 2186 6221
rect 2152 6119 2186 6153
rect 2152 6051 2186 6085
rect 2152 5983 2186 6017
rect 2152 5915 2186 5949
rect 2152 5847 2186 5881
rect 2152 5779 2186 5813
rect 2152 5711 2186 5745
rect 2152 5643 2186 5677
rect 2248 6527 2282 6561
rect 2248 6459 2282 6493
rect 2248 6391 2282 6425
rect 2248 6323 2282 6357
rect 2248 6255 2282 6289
rect 2248 6187 2282 6221
rect 2248 6119 2282 6153
rect 2248 6051 2282 6085
rect 2248 5983 2282 6017
rect 2248 5915 2282 5949
rect 2248 5847 2282 5881
rect 2248 5779 2282 5813
rect 2248 5711 2282 5745
rect 2248 5643 2282 5677
rect 2344 6527 2378 6561
rect 2344 6459 2378 6493
rect 2344 6391 2378 6425
rect 2344 6323 2378 6357
rect 2344 6255 2378 6289
rect 2344 6187 2378 6221
rect 2344 6119 2378 6153
rect 2344 6051 2378 6085
rect 2344 5983 2378 6017
rect 2344 5915 2378 5949
rect 2344 5847 2378 5881
rect 2344 5779 2378 5813
rect 2344 5711 2378 5745
rect 2344 5643 2378 5677
rect 2440 6527 2474 6561
rect 2440 6459 2474 6493
rect 2440 6391 2474 6425
rect 2440 6323 2474 6357
rect 2440 6255 2474 6289
rect 2440 6187 2474 6221
rect 2440 6119 2474 6153
rect 2440 6051 2474 6085
rect 2440 5983 2474 6017
rect 2440 5915 2474 5949
rect 2440 5847 2474 5881
rect 2440 5779 2474 5813
rect 2440 5711 2474 5745
rect 2440 5643 2474 5677
rect 2536 6527 2570 6561
rect 2536 6459 2570 6493
rect 2536 6391 2570 6425
rect 2536 6323 2570 6357
rect 2536 6255 2570 6289
rect 2536 6187 2570 6221
rect 2536 6119 2570 6153
rect 2536 6051 2570 6085
rect 2536 5983 2570 6017
rect 2536 5915 2570 5949
rect 2536 5847 2570 5881
rect 2536 5779 2570 5813
rect 2536 5711 2570 5745
rect 2536 5643 2570 5677
rect 2632 6527 2666 6561
rect 2632 6459 2666 6493
rect 2632 6391 2666 6425
rect 2632 6323 2666 6357
rect 2632 6255 2666 6289
rect 2632 6187 2666 6221
rect 2632 6119 2666 6153
rect 2632 6051 2666 6085
rect 2632 5983 2666 6017
rect 2632 5915 2666 5949
rect 2632 5847 2666 5881
rect 2632 5779 2666 5813
rect 2632 5711 2666 5745
rect 2632 5643 2666 5677
rect 2728 6527 2762 6561
rect 2728 6459 2762 6493
rect 2728 6391 2762 6425
rect 2728 6323 2762 6357
rect 2728 6255 2762 6289
rect 2728 6187 2762 6221
rect 2728 6119 2762 6153
rect 2728 6051 2762 6085
rect 2728 5983 2762 6017
rect 2728 5915 2762 5949
rect 2728 5847 2762 5881
rect 2728 5779 2762 5813
rect 2728 5711 2762 5745
rect 2728 5643 2762 5677
rect 3150 6515 3184 6549
rect 3150 6447 3184 6481
rect 3150 6379 3184 6413
rect 3150 6311 3184 6345
rect 3150 6243 3184 6277
rect 3150 6175 3184 6209
rect 3150 6107 3184 6141
rect 3150 6039 3184 6073
rect 3150 5971 3184 6005
rect 3150 5903 3184 5937
rect 3150 5835 3184 5869
rect 3150 5767 3184 5801
rect 3150 5699 3184 5733
rect 3150 5631 3184 5665
rect 3246 6515 3280 6549
rect 3246 6447 3280 6481
rect 3246 6379 3280 6413
rect 3246 6311 3280 6345
rect 3246 6243 3280 6277
rect 3246 6175 3280 6209
rect 3246 6107 3280 6141
rect 3246 6039 3280 6073
rect 3246 5971 3280 6005
rect 3246 5903 3280 5937
rect 3246 5835 3280 5869
rect 3246 5767 3280 5801
rect 3246 5699 3280 5733
rect 3246 5631 3280 5665
rect 3342 6515 3376 6549
rect 3342 6447 3376 6481
rect 3342 6379 3376 6413
rect 3342 6311 3376 6345
rect 3342 6243 3376 6277
rect 3342 6175 3376 6209
rect 3342 6107 3376 6141
rect 3342 6039 3376 6073
rect 3342 5971 3376 6005
rect 3342 5903 3376 5937
rect 3342 5835 3376 5869
rect 3342 5767 3376 5801
rect 3342 5699 3376 5733
rect 3342 5631 3376 5665
rect 3438 6515 3472 6549
rect 3438 6447 3472 6481
rect 3438 6379 3472 6413
rect 3438 6311 3472 6345
rect 3438 6243 3472 6277
rect 3438 6175 3472 6209
rect 3438 6107 3472 6141
rect 3438 6039 3472 6073
rect 3438 5971 3472 6005
rect 3438 5903 3472 5937
rect 3438 5835 3472 5869
rect 3438 5767 3472 5801
rect 3438 5699 3472 5733
rect 3438 5631 3472 5665
rect 3534 6515 3568 6549
rect 3534 6447 3568 6481
rect 3534 6379 3568 6413
rect 3534 6311 3568 6345
rect 3534 6243 3568 6277
rect 3534 6175 3568 6209
rect 3534 6107 3568 6141
rect 3534 6039 3568 6073
rect 3534 5971 3568 6005
rect 3534 5903 3568 5937
rect 3534 5835 3568 5869
rect 3534 5767 3568 5801
rect 3534 5699 3568 5733
rect 3534 5631 3568 5665
rect 3630 6515 3664 6549
rect 3630 6447 3664 6481
rect 3630 6379 3664 6413
rect 3630 6311 3664 6345
rect 3630 6243 3664 6277
rect 3630 6175 3664 6209
rect 3630 6107 3664 6141
rect 3630 6039 3664 6073
rect 3630 5971 3664 6005
rect 3630 5903 3664 5937
rect 3630 5835 3664 5869
rect 3630 5767 3664 5801
rect 3630 5699 3664 5733
rect 3630 5631 3664 5665
rect 3726 6515 3760 6549
rect 3726 6447 3760 6481
rect 3726 6379 3760 6413
rect 3726 6311 3760 6345
rect 3726 6243 3760 6277
rect 3726 6175 3760 6209
rect 3726 6107 3760 6141
rect 3726 6039 3760 6073
rect 3726 5971 3760 6005
rect 3726 5903 3760 5937
rect 3726 5835 3760 5869
rect 3726 5767 3760 5801
rect 3726 5699 3760 5733
rect 3726 5631 3760 5665
rect 3822 6515 3856 6549
rect 3822 6447 3856 6481
rect 3822 6379 3856 6413
rect 3822 6311 3856 6345
rect 3822 6243 3856 6277
rect 3822 6175 3856 6209
rect 3822 6107 3856 6141
rect 3822 6039 3856 6073
rect 3822 5971 3856 6005
rect 3822 5903 3856 5937
rect 3822 5835 3856 5869
rect 3822 5767 3856 5801
rect 3822 5699 3856 5733
rect 3822 5631 3856 5665
rect 3918 6515 3952 6549
rect 3918 6447 3952 6481
rect 3918 6379 3952 6413
rect 3918 6311 3952 6345
rect 3918 6243 3952 6277
rect 3918 6175 3952 6209
rect 3918 6107 3952 6141
rect 3918 6039 3952 6073
rect 3918 5971 3952 6005
rect 3918 5903 3952 5937
rect 3918 5835 3952 5869
rect 3918 5767 3952 5801
rect 3918 5699 3952 5733
rect 3918 5631 3952 5665
rect 4014 6515 4048 6549
rect 4014 6447 4048 6481
rect 4014 6379 4048 6413
rect 4014 6311 4048 6345
rect 4014 6243 4048 6277
rect 4014 6175 4048 6209
rect 4014 6107 4048 6141
rect 4014 6039 4048 6073
rect 4014 5971 4048 6005
rect 4014 5903 4048 5937
rect 4014 5835 4048 5869
rect 4014 5767 4048 5801
rect 4014 5699 4048 5733
rect 4014 5631 4048 5665
rect 4110 6515 4144 6549
rect 4110 6447 4144 6481
rect 4110 6379 4144 6413
rect 4110 6311 4144 6345
rect 4110 6243 4144 6277
rect 4110 6175 4144 6209
rect 4110 6107 4144 6141
rect 4110 6039 4144 6073
rect 4110 5971 4144 6005
rect 4110 5903 4144 5937
rect 4110 5835 4144 5869
rect 4110 5767 4144 5801
rect 4110 5699 4144 5733
rect 4110 5631 4144 5665
rect 4206 6515 4240 6549
rect 4206 6447 4240 6481
rect 4206 6379 4240 6413
rect 4206 6311 4240 6345
rect 4206 6243 4240 6277
rect 4206 6175 4240 6209
rect 4206 6107 4240 6141
rect 4206 6039 4240 6073
rect 4206 5971 4240 6005
rect 4206 5903 4240 5937
rect 4206 5835 4240 5869
rect 4206 5767 4240 5801
rect 4206 5699 4240 5733
rect 4206 5631 4240 5665
rect 4302 6515 4336 6549
rect 4302 6447 4336 6481
rect 4302 6379 4336 6413
rect 4302 6311 4336 6345
rect 4302 6243 4336 6277
rect 4302 6175 4336 6209
rect 4302 6107 4336 6141
rect 4302 6039 4336 6073
rect 4302 5971 4336 6005
rect 4302 5903 4336 5937
rect 4302 5835 4336 5869
rect 4302 5767 4336 5801
rect 4302 5699 4336 5733
rect 4302 5631 4336 5665
rect 4916 6511 4950 6545
rect 4916 6443 4950 6477
rect 4916 6375 4950 6409
rect 4916 6307 4950 6341
rect 4916 6239 4950 6273
rect 4916 6171 4950 6205
rect 4916 6103 4950 6137
rect 4916 6035 4950 6069
rect 4916 5967 4950 6001
rect 4916 5899 4950 5933
rect 4916 5831 4950 5865
rect 4916 5763 4950 5797
rect 4916 5695 4950 5729
rect 4916 5627 4950 5661
rect 5012 6511 5046 6545
rect 5012 6443 5046 6477
rect 5012 6375 5046 6409
rect 5012 6307 5046 6341
rect 5012 6239 5046 6273
rect 5012 6171 5046 6205
rect 5012 6103 5046 6137
rect 5012 6035 5046 6069
rect 5012 5967 5046 6001
rect 5012 5899 5046 5933
rect 5012 5831 5046 5865
rect 5012 5763 5046 5797
rect 5012 5695 5046 5729
rect 5012 5627 5046 5661
rect 5108 6511 5142 6545
rect 5108 6443 5142 6477
rect 5108 6375 5142 6409
rect 5108 6307 5142 6341
rect 5108 6239 5142 6273
rect 5108 6171 5142 6205
rect 5108 6103 5142 6137
rect 5108 6035 5142 6069
rect 5108 5967 5142 6001
rect 5108 5899 5142 5933
rect 5108 5831 5142 5865
rect 5108 5763 5142 5797
rect 5108 5695 5142 5729
rect 5108 5627 5142 5661
rect 5204 6511 5238 6545
rect 5204 6443 5238 6477
rect 5204 6375 5238 6409
rect 5204 6307 5238 6341
rect 5204 6239 5238 6273
rect 5204 6171 5238 6205
rect 5204 6103 5238 6137
rect 5204 6035 5238 6069
rect 5204 5967 5238 6001
rect 5204 5899 5238 5933
rect 5204 5831 5238 5865
rect 5204 5763 5238 5797
rect 5204 5695 5238 5729
rect 5204 5627 5238 5661
rect 5300 6511 5334 6545
rect 5300 6443 5334 6477
rect 5300 6375 5334 6409
rect 5300 6307 5334 6341
rect 5300 6239 5334 6273
rect 5300 6171 5334 6205
rect 5300 6103 5334 6137
rect 5300 6035 5334 6069
rect 5300 5967 5334 6001
rect 5300 5899 5334 5933
rect 5300 5831 5334 5865
rect 5300 5763 5334 5797
rect 5300 5695 5334 5729
rect 5300 5627 5334 5661
rect 5396 6511 5430 6545
rect 5396 6443 5430 6477
rect 5396 6375 5430 6409
rect 5396 6307 5430 6341
rect 5396 6239 5430 6273
rect 5396 6171 5430 6205
rect 5396 6103 5430 6137
rect 5396 6035 5430 6069
rect 5396 5967 5430 6001
rect 5396 5899 5430 5933
rect 5396 5831 5430 5865
rect 5396 5763 5430 5797
rect 5396 5695 5430 5729
rect 5396 5627 5430 5661
rect 5492 6511 5526 6545
rect 5492 6443 5526 6477
rect 5492 6375 5526 6409
rect 5492 6307 5526 6341
rect 5492 6239 5526 6273
rect 5492 6171 5526 6205
rect 5492 6103 5526 6137
rect 5492 6035 5526 6069
rect 5492 5967 5526 6001
rect 5492 5899 5526 5933
rect 5492 5831 5526 5865
rect 5492 5763 5526 5797
rect 5492 5695 5526 5729
rect 5492 5627 5526 5661
rect 5588 6511 5622 6545
rect 5588 6443 5622 6477
rect 5588 6375 5622 6409
rect 5588 6307 5622 6341
rect 5588 6239 5622 6273
rect 5588 6171 5622 6205
rect 5588 6103 5622 6137
rect 5588 6035 5622 6069
rect 5588 5967 5622 6001
rect 5588 5899 5622 5933
rect 5588 5831 5622 5865
rect 5588 5763 5622 5797
rect 5588 5695 5622 5729
rect 5588 5627 5622 5661
rect 5684 6511 5718 6545
rect 5684 6443 5718 6477
rect 5684 6375 5718 6409
rect 5684 6307 5718 6341
rect 5684 6239 5718 6273
rect 5684 6171 5718 6205
rect 5684 6103 5718 6137
rect 5684 6035 5718 6069
rect 5684 5967 5718 6001
rect 5684 5899 5718 5933
rect 5684 5831 5718 5865
rect 5684 5763 5718 5797
rect 5684 5695 5718 5729
rect 5684 5627 5718 5661
rect 6180 6515 6214 6549
rect 6180 6447 6214 6481
rect 6180 6379 6214 6413
rect 6180 6311 6214 6345
rect 6180 6243 6214 6277
rect 6180 6175 6214 6209
rect 6180 6107 6214 6141
rect 6180 6039 6214 6073
rect 6180 5971 6214 6005
rect 6180 5903 6214 5937
rect 6180 5835 6214 5869
rect 6180 5767 6214 5801
rect 6180 5699 6214 5733
rect 6180 5631 6214 5665
rect 6276 6515 6310 6549
rect 6276 6447 6310 6481
rect 6276 6379 6310 6413
rect 6276 6311 6310 6345
rect 6276 6243 6310 6277
rect 6276 6175 6310 6209
rect 6276 6107 6310 6141
rect 6276 6039 6310 6073
rect 6276 5971 6310 6005
rect 6276 5903 6310 5937
rect 6276 5835 6310 5869
rect 6276 5767 6310 5801
rect 6276 5699 6310 5733
rect 6276 5631 6310 5665
rect 6372 6515 6406 6549
rect 6372 6447 6406 6481
rect 6372 6379 6406 6413
rect 6372 6311 6406 6345
rect 6372 6243 6406 6277
rect 6372 6175 6406 6209
rect 6372 6107 6406 6141
rect 6372 6039 6406 6073
rect 6372 5971 6406 6005
rect 6372 5903 6406 5937
rect 6372 5835 6406 5869
rect 6372 5767 6406 5801
rect 6372 5699 6406 5733
rect 6372 5631 6406 5665
rect 6468 6515 6502 6549
rect 6468 6447 6502 6481
rect 6468 6379 6502 6413
rect 6468 6311 6502 6345
rect 6468 6243 6502 6277
rect 6468 6175 6502 6209
rect 6468 6107 6502 6141
rect 6468 6039 6502 6073
rect 6468 5971 6502 6005
rect 6468 5903 6502 5937
rect 6468 5835 6502 5869
rect 6468 5767 6502 5801
rect 6468 5699 6502 5733
rect 6468 5631 6502 5665
rect 6564 6515 6598 6549
rect 6564 6447 6598 6481
rect 6564 6379 6598 6413
rect 6564 6311 6598 6345
rect 6564 6243 6598 6277
rect 6564 6175 6598 6209
rect 6564 6107 6598 6141
rect 6564 6039 6598 6073
rect 6564 5971 6598 6005
rect 6564 5903 6598 5937
rect 6564 5835 6598 5869
rect 6564 5767 6598 5801
rect 6564 5699 6598 5733
rect 6564 5631 6598 5665
rect 6660 6515 6694 6549
rect 6660 6447 6694 6481
rect 6660 6379 6694 6413
rect 6660 6311 6694 6345
rect 6660 6243 6694 6277
rect 6660 6175 6694 6209
rect 6660 6107 6694 6141
rect 6660 6039 6694 6073
rect 6660 5971 6694 6005
rect 6660 5903 6694 5937
rect 6660 5835 6694 5869
rect 6660 5767 6694 5801
rect 6660 5699 6694 5733
rect 6660 5631 6694 5665
rect 6756 6515 6790 6549
rect 6756 6447 6790 6481
rect 6756 6379 6790 6413
rect 6756 6311 6790 6345
rect 6756 6243 6790 6277
rect 6756 6175 6790 6209
rect 6756 6107 6790 6141
rect 6756 6039 6790 6073
rect 6756 5971 6790 6005
rect 6756 5903 6790 5937
rect 6756 5835 6790 5869
rect 6756 5767 6790 5801
rect 6756 5699 6790 5733
rect 6756 5631 6790 5665
rect 6852 6515 6886 6549
rect 6852 6447 6886 6481
rect 6852 6379 6886 6413
rect 6852 6311 6886 6345
rect 6852 6243 6886 6277
rect 6852 6175 6886 6209
rect 6852 6107 6886 6141
rect 6852 6039 6886 6073
rect 6852 5971 6886 6005
rect 6852 5903 6886 5937
rect 6852 5835 6886 5869
rect 6852 5767 6886 5801
rect 6852 5699 6886 5733
rect 6852 5631 6886 5665
rect 6948 6515 6982 6549
rect 6948 6447 6982 6481
rect 6948 6379 6982 6413
rect 6948 6311 6982 6345
rect 6948 6243 6982 6277
rect 6948 6175 6982 6209
rect 6948 6107 6982 6141
rect 6948 6039 6982 6073
rect 6948 5971 6982 6005
rect 6948 5903 6982 5937
rect 6948 5835 6982 5869
rect 6948 5767 6982 5801
rect 6948 5699 6982 5733
rect 6948 5631 6982 5665
rect 7044 6515 7078 6549
rect 7044 6447 7078 6481
rect 7044 6379 7078 6413
rect 7044 6311 7078 6345
rect 7044 6243 7078 6277
rect 7044 6175 7078 6209
rect 7044 6107 7078 6141
rect 7044 6039 7078 6073
rect 7044 5971 7078 6005
rect 7044 5903 7078 5937
rect 7044 5835 7078 5869
rect 7044 5767 7078 5801
rect 7044 5699 7078 5733
rect 7044 5631 7078 5665
rect 7140 6515 7174 6549
rect 7140 6447 7174 6481
rect 7140 6379 7174 6413
rect 7140 6311 7174 6345
rect 7140 6243 7174 6277
rect 7140 6175 7174 6209
rect 7140 6107 7174 6141
rect 7140 6039 7174 6073
rect 7140 5971 7174 6005
rect 7140 5903 7174 5937
rect 7140 5835 7174 5869
rect 7140 5767 7174 5801
rect 7140 5699 7174 5733
rect 7140 5631 7174 5665
rect 7236 6515 7270 6549
rect 7236 6447 7270 6481
rect 7236 6379 7270 6413
rect 7236 6311 7270 6345
rect 7236 6243 7270 6277
rect 7236 6175 7270 6209
rect 7236 6107 7270 6141
rect 7236 6039 7270 6073
rect 7236 5971 7270 6005
rect 7236 5903 7270 5937
rect 7236 5835 7270 5869
rect 7236 5767 7270 5801
rect 7236 5699 7270 5733
rect 7236 5631 7270 5665
rect 7332 6515 7366 6549
rect 7332 6447 7366 6481
rect 7332 6379 7366 6413
rect 7332 6311 7366 6345
rect 7332 6243 7366 6277
rect 7332 6175 7366 6209
rect 7332 6107 7366 6141
rect 7332 6039 7366 6073
rect 7332 5971 7366 6005
rect 7332 5903 7366 5937
rect 7332 5835 7366 5869
rect 7332 5767 7366 5801
rect 7332 5699 7366 5733
rect 7332 5631 7366 5665
rect 7946 6511 7980 6545
rect 7946 6443 7980 6477
rect 7946 6375 7980 6409
rect 7946 6307 7980 6341
rect 7946 6239 7980 6273
rect 7946 6171 7980 6205
rect 7946 6103 7980 6137
rect 7946 6035 7980 6069
rect 7946 5967 7980 6001
rect 7946 5899 7980 5933
rect 7946 5831 7980 5865
rect 7946 5763 7980 5797
rect 7946 5695 7980 5729
rect 7946 5627 7980 5661
rect 8042 6511 8076 6545
rect 8042 6443 8076 6477
rect 8042 6375 8076 6409
rect 8042 6307 8076 6341
rect 8042 6239 8076 6273
rect 8042 6171 8076 6205
rect 8042 6103 8076 6137
rect 8042 6035 8076 6069
rect 8042 5967 8076 6001
rect 8042 5899 8076 5933
rect 8042 5831 8076 5865
rect 8042 5763 8076 5797
rect 8042 5695 8076 5729
rect 8042 5627 8076 5661
rect 8138 6511 8172 6545
rect 8138 6443 8172 6477
rect 8138 6375 8172 6409
rect 8138 6307 8172 6341
rect 8138 6239 8172 6273
rect 8138 6171 8172 6205
rect 8138 6103 8172 6137
rect 8138 6035 8172 6069
rect 8138 5967 8172 6001
rect 8138 5899 8172 5933
rect 8138 5831 8172 5865
rect 8138 5763 8172 5797
rect 8138 5695 8172 5729
rect 8138 5627 8172 5661
rect 8234 6511 8268 6545
rect 8234 6443 8268 6477
rect 8234 6375 8268 6409
rect 8234 6307 8268 6341
rect 8234 6239 8268 6273
rect 8234 6171 8268 6205
rect 8234 6103 8268 6137
rect 8234 6035 8268 6069
rect 8234 5967 8268 6001
rect 8234 5899 8268 5933
rect 8234 5831 8268 5865
rect 8234 5763 8268 5797
rect 8234 5695 8268 5729
rect 8234 5627 8268 5661
rect 8330 6511 8364 6545
rect 8330 6443 8364 6477
rect 8330 6375 8364 6409
rect 8330 6307 8364 6341
rect 8330 6239 8364 6273
rect 8330 6171 8364 6205
rect 8330 6103 8364 6137
rect 8330 6035 8364 6069
rect 8330 5967 8364 6001
rect 8330 5899 8364 5933
rect 8330 5831 8364 5865
rect 8330 5763 8364 5797
rect 8330 5695 8364 5729
rect 8330 5627 8364 5661
rect 8426 6511 8460 6545
rect 8426 6443 8460 6477
rect 8426 6375 8460 6409
rect 8426 6307 8460 6341
rect 8426 6239 8460 6273
rect 8426 6171 8460 6205
rect 8426 6103 8460 6137
rect 8426 6035 8460 6069
rect 8426 5967 8460 6001
rect 8426 5899 8460 5933
rect 8426 5831 8460 5865
rect 8426 5763 8460 5797
rect 8426 5695 8460 5729
rect 8426 5627 8460 5661
rect 8522 6511 8556 6545
rect 8522 6443 8556 6477
rect 8522 6375 8556 6409
rect 8522 6307 8556 6341
rect 8522 6239 8556 6273
rect 8522 6171 8556 6205
rect 8522 6103 8556 6137
rect 8522 6035 8556 6069
rect 8522 5967 8556 6001
rect 8522 5899 8556 5933
rect 8522 5831 8556 5865
rect 8522 5763 8556 5797
rect 8522 5695 8556 5729
rect 8522 5627 8556 5661
rect 8618 6511 8652 6545
rect 8618 6443 8652 6477
rect 8618 6375 8652 6409
rect 8618 6307 8652 6341
rect 8618 6239 8652 6273
rect 8618 6171 8652 6205
rect 8618 6103 8652 6137
rect 8618 6035 8652 6069
rect 8618 5967 8652 6001
rect 8618 5899 8652 5933
rect 8618 5831 8652 5865
rect 8618 5763 8652 5797
rect 8618 5695 8652 5729
rect 8618 5627 8652 5661
rect 8714 6511 8748 6545
rect 8714 6443 8748 6477
rect 8714 6375 8748 6409
rect 8714 6307 8748 6341
rect 8714 6239 8748 6273
rect 8714 6171 8748 6205
rect 8714 6103 8748 6137
rect 8714 6035 8748 6069
rect 8714 5967 8748 6001
rect 8714 5899 8748 5933
rect 8714 5831 8748 5865
rect 8714 5763 8748 5797
rect 8714 5695 8748 5729
rect 8714 5627 8748 5661
rect 9268 6513 9302 6547
rect 9268 6445 9302 6479
rect 9268 6377 9302 6411
rect 9268 6309 9302 6343
rect 9268 6241 9302 6275
rect 9268 6173 9302 6207
rect 9268 6105 9302 6139
rect 9268 6037 9302 6071
rect 9268 5969 9302 6003
rect 9268 5901 9302 5935
rect 9268 5833 9302 5867
rect 9268 5765 9302 5799
rect 9268 5697 9302 5731
rect 9268 5629 9302 5663
rect 9364 6513 9398 6547
rect 9364 6445 9398 6479
rect 9364 6377 9398 6411
rect 9364 6309 9398 6343
rect 9364 6241 9398 6275
rect 9364 6173 9398 6207
rect 9364 6105 9398 6139
rect 9364 6037 9398 6071
rect 9364 5969 9398 6003
rect 9364 5901 9398 5935
rect 9364 5833 9398 5867
rect 9364 5765 9398 5799
rect 9364 5697 9398 5731
rect 9364 5629 9398 5663
rect 9460 6513 9494 6547
rect 9460 6445 9494 6479
rect 9460 6377 9494 6411
rect 9460 6309 9494 6343
rect 9460 6241 9494 6275
rect 9460 6173 9494 6207
rect 9460 6105 9494 6139
rect 9460 6037 9494 6071
rect 9460 5969 9494 6003
rect 9460 5901 9494 5935
rect 9460 5833 9494 5867
rect 9460 5765 9494 5799
rect 9460 5697 9494 5731
rect 9460 5629 9494 5663
rect 9556 6513 9590 6547
rect 9556 6445 9590 6479
rect 9556 6377 9590 6411
rect 9556 6309 9590 6343
rect 9556 6241 9590 6275
rect 9556 6173 9590 6207
rect 9556 6105 9590 6139
rect 9556 6037 9590 6071
rect 9556 5969 9590 6003
rect 9556 5901 9590 5935
rect 9556 5833 9590 5867
rect 9556 5765 9590 5799
rect 9556 5697 9590 5731
rect 9556 5629 9590 5663
rect 9652 6513 9686 6547
rect 9652 6445 9686 6479
rect 9652 6377 9686 6411
rect 9652 6309 9686 6343
rect 9652 6241 9686 6275
rect 9652 6173 9686 6207
rect 9652 6105 9686 6139
rect 9652 6037 9686 6071
rect 9652 5969 9686 6003
rect 9652 5901 9686 5935
rect 9652 5833 9686 5867
rect 9652 5765 9686 5799
rect 9652 5697 9686 5731
rect 9652 5629 9686 5663
rect 9748 6513 9782 6547
rect 9748 6445 9782 6479
rect 9748 6377 9782 6411
rect 9748 6309 9782 6343
rect 9748 6241 9782 6275
rect 9748 6173 9782 6207
rect 9748 6105 9782 6139
rect 9748 6037 9782 6071
rect 9748 5969 9782 6003
rect 9748 5901 9782 5935
rect 9748 5833 9782 5867
rect 9748 5765 9782 5799
rect 9748 5697 9782 5731
rect 9748 5629 9782 5663
rect 9844 6513 9878 6547
rect 9844 6445 9878 6479
rect 9844 6377 9878 6411
rect 9844 6309 9878 6343
rect 9844 6241 9878 6275
rect 9844 6173 9878 6207
rect 9844 6105 9878 6139
rect 9844 6037 9878 6071
rect 9844 5969 9878 6003
rect 9844 5901 9878 5935
rect 9844 5833 9878 5867
rect 9844 5765 9878 5799
rect 9844 5697 9878 5731
rect 9844 5629 9878 5663
rect 9940 6513 9974 6547
rect 9940 6445 9974 6479
rect 9940 6377 9974 6411
rect 9940 6309 9974 6343
rect 9940 6241 9974 6275
rect 9940 6173 9974 6207
rect 9940 6105 9974 6139
rect 9940 6037 9974 6071
rect 9940 5969 9974 6003
rect 9940 5901 9974 5935
rect 9940 5833 9974 5867
rect 9940 5765 9974 5799
rect 9940 5697 9974 5731
rect 9940 5629 9974 5663
rect 10036 6513 10070 6547
rect 10036 6445 10070 6479
rect 10036 6377 10070 6411
rect 10036 6309 10070 6343
rect 10036 6241 10070 6275
rect 10036 6173 10070 6207
rect 10036 6105 10070 6139
rect 10036 6037 10070 6071
rect 10036 5969 10070 6003
rect 10036 5901 10070 5935
rect 10036 5833 10070 5867
rect 10036 5765 10070 5799
rect 10036 5697 10070 5731
rect 10036 5629 10070 5663
rect 10132 6513 10166 6547
rect 10132 6445 10166 6479
rect 10132 6377 10166 6411
rect 10132 6309 10166 6343
rect 10132 6241 10166 6275
rect 10132 6173 10166 6207
rect 10132 6105 10166 6139
rect 10132 6037 10166 6071
rect 10132 5969 10166 6003
rect 10132 5901 10166 5935
rect 10132 5833 10166 5867
rect 10132 5765 10166 5799
rect 10132 5697 10166 5731
rect 10132 5629 10166 5663
rect 10228 6513 10262 6547
rect 10228 6445 10262 6479
rect 10228 6377 10262 6411
rect 10228 6309 10262 6343
rect 10228 6241 10262 6275
rect 10228 6173 10262 6207
rect 10228 6105 10262 6139
rect 10228 6037 10262 6071
rect 10228 5969 10262 6003
rect 10228 5901 10262 5935
rect 10228 5833 10262 5867
rect 10228 5765 10262 5799
rect 10228 5697 10262 5731
rect 10228 5629 10262 5663
rect 10324 6513 10358 6547
rect 10324 6445 10358 6479
rect 10324 6377 10358 6411
rect 10324 6309 10358 6343
rect 10324 6241 10358 6275
rect 10324 6173 10358 6207
rect 10324 6105 10358 6139
rect 10324 6037 10358 6071
rect 10324 5969 10358 6003
rect 10324 5901 10358 5935
rect 10324 5833 10358 5867
rect 10324 5765 10358 5799
rect 10324 5697 10358 5731
rect 10324 5629 10358 5663
rect 10420 6513 10454 6547
rect 10420 6445 10454 6479
rect 10420 6377 10454 6411
rect 10420 6309 10454 6343
rect 10420 6241 10454 6275
rect 10420 6173 10454 6207
rect 10420 6105 10454 6139
rect 10420 6037 10454 6071
rect 10420 5969 10454 6003
rect 10420 5901 10454 5935
rect 10420 5833 10454 5867
rect 10420 5765 10454 5799
rect 10420 5697 10454 5731
rect 10420 5629 10454 5663
rect 11034 6509 11068 6543
rect 11034 6441 11068 6475
rect 11034 6373 11068 6407
rect 11034 6305 11068 6339
rect 11034 6237 11068 6271
rect 11034 6169 11068 6203
rect 11034 6101 11068 6135
rect 11034 6033 11068 6067
rect 11034 5965 11068 5999
rect 11034 5897 11068 5931
rect 11034 5829 11068 5863
rect 11034 5761 11068 5795
rect 11034 5693 11068 5727
rect 11034 5625 11068 5659
rect 11130 6509 11164 6543
rect 11130 6441 11164 6475
rect 11130 6373 11164 6407
rect 11130 6305 11164 6339
rect 11130 6237 11164 6271
rect 11130 6169 11164 6203
rect 11130 6101 11164 6135
rect 11130 6033 11164 6067
rect 11130 5965 11164 5999
rect 11130 5897 11164 5931
rect 11130 5829 11164 5863
rect 11130 5761 11164 5795
rect 11130 5693 11164 5727
rect 11130 5625 11164 5659
rect 11226 6509 11260 6543
rect 11226 6441 11260 6475
rect 11226 6373 11260 6407
rect 11226 6305 11260 6339
rect 11226 6237 11260 6271
rect 11226 6169 11260 6203
rect 11226 6101 11260 6135
rect 11226 6033 11260 6067
rect 11226 5965 11260 5999
rect 11226 5897 11260 5931
rect 11226 5829 11260 5863
rect 11226 5761 11260 5795
rect 11226 5693 11260 5727
rect 11226 5625 11260 5659
rect 11322 6509 11356 6543
rect 11322 6441 11356 6475
rect 11322 6373 11356 6407
rect 11322 6305 11356 6339
rect 11322 6237 11356 6271
rect 11322 6169 11356 6203
rect 11322 6101 11356 6135
rect 11322 6033 11356 6067
rect 11322 5965 11356 5999
rect 11322 5897 11356 5931
rect 11322 5829 11356 5863
rect 11322 5761 11356 5795
rect 11322 5693 11356 5727
rect 11322 5625 11356 5659
rect 11418 6509 11452 6543
rect 11418 6441 11452 6475
rect 11418 6373 11452 6407
rect 11418 6305 11452 6339
rect 11418 6237 11452 6271
rect 11418 6169 11452 6203
rect 11418 6101 11452 6135
rect 11418 6033 11452 6067
rect 11418 5965 11452 5999
rect 11418 5897 11452 5931
rect 11418 5829 11452 5863
rect 11418 5761 11452 5795
rect 11418 5693 11452 5727
rect 11418 5625 11452 5659
rect 11514 6509 11548 6543
rect 11514 6441 11548 6475
rect 11514 6373 11548 6407
rect 11514 6305 11548 6339
rect 11514 6237 11548 6271
rect 11514 6169 11548 6203
rect 11514 6101 11548 6135
rect 11514 6033 11548 6067
rect 11514 5965 11548 5999
rect 11514 5897 11548 5931
rect 11514 5829 11548 5863
rect 11514 5761 11548 5795
rect 11514 5693 11548 5727
rect 11514 5625 11548 5659
rect 11610 6509 11644 6543
rect 11610 6441 11644 6475
rect 11610 6373 11644 6407
rect 11610 6305 11644 6339
rect 11610 6237 11644 6271
rect 11610 6169 11644 6203
rect 11610 6101 11644 6135
rect 11610 6033 11644 6067
rect 11610 5965 11644 5999
rect 11610 5897 11644 5931
rect 11610 5829 11644 5863
rect 11610 5761 11644 5795
rect 11610 5693 11644 5727
rect 11610 5625 11644 5659
rect 11706 6509 11740 6543
rect 11706 6441 11740 6475
rect 11706 6373 11740 6407
rect 11706 6305 11740 6339
rect 11706 6237 11740 6271
rect 11706 6169 11740 6203
rect 11706 6101 11740 6135
rect 11706 6033 11740 6067
rect 11706 5965 11740 5999
rect 11706 5897 11740 5931
rect 11706 5829 11740 5863
rect 11706 5761 11740 5795
rect 11706 5693 11740 5727
rect 11706 5625 11740 5659
rect 11802 6509 11836 6543
rect 11802 6441 11836 6475
rect 11802 6373 11836 6407
rect 11802 6305 11836 6339
rect 11802 6237 11836 6271
rect 11802 6169 11836 6203
rect 11802 6101 11836 6135
rect 11802 6033 11836 6067
rect 11802 5965 11836 5999
rect 11802 5897 11836 5931
rect 11802 5829 11836 5863
rect 11802 5761 11836 5795
rect 11802 5693 11836 5727
rect 11802 5625 11836 5659
rect 12424 6487 12458 6521
rect 12424 6419 12458 6453
rect 12424 6351 12458 6385
rect 12424 6283 12458 6317
rect 12424 6215 12458 6249
rect 12424 6147 12458 6181
rect 12424 6079 12458 6113
rect 12424 6011 12458 6045
rect 12424 5943 12458 5977
rect 12424 5875 12458 5909
rect 12424 5807 12458 5841
rect 12424 5739 12458 5773
rect 12424 5671 12458 5705
rect 12424 5603 12458 5637
rect 12520 6487 12554 6521
rect 12520 6419 12554 6453
rect 12520 6351 12554 6385
rect 12520 6283 12554 6317
rect 12520 6215 12554 6249
rect 12520 6147 12554 6181
rect 12520 6079 12554 6113
rect 12520 6011 12554 6045
rect 12520 5943 12554 5977
rect 12520 5875 12554 5909
rect 12520 5807 12554 5841
rect 12520 5739 12554 5773
rect 12520 5671 12554 5705
rect 12520 5603 12554 5637
rect 12616 6487 12650 6521
rect 12616 6419 12650 6453
rect 12616 6351 12650 6385
rect 12616 6283 12650 6317
rect 12616 6215 12650 6249
rect 12616 6147 12650 6181
rect 12616 6079 12650 6113
rect 12616 6011 12650 6045
rect 12616 5943 12650 5977
rect 12616 5875 12650 5909
rect 12616 5807 12650 5841
rect 12616 5739 12650 5773
rect 12616 5671 12650 5705
rect 12616 5603 12650 5637
rect 12712 6487 12746 6521
rect 12712 6419 12746 6453
rect 12712 6351 12746 6385
rect 12712 6283 12746 6317
rect 12712 6215 12746 6249
rect 12712 6147 12746 6181
rect 12712 6079 12746 6113
rect 12712 6011 12746 6045
rect 12712 5943 12746 5977
rect 12712 5875 12746 5909
rect 12712 5807 12746 5841
rect 12712 5739 12746 5773
rect 12712 5671 12746 5705
rect 12712 5603 12746 5637
rect 12808 6487 12842 6521
rect 12808 6419 12842 6453
rect 12808 6351 12842 6385
rect 12808 6283 12842 6317
rect 12808 6215 12842 6249
rect 12808 6147 12842 6181
rect 12808 6079 12842 6113
rect 12808 6011 12842 6045
rect 12808 5943 12842 5977
rect 12808 5875 12842 5909
rect 12808 5807 12842 5841
rect 12808 5739 12842 5773
rect 12808 5671 12842 5705
rect 12808 5603 12842 5637
rect 12904 6487 12938 6521
rect 12904 6419 12938 6453
rect 12904 6351 12938 6385
rect 12904 6283 12938 6317
rect 12904 6215 12938 6249
rect 12904 6147 12938 6181
rect 12904 6079 12938 6113
rect 12904 6011 12938 6045
rect 12904 5943 12938 5977
rect 12904 5875 12938 5909
rect 12904 5807 12938 5841
rect 12904 5739 12938 5773
rect 12904 5671 12938 5705
rect 12904 5603 12938 5637
rect 13000 6487 13034 6521
rect 13000 6419 13034 6453
rect 13000 6351 13034 6385
rect 13000 6283 13034 6317
rect 13000 6215 13034 6249
rect 13000 6147 13034 6181
rect 13000 6079 13034 6113
rect 13000 6011 13034 6045
rect 13000 5943 13034 5977
rect 13000 5875 13034 5909
rect 13000 5807 13034 5841
rect 13000 5739 13034 5773
rect 13000 5671 13034 5705
rect 13000 5603 13034 5637
rect 13096 6487 13130 6521
rect 13096 6419 13130 6453
rect 13096 6351 13130 6385
rect 13096 6283 13130 6317
rect 13096 6215 13130 6249
rect 13096 6147 13130 6181
rect 13096 6079 13130 6113
rect 13096 6011 13130 6045
rect 13096 5943 13130 5977
rect 13096 5875 13130 5909
rect 13096 5807 13130 5841
rect 13096 5739 13130 5773
rect 13096 5671 13130 5705
rect 13096 5603 13130 5637
rect 13192 6487 13226 6521
rect 13192 6419 13226 6453
rect 13192 6351 13226 6385
rect 13192 6283 13226 6317
rect 13192 6215 13226 6249
rect 13192 6147 13226 6181
rect 13192 6079 13226 6113
rect 13192 6011 13226 6045
rect 13192 5943 13226 5977
rect 13192 5875 13226 5909
rect 13192 5807 13226 5841
rect 13192 5739 13226 5773
rect 13192 5671 13226 5705
rect 13192 5603 13226 5637
rect 13288 6487 13322 6521
rect 13288 6419 13322 6453
rect 13288 6351 13322 6385
rect 13288 6283 13322 6317
rect 13288 6215 13322 6249
rect 13288 6147 13322 6181
rect 13288 6079 13322 6113
rect 13288 6011 13322 6045
rect 13288 5943 13322 5977
rect 13288 5875 13322 5909
rect 13288 5807 13322 5841
rect 13288 5739 13322 5773
rect 13288 5671 13322 5705
rect 13288 5603 13322 5637
rect 13384 6487 13418 6521
rect 13384 6419 13418 6453
rect 13384 6351 13418 6385
rect 13384 6283 13418 6317
rect 13384 6215 13418 6249
rect 13384 6147 13418 6181
rect 13384 6079 13418 6113
rect 13384 6011 13418 6045
rect 13384 5943 13418 5977
rect 13384 5875 13418 5909
rect 13384 5807 13418 5841
rect 13384 5739 13418 5773
rect 13384 5671 13418 5705
rect 13384 5603 13418 5637
rect 13480 6487 13514 6521
rect 13480 6419 13514 6453
rect 13480 6351 13514 6385
rect 13480 6283 13514 6317
rect 13480 6215 13514 6249
rect 13480 6147 13514 6181
rect 13480 6079 13514 6113
rect 13480 6011 13514 6045
rect 13480 5943 13514 5977
rect 13480 5875 13514 5909
rect 13480 5807 13514 5841
rect 13480 5739 13514 5773
rect 13480 5671 13514 5705
rect 13480 5603 13514 5637
rect 13576 6487 13610 6521
rect 13576 6419 13610 6453
rect 13576 6351 13610 6385
rect 13576 6283 13610 6317
rect 13576 6215 13610 6249
rect 13576 6147 13610 6181
rect 13576 6079 13610 6113
rect 13576 6011 13610 6045
rect 13576 5943 13610 5977
rect 13576 5875 13610 5909
rect 13576 5807 13610 5841
rect 13576 5739 13610 5773
rect 13576 5671 13610 5705
rect 13576 5603 13610 5637
rect 14190 6483 14224 6517
rect 14190 6415 14224 6449
rect 14190 6347 14224 6381
rect 14190 6279 14224 6313
rect 14190 6211 14224 6245
rect 14190 6143 14224 6177
rect 14190 6075 14224 6109
rect 14190 6007 14224 6041
rect 14190 5939 14224 5973
rect 14190 5871 14224 5905
rect 14190 5803 14224 5837
rect 14190 5735 14224 5769
rect 14190 5667 14224 5701
rect 14190 5599 14224 5633
rect -868 5521 -834 5555
rect 14286 6483 14320 6517
rect 14286 6415 14320 6449
rect 14286 6347 14320 6381
rect 14286 6279 14320 6313
rect 14286 6211 14320 6245
rect 14286 6143 14320 6177
rect 14286 6075 14320 6109
rect 14286 6007 14320 6041
rect 14286 5939 14320 5973
rect 14286 5871 14320 5905
rect 14286 5803 14320 5837
rect 14286 5735 14320 5769
rect 14286 5667 14320 5701
rect 14286 5599 14320 5633
rect 14382 6483 14416 6517
rect 14382 6415 14416 6449
rect 14382 6347 14416 6381
rect 14382 6279 14416 6313
rect 14382 6211 14416 6245
rect 14382 6143 14416 6177
rect 14382 6075 14416 6109
rect 14382 6007 14416 6041
rect 14382 5939 14416 5973
rect 14382 5871 14416 5905
rect 14382 5803 14416 5837
rect 14382 5735 14416 5769
rect 14382 5667 14416 5701
rect 14382 5599 14416 5633
rect 14478 6483 14512 6517
rect 14478 6415 14512 6449
rect 14478 6347 14512 6381
rect 14478 6279 14512 6313
rect 14478 6211 14512 6245
rect 14478 6143 14512 6177
rect 14478 6075 14512 6109
rect 14478 6007 14512 6041
rect 14478 5939 14512 5973
rect 14478 5871 14512 5905
rect 14478 5803 14512 5837
rect 14478 5735 14512 5769
rect 14478 5667 14512 5701
rect 14478 5599 14512 5633
rect 14574 6483 14608 6517
rect 14574 6415 14608 6449
rect 14574 6347 14608 6381
rect 14574 6279 14608 6313
rect 14574 6211 14608 6245
rect 14574 6143 14608 6177
rect 14574 6075 14608 6109
rect 14574 6007 14608 6041
rect 14574 5939 14608 5973
rect 14574 5871 14608 5905
rect 14574 5803 14608 5837
rect 14574 5735 14608 5769
rect 14574 5667 14608 5701
rect 14574 5599 14608 5633
rect 14670 6483 14704 6517
rect 14670 6415 14704 6449
rect 14670 6347 14704 6381
rect 14670 6279 14704 6313
rect 14670 6211 14704 6245
rect 14670 6143 14704 6177
rect 14670 6075 14704 6109
rect 14670 6007 14704 6041
rect 14670 5939 14704 5973
rect 14670 5871 14704 5905
rect 14670 5803 14704 5837
rect 14670 5735 14704 5769
rect 14670 5667 14704 5701
rect 14670 5599 14704 5633
rect 14766 6483 14800 6517
rect 14766 6415 14800 6449
rect 14766 6347 14800 6381
rect 14766 6279 14800 6313
rect 14766 6211 14800 6245
rect 14766 6143 14800 6177
rect 14766 6075 14800 6109
rect 14766 6007 14800 6041
rect 14766 5939 14800 5973
rect 14766 5871 14800 5905
rect 14766 5803 14800 5837
rect 14766 5735 14800 5769
rect 14766 5667 14800 5701
rect 14766 5599 14800 5633
rect 14862 6483 14896 6517
rect 14862 6415 14896 6449
rect 14862 6347 14896 6381
rect 14862 6279 14896 6313
rect 14862 6211 14896 6245
rect 14862 6143 14896 6177
rect 14862 6075 14896 6109
rect 14862 6007 14896 6041
rect 14862 5939 14896 5973
rect 14862 5871 14896 5905
rect 14862 5803 14896 5837
rect 14862 5735 14896 5769
rect 14862 5667 14896 5701
rect 14862 5599 14896 5633
rect 14958 6483 14992 6517
rect 14958 6415 14992 6449
rect 14958 6347 14992 6381
rect 14958 6279 14992 6313
rect 14958 6211 14992 6245
rect 14958 6143 14992 6177
rect 14958 6075 14992 6109
rect 14958 6007 14992 6041
rect 14958 5939 14992 5973
rect 14958 5871 14992 5905
rect 14958 5803 14992 5837
rect 14958 5735 14992 5769
rect 14958 5667 14992 5701
rect 14958 5599 14992 5633
rect 15518 5861 15552 5895
rect 15518 5793 15552 5827
rect 15518 5725 15552 5759
rect 15518 5657 15552 5691
rect 15518 5589 15552 5623
rect -868 5453 -834 5487
rect -868 5385 -834 5419
rect -868 5317 -834 5351
rect -868 5249 -834 5283
rect -868 5181 -834 5215
rect -868 5113 -834 5147
rect -868 5045 -834 5079
rect 15518 5521 15552 5555
rect 15518 5453 15552 5487
rect 15518 5385 15552 5419
rect 15518 5317 15552 5351
rect 15518 5249 15552 5283
rect 15518 5181 15552 5215
rect 15518 5113 15552 5147
rect 15518 5045 15552 5079
rect -868 4977 -834 5011
rect 1484 4869 1518 4903
rect 1484 4801 1518 4835
rect 1484 4733 1518 4767
rect 1484 4665 1518 4699
rect 1484 4597 1518 4631
rect 1484 4529 1518 4563
rect -23586 4367 -23552 4401
rect -23586 4299 -23552 4333
rect -23586 4231 -23552 4265
rect -23586 4163 -23552 4197
rect -23586 4095 -23552 4129
rect -23586 4027 -23552 4061
rect -23586 3959 -23552 3993
rect -23586 3891 -23552 3925
rect -23586 3823 -23552 3857
rect -23586 3755 -23552 3789
rect -23586 3687 -23552 3721
rect -23586 3619 -23552 3653
rect -23586 3551 -23552 3585
rect -23586 3483 -23552 3517
rect -23490 4367 -23456 4401
rect -23490 4299 -23456 4333
rect -23490 4231 -23456 4265
rect -23490 4163 -23456 4197
rect -23490 4095 -23456 4129
rect -23490 4027 -23456 4061
rect -23490 3959 -23456 3993
rect -23490 3891 -23456 3925
rect -23490 3823 -23456 3857
rect -23490 3755 -23456 3789
rect -23490 3687 -23456 3721
rect -23490 3619 -23456 3653
rect -23490 3551 -23456 3585
rect -23490 3483 -23456 3517
rect -23394 4367 -23360 4401
rect -23394 4299 -23360 4333
rect -23394 4231 -23360 4265
rect -23394 4163 -23360 4197
rect -23394 4095 -23360 4129
rect -23394 4027 -23360 4061
rect -23394 3959 -23360 3993
rect -23394 3891 -23360 3925
rect -23394 3823 -23360 3857
rect -23394 3755 -23360 3789
rect -23394 3687 -23360 3721
rect -23394 3619 -23360 3653
rect -23394 3551 -23360 3585
rect -23394 3483 -23360 3517
rect -23298 4367 -23264 4401
rect -23298 4299 -23264 4333
rect -23298 4231 -23264 4265
rect -23298 4163 -23264 4197
rect -23298 4095 -23264 4129
rect -23298 4027 -23264 4061
rect -23298 3959 -23264 3993
rect -23298 3891 -23264 3925
rect -23298 3823 -23264 3857
rect -23298 3755 -23264 3789
rect -23298 3687 -23264 3721
rect -23298 3619 -23264 3653
rect -23298 3551 -23264 3585
rect -23298 3483 -23264 3517
rect -23202 4367 -23168 4401
rect -23202 4299 -23168 4333
rect -23202 4231 -23168 4265
rect -23202 4163 -23168 4197
rect -23202 4095 -23168 4129
rect -23202 4027 -23168 4061
rect -23202 3959 -23168 3993
rect -23202 3891 -23168 3925
rect -23202 3823 -23168 3857
rect -23202 3755 -23168 3789
rect -23202 3687 -23168 3721
rect -23202 3619 -23168 3653
rect -23202 3551 -23168 3585
rect -23202 3483 -23168 3517
rect -23106 4367 -23072 4401
rect -23106 4299 -23072 4333
rect -23106 4231 -23072 4265
rect -23106 4163 -23072 4197
rect -23106 4095 -23072 4129
rect -23106 4027 -23072 4061
rect -23106 3959 -23072 3993
rect -23106 3891 -23072 3925
rect -23106 3823 -23072 3857
rect -23106 3755 -23072 3789
rect -23106 3687 -23072 3721
rect -23106 3619 -23072 3653
rect -23106 3551 -23072 3585
rect -23106 3483 -23072 3517
rect -23010 4367 -22976 4401
rect -23010 4299 -22976 4333
rect -23010 4231 -22976 4265
rect -23010 4163 -22976 4197
rect -23010 4095 -22976 4129
rect -23010 4027 -22976 4061
rect -23010 3959 -22976 3993
rect -23010 3891 -22976 3925
rect -23010 3823 -22976 3857
rect -23010 3755 -22976 3789
rect -23010 3687 -22976 3721
rect -23010 3619 -22976 3653
rect -23010 3551 -22976 3585
rect -23010 3483 -22976 3517
rect -22914 4367 -22880 4401
rect -22914 4299 -22880 4333
rect -22914 4231 -22880 4265
rect -22914 4163 -22880 4197
rect -22914 4095 -22880 4129
rect -22914 4027 -22880 4061
rect -22914 3959 -22880 3993
rect -22914 3891 -22880 3925
rect -22914 3823 -22880 3857
rect -22914 3755 -22880 3789
rect -22914 3687 -22880 3721
rect -22914 3619 -22880 3653
rect -22914 3551 -22880 3585
rect -22914 3483 -22880 3517
rect -22818 4367 -22784 4401
rect -22818 4299 -22784 4333
rect -22818 4231 -22784 4265
rect -22818 4163 -22784 4197
rect -22818 4095 -22784 4129
rect -22818 4027 -22784 4061
rect -22818 3959 -22784 3993
rect -22818 3891 -22784 3925
rect -22818 3823 -22784 3857
rect -22818 3755 -22784 3789
rect -22818 3687 -22784 3721
rect -22818 3619 -22784 3653
rect -22818 3551 -22784 3585
rect -22818 3483 -22784 3517
rect -22722 4367 -22688 4401
rect -22722 4299 -22688 4333
rect -22722 4231 -22688 4265
rect -22722 4163 -22688 4197
rect -22722 4095 -22688 4129
rect -22722 4027 -22688 4061
rect -22722 3959 -22688 3993
rect -22722 3891 -22688 3925
rect -22722 3823 -22688 3857
rect -22722 3755 -22688 3789
rect -22722 3687 -22688 3721
rect -22722 3619 -22688 3653
rect -22722 3551 -22688 3585
rect -22722 3483 -22688 3517
rect -22626 4367 -22592 4401
rect -22626 4299 -22592 4333
rect -22626 4231 -22592 4265
rect -22626 4163 -22592 4197
rect -22626 4095 -22592 4129
rect -22626 4027 -22592 4061
rect -22626 3959 -22592 3993
rect -22626 3891 -22592 3925
rect -22626 3823 -22592 3857
rect -22626 3755 -22592 3789
rect -22626 3687 -22592 3721
rect -22626 3619 -22592 3653
rect -22626 3551 -22592 3585
rect -22626 3483 -22592 3517
rect -22530 4367 -22496 4401
rect -22530 4299 -22496 4333
rect -22530 4231 -22496 4265
rect -22530 4163 -22496 4197
rect -22530 4095 -22496 4129
rect -22530 4027 -22496 4061
rect -22530 3959 -22496 3993
rect -22530 3891 -22496 3925
rect -22530 3823 -22496 3857
rect -22530 3755 -22496 3789
rect -22530 3687 -22496 3721
rect -22530 3619 -22496 3653
rect -22530 3551 -22496 3585
rect -22530 3483 -22496 3517
rect -22434 4367 -22400 4401
rect -22434 4299 -22400 4333
rect -22434 4231 -22400 4265
rect -22434 4163 -22400 4197
rect -22434 4095 -22400 4129
rect -22434 4027 -22400 4061
rect -22434 3959 -22400 3993
rect -22434 3891 -22400 3925
rect -22434 3823 -22400 3857
rect -22434 3755 -22400 3789
rect -22434 3687 -22400 3721
rect -22434 3619 -22400 3653
rect -22434 3551 -22400 3585
rect -22434 3483 -22400 3517
rect -22338 4367 -22304 4401
rect -22338 4299 -22304 4333
rect -22338 4231 -22304 4265
rect -22338 4163 -22304 4197
rect -22338 4095 -22304 4129
rect -22338 4027 -22304 4061
rect -22338 3959 -22304 3993
rect -22338 3891 -22304 3925
rect -22338 3823 -22304 3857
rect -22338 3755 -22304 3789
rect -22338 3687 -22304 3721
rect -22338 3619 -22304 3653
rect -22338 3551 -22304 3585
rect -22338 3483 -22304 3517
rect -22242 4367 -22208 4401
rect -22242 4299 -22208 4333
rect -22242 4231 -22208 4265
rect -22242 4163 -22208 4197
rect -22242 4095 -22208 4129
rect -22242 4027 -22208 4061
rect -22242 3959 -22208 3993
rect -22242 3891 -22208 3925
rect -22242 3823 -22208 3857
rect -22242 3755 -22208 3789
rect -22242 3687 -22208 3721
rect -22242 3619 -22208 3653
rect -22242 3551 -22208 3585
rect -22242 3483 -22208 3517
rect -22146 4367 -22112 4401
rect -22146 4299 -22112 4333
rect -22146 4231 -22112 4265
rect -22146 4163 -22112 4197
rect -22146 4095 -22112 4129
rect -22146 4027 -22112 4061
rect -22146 3959 -22112 3993
rect -22146 3891 -22112 3925
rect -22146 3823 -22112 3857
rect -22146 3755 -22112 3789
rect -22146 3687 -22112 3721
rect -22146 3619 -22112 3653
rect -22146 3551 -22112 3585
rect -22146 3483 -22112 3517
rect -22050 4367 -22016 4401
rect -22050 4299 -22016 4333
rect -22050 4231 -22016 4265
rect -22050 4163 -22016 4197
rect -22050 4095 -22016 4129
rect -22050 4027 -22016 4061
rect -22050 3959 -22016 3993
rect -22050 3891 -22016 3925
rect -22050 3823 -22016 3857
rect -22050 3755 -22016 3789
rect -22050 3687 -22016 3721
rect -22050 3619 -22016 3653
rect -22050 3551 -22016 3585
rect -22050 3483 -22016 3517
rect -21954 4367 -21920 4401
rect -21954 4299 -21920 4333
rect -21954 4231 -21920 4265
rect -21954 4163 -21920 4197
rect -21954 4095 -21920 4129
rect -21954 4027 -21920 4061
rect -21954 3959 -21920 3993
rect -21954 3891 -21920 3925
rect -21954 3823 -21920 3857
rect -21954 3755 -21920 3789
rect -21954 3687 -21920 3721
rect -21954 3619 -21920 3653
rect -21954 3551 -21920 3585
rect -21954 3483 -21920 3517
rect -21858 4367 -21824 4401
rect -21858 4299 -21824 4333
rect -21858 4231 -21824 4265
rect -21858 4163 -21824 4197
rect -21858 4095 -21824 4129
rect -21858 4027 -21824 4061
rect -21858 3959 -21824 3993
rect -21858 3891 -21824 3925
rect -21858 3823 -21824 3857
rect -21858 3755 -21824 3789
rect -21858 3687 -21824 3721
rect -21858 3619 -21824 3653
rect -21858 3551 -21824 3585
rect -21858 3483 -21824 3517
rect -21762 4367 -21728 4401
rect -21762 4299 -21728 4333
rect -21762 4231 -21728 4265
rect -21762 4163 -21728 4197
rect -21762 4095 -21728 4129
rect -21762 4027 -21728 4061
rect -21762 3959 -21728 3993
rect -21762 3891 -21728 3925
rect -21762 3823 -21728 3857
rect -21762 3755 -21728 3789
rect -21762 3687 -21728 3721
rect -21762 3619 -21728 3653
rect -21762 3551 -21728 3585
rect -21762 3483 -21728 3517
rect -21666 4367 -21632 4401
rect -21666 4299 -21632 4333
rect -21666 4231 -21632 4265
rect -21666 4163 -21632 4197
rect -21666 4095 -21632 4129
rect -21666 4027 -21632 4061
rect -21666 3959 -21632 3993
rect -21666 3891 -21632 3925
rect -21666 3823 -21632 3857
rect -21666 3755 -21632 3789
rect -21666 3687 -21632 3721
rect -21666 3619 -21632 3653
rect -21666 3551 -21632 3585
rect -21666 3483 -21632 3517
rect -21442 4373 -21408 4407
rect -21442 4305 -21408 4339
rect -21442 4237 -21408 4271
rect -21442 4169 -21408 4203
rect -21442 4101 -21408 4135
rect -21442 4033 -21408 4067
rect -21442 3965 -21408 3999
rect -21442 3897 -21408 3931
rect -21442 3829 -21408 3863
rect -21442 3761 -21408 3795
rect -21442 3693 -21408 3727
rect -21442 3625 -21408 3659
rect -21442 3557 -21408 3591
rect -21442 3489 -21408 3523
rect -21346 4373 -21312 4407
rect -21346 4305 -21312 4339
rect -21346 4237 -21312 4271
rect -21346 4169 -21312 4203
rect -21346 4101 -21312 4135
rect -21346 4033 -21312 4067
rect -21346 3965 -21312 3999
rect -21346 3897 -21312 3931
rect -21346 3829 -21312 3863
rect -21346 3761 -21312 3795
rect -21346 3693 -21312 3727
rect -21346 3625 -21312 3659
rect -21346 3557 -21312 3591
rect -21346 3489 -21312 3523
rect -21250 4373 -21216 4407
rect -21250 4305 -21216 4339
rect -21250 4237 -21216 4271
rect -21250 4169 -21216 4203
rect -21250 4101 -21216 4135
rect -21250 4033 -21216 4067
rect -21250 3965 -21216 3999
rect -21250 3897 -21216 3931
rect -21250 3829 -21216 3863
rect -21250 3761 -21216 3795
rect -21250 3693 -21216 3727
rect -21250 3625 -21216 3659
rect -21250 3557 -21216 3591
rect -21250 3489 -21216 3523
rect -21154 4373 -21120 4407
rect -21154 4305 -21120 4339
rect -21154 4237 -21120 4271
rect -21154 4169 -21120 4203
rect -21154 4101 -21120 4135
rect -21154 4033 -21120 4067
rect -21154 3965 -21120 3999
rect -21154 3897 -21120 3931
rect -21154 3829 -21120 3863
rect -21154 3761 -21120 3795
rect -21154 3693 -21120 3727
rect -21154 3625 -21120 3659
rect -21154 3557 -21120 3591
rect -21154 3489 -21120 3523
rect -21058 4373 -21024 4407
rect -21058 4305 -21024 4339
rect -21058 4237 -21024 4271
rect -21058 4169 -21024 4203
rect -21058 4101 -21024 4135
rect -21058 4033 -21024 4067
rect -21058 3965 -21024 3999
rect -21058 3897 -21024 3931
rect -21058 3829 -21024 3863
rect -21058 3761 -21024 3795
rect -21058 3693 -21024 3727
rect -21058 3625 -21024 3659
rect -21058 3557 -21024 3591
rect -21058 3489 -21024 3523
rect -20962 4373 -20928 4407
rect -20962 4305 -20928 4339
rect -20962 4237 -20928 4271
rect -20962 4169 -20928 4203
rect -20962 4101 -20928 4135
rect -20962 4033 -20928 4067
rect -20962 3965 -20928 3999
rect -20962 3897 -20928 3931
rect -20962 3829 -20928 3863
rect -20962 3761 -20928 3795
rect -20962 3693 -20928 3727
rect -20962 3625 -20928 3659
rect -20962 3557 -20928 3591
rect -20962 3489 -20928 3523
rect -20866 4373 -20832 4407
rect -20866 4305 -20832 4339
rect -20866 4237 -20832 4271
rect -20866 4169 -20832 4203
rect -20866 4101 -20832 4135
rect -20866 4033 -20832 4067
rect -20866 3965 -20832 3999
rect -20866 3897 -20832 3931
rect -20866 3829 -20832 3863
rect -20866 3761 -20832 3795
rect -20866 3693 -20832 3727
rect -20866 3625 -20832 3659
rect -20866 3557 -20832 3591
rect -20866 3489 -20832 3523
rect -20770 4373 -20736 4407
rect -20770 4305 -20736 4339
rect -20770 4237 -20736 4271
rect -20770 4169 -20736 4203
rect -20770 4101 -20736 4135
rect -20770 4033 -20736 4067
rect -20770 3965 -20736 3999
rect -20770 3897 -20736 3931
rect -20770 3829 -20736 3863
rect -20770 3761 -20736 3795
rect -20770 3693 -20736 3727
rect -20770 3625 -20736 3659
rect -20770 3557 -20736 3591
rect -20770 3489 -20736 3523
rect -20674 4373 -20640 4407
rect -20674 4305 -20640 4339
rect -20674 4237 -20640 4271
rect -20674 4169 -20640 4203
rect -20674 4101 -20640 4135
rect -20674 4033 -20640 4067
rect -20674 3965 -20640 3999
rect -20674 3897 -20640 3931
rect -20674 3829 -20640 3863
rect -20674 3761 -20640 3795
rect -20674 3693 -20640 3727
rect -20674 3625 -20640 3659
rect -20674 3557 -20640 3591
rect -20674 3489 -20640 3523
rect -20578 4373 -20544 4407
rect -20578 4305 -20544 4339
rect -20578 4237 -20544 4271
rect -20578 4169 -20544 4203
rect -20578 4101 -20544 4135
rect -20578 4033 -20544 4067
rect -20578 3965 -20544 3999
rect -20578 3897 -20544 3931
rect -20578 3829 -20544 3863
rect -20578 3761 -20544 3795
rect -20578 3693 -20544 3727
rect -20578 3625 -20544 3659
rect -20578 3557 -20544 3591
rect -20578 3489 -20544 3523
rect -20482 4373 -20448 4407
rect -20482 4305 -20448 4339
rect -20482 4237 -20448 4271
rect -20482 4169 -20448 4203
rect -20482 4101 -20448 4135
rect -20482 4033 -20448 4067
rect -20482 3965 -20448 3999
rect -20482 3897 -20448 3931
rect -20482 3829 -20448 3863
rect -20482 3761 -20448 3795
rect -20482 3693 -20448 3727
rect -20482 3625 -20448 3659
rect -20482 3557 -20448 3591
rect -20482 3489 -20448 3523
rect -20386 4373 -20352 4407
rect -20386 4305 -20352 4339
rect -20386 4237 -20352 4271
rect -20386 4169 -20352 4203
rect -20386 4101 -20352 4135
rect -20386 4033 -20352 4067
rect -20386 3965 -20352 3999
rect -20386 3897 -20352 3931
rect -20386 3829 -20352 3863
rect -20386 3761 -20352 3795
rect -20386 3693 -20352 3727
rect -20386 3625 -20352 3659
rect -20386 3557 -20352 3591
rect -20386 3489 -20352 3523
rect -20290 4373 -20256 4407
rect -20290 4305 -20256 4339
rect -20290 4237 -20256 4271
rect -20290 4169 -20256 4203
rect -20290 4101 -20256 4135
rect -20290 4033 -20256 4067
rect -20290 3965 -20256 3999
rect -20290 3897 -20256 3931
rect -20290 3829 -20256 3863
rect -20290 3761 -20256 3795
rect -20290 3693 -20256 3727
rect -20290 3625 -20256 3659
rect -20290 3557 -20256 3591
rect -20290 3489 -20256 3523
rect -20194 4373 -20160 4407
rect -20194 4305 -20160 4339
rect -20194 4237 -20160 4271
rect -20194 4169 -20160 4203
rect -20194 4101 -20160 4135
rect -20194 4033 -20160 4067
rect -20194 3965 -20160 3999
rect -20194 3897 -20160 3931
rect -20194 3829 -20160 3863
rect -20194 3761 -20160 3795
rect -20194 3693 -20160 3727
rect -20194 3625 -20160 3659
rect -20194 3557 -20160 3591
rect -20194 3489 -20160 3523
rect -20098 4373 -20064 4407
rect -20098 4305 -20064 4339
rect -20098 4237 -20064 4271
rect -20098 4169 -20064 4203
rect -20098 4101 -20064 4135
rect -20098 4033 -20064 4067
rect -20098 3965 -20064 3999
rect -20098 3897 -20064 3931
rect -20098 3829 -20064 3863
rect -20098 3761 -20064 3795
rect -20098 3693 -20064 3727
rect -20098 3625 -20064 3659
rect -20098 3557 -20064 3591
rect -20098 3489 -20064 3523
rect -20002 4373 -19968 4407
rect -20002 4305 -19968 4339
rect -20002 4237 -19968 4271
rect -20002 4169 -19968 4203
rect -20002 4101 -19968 4135
rect -20002 4033 -19968 4067
rect -20002 3965 -19968 3999
rect -20002 3897 -19968 3931
rect -20002 3829 -19968 3863
rect -20002 3761 -19968 3795
rect -20002 3693 -19968 3727
rect -20002 3625 -19968 3659
rect -20002 3557 -19968 3591
rect -20002 3489 -19968 3523
rect -19758 4379 -19724 4413
rect -19758 4311 -19724 4345
rect -19758 4243 -19724 4277
rect -19758 4175 -19724 4209
rect -19758 4107 -19724 4141
rect -19758 4039 -19724 4073
rect -19758 3971 -19724 4005
rect -19758 3903 -19724 3937
rect -19758 3835 -19724 3869
rect -19758 3767 -19724 3801
rect -19758 3699 -19724 3733
rect -19758 3631 -19724 3665
rect -19758 3563 -19724 3597
rect -19758 3495 -19724 3529
rect -19662 4379 -19628 4413
rect -19662 4311 -19628 4345
rect -19662 4243 -19628 4277
rect -19662 4175 -19628 4209
rect -19662 4107 -19628 4141
rect -19662 4039 -19628 4073
rect -19662 3971 -19628 4005
rect -19662 3903 -19628 3937
rect -19662 3835 -19628 3869
rect -19662 3767 -19628 3801
rect -19662 3699 -19628 3733
rect -19662 3631 -19628 3665
rect -19662 3563 -19628 3597
rect -19662 3495 -19628 3529
rect -19566 4379 -19532 4413
rect -19566 4311 -19532 4345
rect -19566 4243 -19532 4277
rect -19566 4175 -19532 4209
rect -19566 4107 -19532 4141
rect -19566 4039 -19532 4073
rect -19566 3971 -19532 4005
rect -19566 3903 -19532 3937
rect -19566 3835 -19532 3869
rect -19566 3767 -19532 3801
rect -19566 3699 -19532 3733
rect -19566 3631 -19532 3665
rect -19566 3563 -19532 3597
rect -19566 3495 -19532 3529
rect -19470 4379 -19436 4413
rect -19470 4311 -19436 4345
rect -19470 4243 -19436 4277
rect -19470 4175 -19436 4209
rect -19470 4107 -19436 4141
rect -19470 4039 -19436 4073
rect -19470 3971 -19436 4005
rect -19470 3903 -19436 3937
rect -19470 3835 -19436 3869
rect -19470 3767 -19436 3801
rect -19470 3699 -19436 3733
rect -19470 3631 -19436 3665
rect -19470 3563 -19436 3597
rect -19470 3495 -19436 3529
rect -19374 4379 -19340 4413
rect -19374 4311 -19340 4345
rect -19374 4243 -19340 4277
rect -19374 4175 -19340 4209
rect -19374 4107 -19340 4141
rect -19374 4039 -19340 4073
rect -19374 3971 -19340 4005
rect -19374 3903 -19340 3937
rect -19374 3835 -19340 3869
rect -19374 3767 -19340 3801
rect -19374 3699 -19340 3733
rect -19374 3631 -19340 3665
rect -19374 3563 -19340 3597
rect -19374 3495 -19340 3529
rect -19278 4379 -19244 4413
rect -19278 4311 -19244 4345
rect -19278 4243 -19244 4277
rect -19278 4175 -19244 4209
rect -19278 4107 -19244 4141
rect -19278 4039 -19244 4073
rect -19278 3971 -19244 4005
rect -19278 3903 -19244 3937
rect -19278 3835 -19244 3869
rect -19278 3767 -19244 3801
rect -19278 3699 -19244 3733
rect -19278 3631 -19244 3665
rect -19278 3563 -19244 3597
rect -19278 3495 -19244 3529
rect -19182 4379 -19148 4413
rect -19182 4311 -19148 4345
rect -19182 4243 -19148 4277
rect -19182 4175 -19148 4209
rect -19182 4107 -19148 4141
rect -19182 4039 -19148 4073
rect -19182 3971 -19148 4005
rect -19182 3903 -19148 3937
rect -19182 3835 -19148 3869
rect -19182 3767 -19148 3801
rect -19182 3699 -19148 3733
rect -19182 3631 -19148 3665
rect -19182 3563 -19148 3597
rect -19182 3495 -19148 3529
rect -19086 4379 -19052 4413
rect -19086 4311 -19052 4345
rect -19086 4243 -19052 4277
rect -19086 4175 -19052 4209
rect -19086 4107 -19052 4141
rect -19086 4039 -19052 4073
rect -19086 3971 -19052 4005
rect -19086 3903 -19052 3937
rect -19086 3835 -19052 3869
rect -19086 3767 -19052 3801
rect -19086 3699 -19052 3733
rect -19086 3631 -19052 3665
rect -19086 3563 -19052 3597
rect -19086 3495 -19052 3529
rect -18990 4379 -18956 4413
rect -18990 4311 -18956 4345
rect -18990 4243 -18956 4277
rect -18990 4175 -18956 4209
rect -18990 4107 -18956 4141
rect -18990 4039 -18956 4073
rect -18990 3971 -18956 4005
rect -18990 3903 -18956 3937
rect -18990 3835 -18956 3869
rect -18990 3767 -18956 3801
rect -18990 3699 -18956 3733
rect -18990 3631 -18956 3665
rect -18990 3563 -18956 3597
rect -18990 3495 -18956 3529
rect -18894 4379 -18860 4413
rect -18894 4311 -18860 4345
rect -18894 4243 -18860 4277
rect -18894 4175 -18860 4209
rect -18894 4107 -18860 4141
rect -18894 4039 -18860 4073
rect -18894 3971 -18860 4005
rect -18894 3903 -18860 3937
rect -18894 3835 -18860 3869
rect -18894 3767 -18860 3801
rect -18894 3699 -18860 3733
rect -18894 3631 -18860 3665
rect -18894 3563 -18860 3597
rect -18894 3495 -18860 3529
rect -18798 4379 -18764 4413
rect -18798 4311 -18764 4345
rect -18798 4243 -18764 4277
rect -18798 4175 -18764 4209
rect -18798 4107 -18764 4141
rect -18798 4039 -18764 4073
rect -18798 3971 -18764 4005
rect -18798 3903 -18764 3937
rect -18798 3835 -18764 3869
rect -18798 3767 -18764 3801
rect -18798 3699 -18764 3733
rect -18798 3631 -18764 3665
rect -18798 3563 -18764 3597
rect -18798 3495 -18764 3529
rect -18590 4381 -18556 4415
rect -18590 4313 -18556 4347
rect -18590 4245 -18556 4279
rect -18590 4177 -18556 4211
rect -18590 4109 -18556 4143
rect -18590 4041 -18556 4075
rect -18590 3973 -18556 4007
rect -18590 3905 -18556 3939
rect -18590 3837 -18556 3871
rect -18590 3769 -18556 3803
rect -18590 3701 -18556 3735
rect -18590 3633 -18556 3667
rect -18590 3565 -18556 3599
rect -18590 3497 -18556 3531
rect -18494 4381 -18460 4415
rect -18494 4313 -18460 4347
rect -18494 4245 -18460 4279
rect -18494 4177 -18460 4211
rect -18494 4109 -18460 4143
rect -18494 4041 -18460 4075
rect -18494 3973 -18460 4007
rect -18494 3905 -18460 3939
rect -18494 3837 -18460 3871
rect -18494 3769 -18460 3803
rect -18494 3701 -18460 3735
rect -18494 3633 -18460 3667
rect -18494 3565 -18460 3599
rect -18494 3497 -18460 3531
rect -18398 4381 -18364 4415
rect -18398 4313 -18364 4347
rect -18398 4245 -18364 4279
rect -18398 4177 -18364 4211
rect -18398 4109 -18364 4143
rect -18398 4041 -18364 4075
rect -18398 3973 -18364 4007
rect -18398 3905 -18364 3939
rect -18398 3837 -18364 3871
rect -18398 3769 -18364 3803
rect -18398 3701 -18364 3735
rect -18398 3633 -18364 3667
rect -18398 3565 -18364 3599
rect -18398 3497 -18364 3531
rect -18302 4381 -18268 4415
rect -18302 4313 -18268 4347
rect -18302 4245 -18268 4279
rect -18302 4177 -18268 4211
rect -18302 4109 -18268 4143
rect -18302 4041 -18268 4075
rect -18302 3973 -18268 4007
rect -18302 3905 -18268 3939
rect -18302 3837 -18268 3871
rect -18302 3769 -18268 3803
rect -18302 3701 -18268 3735
rect -18302 3633 -18268 3667
rect -18302 3565 -18268 3599
rect -18302 3497 -18268 3531
rect -18206 4381 -18172 4415
rect -18206 4313 -18172 4347
rect -18206 4245 -18172 4279
rect -18206 4177 -18172 4211
rect -18206 4109 -18172 4143
rect -18206 4041 -18172 4075
rect -18206 3973 -18172 4007
rect -18206 3905 -18172 3939
rect -18206 3837 -18172 3871
rect -18206 3769 -18172 3803
rect -18206 3701 -18172 3735
rect -18206 3633 -18172 3667
rect -18206 3565 -18172 3599
rect -18206 3497 -18172 3531
rect -18110 4381 -18076 4415
rect -18110 4313 -18076 4347
rect -18110 4245 -18076 4279
rect -18110 4177 -18076 4211
rect -18110 4109 -18076 4143
rect -18110 4041 -18076 4075
rect -18110 3973 -18076 4007
rect -18110 3905 -18076 3939
rect -18110 3837 -18076 3871
rect -18110 3769 -18076 3803
rect -18110 3701 -18076 3735
rect -18110 3633 -18076 3667
rect -18110 3565 -18076 3599
rect -18110 3497 -18076 3531
rect -16756 4379 -16722 4413
rect -16756 4311 -16722 4345
rect -16756 4243 -16722 4277
rect -16756 4175 -16722 4209
rect -16756 4107 -16722 4141
rect -16756 4039 -16722 4073
rect -16756 3971 -16722 4005
rect -16756 3903 -16722 3937
rect -16756 3835 -16722 3869
rect -16756 3767 -16722 3801
rect -16756 3699 -16722 3733
rect -16756 3631 -16722 3665
rect -16756 3563 -16722 3597
rect -16756 3495 -16722 3529
rect -16660 4379 -16626 4413
rect -16660 4311 -16626 4345
rect -16660 4243 -16626 4277
rect -16660 4175 -16626 4209
rect -16660 4107 -16626 4141
rect -16660 4039 -16626 4073
rect -16660 3971 -16626 4005
rect -16660 3903 -16626 3937
rect -16660 3835 -16626 3869
rect -16660 3767 -16626 3801
rect -16660 3699 -16626 3733
rect -16660 3631 -16626 3665
rect -16660 3563 -16626 3597
rect -16660 3495 -16626 3529
rect -16564 4379 -16530 4413
rect -16564 4311 -16530 4345
rect -16564 4243 -16530 4277
rect -16564 4175 -16530 4209
rect -16564 4107 -16530 4141
rect -16564 4039 -16530 4073
rect -16564 3971 -16530 4005
rect -16564 3903 -16530 3937
rect -16564 3835 -16530 3869
rect -16564 3767 -16530 3801
rect -16564 3699 -16530 3733
rect -16564 3631 -16530 3665
rect -16564 3563 -16530 3597
rect -16564 3495 -16530 3529
rect -16468 4379 -16434 4413
rect -16468 4311 -16434 4345
rect -16468 4243 -16434 4277
rect -16468 4175 -16434 4209
rect -16468 4107 -16434 4141
rect -16468 4039 -16434 4073
rect -16468 3971 -16434 4005
rect -16468 3903 -16434 3937
rect -16468 3835 -16434 3869
rect -16468 3767 -16434 3801
rect -16468 3699 -16434 3733
rect -16468 3631 -16434 3665
rect -16468 3563 -16434 3597
rect -16468 3495 -16434 3529
rect -16372 4379 -16338 4413
rect -16372 4311 -16338 4345
rect -16372 4243 -16338 4277
rect -16372 4175 -16338 4209
rect -16372 4107 -16338 4141
rect -16372 4039 -16338 4073
rect -16372 3971 -16338 4005
rect -16372 3903 -16338 3937
rect -16372 3835 -16338 3869
rect -16372 3767 -16338 3801
rect -16372 3699 -16338 3733
rect -16372 3631 -16338 3665
rect -16372 3563 -16338 3597
rect -16372 3495 -16338 3529
rect -16276 4379 -16242 4413
rect -16276 4311 -16242 4345
rect -16276 4243 -16242 4277
rect -16276 4175 -16242 4209
rect -16276 4107 -16242 4141
rect -16276 4039 -16242 4073
rect -16276 3971 -16242 4005
rect -16276 3903 -16242 3937
rect -16276 3835 -16242 3869
rect -16276 3767 -16242 3801
rect -16276 3699 -16242 3733
rect -16276 3631 -16242 3665
rect -16276 3563 -16242 3597
rect -16276 3495 -16242 3529
rect -16180 4379 -16146 4413
rect -16180 4311 -16146 4345
rect -16180 4243 -16146 4277
rect -16180 4175 -16146 4209
rect -16180 4107 -16146 4141
rect -16180 4039 -16146 4073
rect -16180 3971 -16146 4005
rect -16180 3903 -16146 3937
rect -16180 3835 -16146 3869
rect -16180 3767 -16146 3801
rect -16180 3699 -16146 3733
rect -16180 3631 -16146 3665
rect -16180 3563 -16146 3597
rect -16180 3495 -16146 3529
rect -16084 4379 -16050 4413
rect -16084 4311 -16050 4345
rect -16084 4243 -16050 4277
rect -16084 4175 -16050 4209
rect -16084 4107 -16050 4141
rect -16084 4039 -16050 4073
rect -16084 3971 -16050 4005
rect -16084 3903 -16050 3937
rect -16084 3835 -16050 3869
rect -16084 3767 -16050 3801
rect -16084 3699 -16050 3733
rect -16084 3631 -16050 3665
rect -16084 3563 -16050 3597
rect -16084 3495 -16050 3529
rect -15988 4379 -15954 4413
rect -15988 4311 -15954 4345
rect -15988 4243 -15954 4277
rect -15988 4175 -15954 4209
rect -15988 4107 -15954 4141
rect -15988 4039 -15954 4073
rect -15988 3971 -15954 4005
rect -15988 3903 -15954 3937
rect -15988 3835 -15954 3869
rect -15988 3767 -15954 3801
rect -15988 3699 -15954 3733
rect -15988 3631 -15954 3665
rect -15988 3563 -15954 3597
rect -15988 3495 -15954 3529
rect -15892 4379 -15858 4413
rect -15892 4311 -15858 4345
rect -15892 4243 -15858 4277
rect -15892 4175 -15858 4209
rect -15892 4107 -15858 4141
rect -15892 4039 -15858 4073
rect -15892 3971 -15858 4005
rect -15892 3903 -15858 3937
rect -15892 3835 -15858 3869
rect -15892 3767 -15858 3801
rect -15892 3699 -15858 3733
rect -15892 3631 -15858 3665
rect -15892 3563 -15858 3597
rect -15892 3495 -15858 3529
rect -15796 4379 -15762 4413
rect -15796 4311 -15762 4345
rect -15796 4243 -15762 4277
rect -15796 4175 -15762 4209
rect -15796 4107 -15762 4141
rect -15796 4039 -15762 4073
rect -15796 3971 -15762 4005
rect -15796 3903 -15762 3937
rect -15796 3835 -15762 3869
rect -15796 3767 -15762 3801
rect -15796 3699 -15762 3733
rect -15796 3631 -15762 3665
rect -15796 3563 -15762 3597
rect -15796 3495 -15762 3529
rect -15700 4379 -15666 4413
rect -15700 4311 -15666 4345
rect -15700 4243 -15666 4277
rect -15700 4175 -15666 4209
rect -15700 4107 -15666 4141
rect -15700 4039 -15666 4073
rect -15700 3971 -15666 4005
rect -15700 3903 -15666 3937
rect -15700 3835 -15666 3869
rect -15700 3767 -15666 3801
rect -15700 3699 -15666 3733
rect -15700 3631 -15666 3665
rect -15700 3563 -15666 3597
rect -15700 3495 -15666 3529
rect -15604 4379 -15570 4413
rect -15604 4311 -15570 4345
rect -15604 4243 -15570 4277
rect -15604 4175 -15570 4209
rect -15604 4107 -15570 4141
rect -15604 4039 -15570 4073
rect -15604 3971 -15570 4005
rect -15604 3903 -15570 3937
rect -15604 3835 -15570 3869
rect -15604 3767 -15570 3801
rect -15604 3699 -15570 3733
rect -15604 3631 -15570 3665
rect -15604 3563 -15570 3597
rect -15604 3495 -15570 3529
rect -15508 4379 -15474 4413
rect -15508 4311 -15474 4345
rect -15508 4243 -15474 4277
rect -15508 4175 -15474 4209
rect -15508 4107 -15474 4141
rect -15508 4039 -15474 4073
rect -15508 3971 -15474 4005
rect -15508 3903 -15474 3937
rect -15508 3835 -15474 3869
rect -15508 3767 -15474 3801
rect -15508 3699 -15474 3733
rect -15508 3631 -15474 3665
rect -15508 3563 -15474 3597
rect -15508 3495 -15474 3529
rect -15412 4379 -15378 4413
rect -15412 4311 -15378 4345
rect -15412 4243 -15378 4277
rect -15412 4175 -15378 4209
rect -15412 4107 -15378 4141
rect -15412 4039 -15378 4073
rect -15412 3971 -15378 4005
rect -15412 3903 -15378 3937
rect -15412 3835 -15378 3869
rect -15412 3767 -15378 3801
rect -15412 3699 -15378 3733
rect -15412 3631 -15378 3665
rect -15412 3563 -15378 3597
rect -15412 3495 -15378 3529
rect -15316 4379 -15282 4413
rect -15316 4311 -15282 4345
rect -15316 4243 -15282 4277
rect -15316 4175 -15282 4209
rect -15316 4107 -15282 4141
rect -15316 4039 -15282 4073
rect -15316 3971 -15282 4005
rect -15316 3903 -15282 3937
rect -15316 3835 -15282 3869
rect -15316 3767 -15282 3801
rect -15316 3699 -15282 3733
rect -15316 3631 -15282 3665
rect -15316 3563 -15282 3597
rect -15316 3495 -15282 3529
rect -15220 4379 -15186 4413
rect -15220 4311 -15186 4345
rect -15220 4243 -15186 4277
rect -15220 4175 -15186 4209
rect -15220 4107 -15186 4141
rect -15220 4039 -15186 4073
rect -15220 3971 -15186 4005
rect -15220 3903 -15186 3937
rect -15220 3835 -15186 3869
rect -15220 3767 -15186 3801
rect -15220 3699 -15186 3733
rect -15220 3631 -15186 3665
rect -15220 3563 -15186 3597
rect -15220 3495 -15186 3529
rect -15124 4379 -15090 4413
rect -15124 4311 -15090 4345
rect -15124 4243 -15090 4277
rect -15124 4175 -15090 4209
rect -15124 4107 -15090 4141
rect -15124 4039 -15090 4073
rect -15124 3971 -15090 4005
rect -15124 3903 -15090 3937
rect -15124 3835 -15090 3869
rect -15124 3767 -15090 3801
rect -15124 3699 -15090 3733
rect -15124 3631 -15090 3665
rect -15124 3563 -15090 3597
rect -15124 3495 -15090 3529
rect -15028 4379 -14994 4413
rect -15028 4311 -14994 4345
rect -15028 4243 -14994 4277
rect -15028 4175 -14994 4209
rect -15028 4107 -14994 4141
rect -15028 4039 -14994 4073
rect -15028 3971 -14994 4005
rect -15028 3903 -14994 3937
rect -15028 3835 -14994 3869
rect -15028 3767 -14994 3801
rect -15028 3699 -14994 3733
rect -15028 3631 -14994 3665
rect -15028 3563 -14994 3597
rect -15028 3495 -14994 3529
rect -14932 4379 -14898 4413
rect -14932 4311 -14898 4345
rect -14932 4243 -14898 4277
rect -14932 4175 -14898 4209
rect -14932 4107 -14898 4141
rect -14932 4039 -14898 4073
rect -14932 3971 -14898 4005
rect -14932 3903 -14898 3937
rect -14932 3835 -14898 3869
rect -14932 3767 -14898 3801
rect -14932 3699 -14898 3733
rect -14932 3631 -14898 3665
rect -14932 3563 -14898 3597
rect -14932 3495 -14898 3529
rect -14836 4379 -14802 4413
rect -14836 4311 -14802 4345
rect -14836 4243 -14802 4277
rect -14836 4175 -14802 4209
rect -14836 4107 -14802 4141
rect -14836 4039 -14802 4073
rect -14836 3971 -14802 4005
rect -14836 3903 -14802 3937
rect -14836 3835 -14802 3869
rect -14836 3767 -14802 3801
rect -14836 3699 -14802 3733
rect -14836 3631 -14802 3665
rect -14836 3563 -14802 3597
rect -14836 3495 -14802 3529
rect -14612 4385 -14578 4419
rect -14612 4317 -14578 4351
rect -14612 4249 -14578 4283
rect -14612 4181 -14578 4215
rect -14612 4113 -14578 4147
rect -14612 4045 -14578 4079
rect -14612 3977 -14578 4011
rect -14612 3909 -14578 3943
rect -14612 3841 -14578 3875
rect -14612 3773 -14578 3807
rect -14612 3705 -14578 3739
rect -14612 3637 -14578 3671
rect -14612 3569 -14578 3603
rect -14612 3501 -14578 3535
rect -14516 4385 -14482 4419
rect -14516 4317 -14482 4351
rect -14516 4249 -14482 4283
rect -14516 4181 -14482 4215
rect -14516 4113 -14482 4147
rect -14516 4045 -14482 4079
rect -14516 3977 -14482 4011
rect -14516 3909 -14482 3943
rect -14516 3841 -14482 3875
rect -14516 3773 -14482 3807
rect -14516 3705 -14482 3739
rect -14516 3637 -14482 3671
rect -14516 3569 -14482 3603
rect -14516 3501 -14482 3535
rect -14420 4385 -14386 4419
rect -14420 4317 -14386 4351
rect -14420 4249 -14386 4283
rect -14420 4181 -14386 4215
rect -14420 4113 -14386 4147
rect -14420 4045 -14386 4079
rect -14420 3977 -14386 4011
rect -14420 3909 -14386 3943
rect -14420 3841 -14386 3875
rect -14420 3773 -14386 3807
rect -14420 3705 -14386 3739
rect -14420 3637 -14386 3671
rect -14420 3569 -14386 3603
rect -14420 3501 -14386 3535
rect -14324 4385 -14290 4419
rect -14324 4317 -14290 4351
rect -14324 4249 -14290 4283
rect -14324 4181 -14290 4215
rect -14324 4113 -14290 4147
rect -14324 4045 -14290 4079
rect -14324 3977 -14290 4011
rect -14324 3909 -14290 3943
rect -14324 3841 -14290 3875
rect -14324 3773 -14290 3807
rect -14324 3705 -14290 3739
rect -14324 3637 -14290 3671
rect -14324 3569 -14290 3603
rect -14324 3501 -14290 3535
rect -14228 4385 -14194 4419
rect -14228 4317 -14194 4351
rect -14228 4249 -14194 4283
rect -14228 4181 -14194 4215
rect -14228 4113 -14194 4147
rect -14228 4045 -14194 4079
rect -14228 3977 -14194 4011
rect -14228 3909 -14194 3943
rect -14228 3841 -14194 3875
rect -14228 3773 -14194 3807
rect -14228 3705 -14194 3739
rect -14228 3637 -14194 3671
rect -14228 3569 -14194 3603
rect -14228 3501 -14194 3535
rect -14132 4385 -14098 4419
rect -14132 4317 -14098 4351
rect -14132 4249 -14098 4283
rect -14132 4181 -14098 4215
rect -14132 4113 -14098 4147
rect -14132 4045 -14098 4079
rect -14132 3977 -14098 4011
rect -14132 3909 -14098 3943
rect -14132 3841 -14098 3875
rect -14132 3773 -14098 3807
rect -14132 3705 -14098 3739
rect -14132 3637 -14098 3671
rect -14132 3569 -14098 3603
rect -14132 3501 -14098 3535
rect -14036 4385 -14002 4419
rect -14036 4317 -14002 4351
rect -14036 4249 -14002 4283
rect -14036 4181 -14002 4215
rect -14036 4113 -14002 4147
rect -14036 4045 -14002 4079
rect -14036 3977 -14002 4011
rect -14036 3909 -14002 3943
rect -14036 3841 -14002 3875
rect -14036 3773 -14002 3807
rect -14036 3705 -14002 3739
rect -14036 3637 -14002 3671
rect -14036 3569 -14002 3603
rect -14036 3501 -14002 3535
rect -13940 4385 -13906 4419
rect -13940 4317 -13906 4351
rect -13940 4249 -13906 4283
rect -13940 4181 -13906 4215
rect -13940 4113 -13906 4147
rect -13940 4045 -13906 4079
rect -13940 3977 -13906 4011
rect -13940 3909 -13906 3943
rect -13940 3841 -13906 3875
rect -13940 3773 -13906 3807
rect -13940 3705 -13906 3739
rect -13940 3637 -13906 3671
rect -13940 3569 -13906 3603
rect -13940 3501 -13906 3535
rect -13844 4385 -13810 4419
rect -13844 4317 -13810 4351
rect -13844 4249 -13810 4283
rect -13844 4181 -13810 4215
rect -13844 4113 -13810 4147
rect -13844 4045 -13810 4079
rect -13844 3977 -13810 4011
rect -13844 3909 -13810 3943
rect -13844 3841 -13810 3875
rect -13844 3773 -13810 3807
rect -13844 3705 -13810 3739
rect -13844 3637 -13810 3671
rect -13844 3569 -13810 3603
rect -13844 3501 -13810 3535
rect -13748 4385 -13714 4419
rect -13748 4317 -13714 4351
rect -13748 4249 -13714 4283
rect -13748 4181 -13714 4215
rect -13748 4113 -13714 4147
rect -13748 4045 -13714 4079
rect -13748 3977 -13714 4011
rect -13748 3909 -13714 3943
rect -13748 3841 -13714 3875
rect -13748 3773 -13714 3807
rect -13748 3705 -13714 3739
rect -13748 3637 -13714 3671
rect -13748 3569 -13714 3603
rect -13748 3501 -13714 3535
rect -13652 4385 -13618 4419
rect -13652 4317 -13618 4351
rect -13652 4249 -13618 4283
rect -13652 4181 -13618 4215
rect -13652 4113 -13618 4147
rect -13652 4045 -13618 4079
rect -13652 3977 -13618 4011
rect -13652 3909 -13618 3943
rect -13652 3841 -13618 3875
rect -13652 3773 -13618 3807
rect -13652 3705 -13618 3739
rect -13652 3637 -13618 3671
rect -13652 3569 -13618 3603
rect -13652 3501 -13618 3535
rect -13556 4385 -13522 4419
rect -13556 4317 -13522 4351
rect -13556 4249 -13522 4283
rect -13556 4181 -13522 4215
rect -13556 4113 -13522 4147
rect -13556 4045 -13522 4079
rect -13556 3977 -13522 4011
rect -13556 3909 -13522 3943
rect -13556 3841 -13522 3875
rect -13556 3773 -13522 3807
rect -13556 3705 -13522 3739
rect -13556 3637 -13522 3671
rect -13556 3569 -13522 3603
rect -13556 3501 -13522 3535
rect -13460 4385 -13426 4419
rect -13460 4317 -13426 4351
rect -13460 4249 -13426 4283
rect -13460 4181 -13426 4215
rect -13460 4113 -13426 4147
rect -13460 4045 -13426 4079
rect -13460 3977 -13426 4011
rect -13460 3909 -13426 3943
rect -13460 3841 -13426 3875
rect -13460 3773 -13426 3807
rect -13460 3705 -13426 3739
rect -13460 3637 -13426 3671
rect -13460 3569 -13426 3603
rect -13460 3501 -13426 3535
rect -13364 4385 -13330 4419
rect -13364 4317 -13330 4351
rect -13364 4249 -13330 4283
rect -13364 4181 -13330 4215
rect -13364 4113 -13330 4147
rect -13364 4045 -13330 4079
rect -13364 3977 -13330 4011
rect -13364 3909 -13330 3943
rect -13364 3841 -13330 3875
rect -13364 3773 -13330 3807
rect -13364 3705 -13330 3739
rect -13364 3637 -13330 3671
rect -13364 3569 -13330 3603
rect -13364 3501 -13330 3535
rect -13268 4385 -13234 4419
rect -13268 4317 -13234 4351
rect -13268 4249 -13234 4283
rect -13268 4181 -13234 4215
rect -13268 4113 -13234 4147
rect -13268 4045 -13234 4079
rect -13268 3977 -13234 4011
rect -13268 3909 -13234 3943
rect -13268 3841 -13234 3875
rect -13268 3773 -13234 3807
rect -13268 3705 -13234 3739
rect -13268 3637 -13234 3671
rect -13268 3569 -13234 3603
rect -13268 3501 -13234 3535
rect -13172 4385 -13138 4419
rect -13172 4317 -13138 4351
rect -13172 4249 -13138 4283
rect -13172 4181 -13138 4215
rect -13172 4113 -13138 4147
rect -13172 4045 -13138 4079
rect -13172 3977 -13138 4011
rect -13172 3909 -13138 3943
rect -13172 3841 -13138 3875
rect -13172 3773 -13138 3807
rect -13172 3705 -13138 3739
rect -13172 3637 -13138 3671
rect -13172 3569 -13138 3603
rect -13172 3501 -13138 3535
rect -12928 4391 -12894 4425
rect -12928 4323 -12894 4357
rect -12928 4255 -12894 4289
rect -12928 4187 -12894 4221
rect -12928 4119 -12894 4153
rect -12928 4051 -12894 4085
rect -12928 3983 -12894 4017
rect -12928 3915 -12894 3949
rect -12928 3847 -12894 3881
rect -12928 3779 -12894 3813
rect -12928 3711 -12894 3745
rect -12928 3643 -12894 3677
rect -12928 3575 -12894 3609
rect -12928 3507 -12894 3541
rect -12832 4391 -12798 4425
rect -12832 4323 -12798 4357
rect -12832 4255 -12798 4289
rect -12832 4187 -12798 4221
rect -12832 4119 -12798 4153
rect -12832 4051 -12798 4085
rect -12832 3983 -12798 4017
rect -12832 3915 -12798 3949
rect -12832 3847 -12798 3881
rect -12832 3779 -12798 3813
rect -12832 3711 -12798 3745
rect -12832 3643 -12798 3677
rect -12832 3575 -12798 3609
rect -12832 3507 -12798 3541
rect -12736 4391 -12702 4425
rect -12736 4323 -12702 4357
rect -12736 4255 -12702 4289
rect -12736 4187 -12702 4221
rect -12736 4119 -12702 4153
rect -12736 4051 -12702 4085
rect -12736 3983 -12702 4017
rect -12736 3915 -12702 3949
rect -12736 3847 -12702 3881
rect -12736 3779 -12702 3813
rect -12736 3711 -12702 3745
rect -12736 3643 -12702 3677
rect -12736 3575 -12702 3609
rect -12736 3507 -12702 3541
rect -12640 4391 -12606 4425
rect -12640 4323 -12606 4357
rect -12640 4255 -12606 4289
rect -12640 4187 -12606 4221
rect -12640 4119 -12606 4153
rect -12640 4051 -12606 4085
rect -12640 3983 -12606 4017
rect -12640 3915 -12606 3949
rect -12640 3847 -12606 3881
rect -12640 3779 -12606 3813
rect -12640 3711 -12606 3745
rect -12640 3643 -12606 3677
rect -12640 3575 -12606 3609
rect -12640 3507 -12606 3541
rect -12544 4391 -12510 4425
rect -12544 4323 -12510 4357
rect -12544 4255 -12510 4289
rect -12544 4187 -12510 4221
rect -12544 4119 -12510 4153
rect -12544 4051 -12510 4085
rect -12544 3983 -12510 4017
rect -12544 3915 -12510 3949
rect -12544 3847 -12510 3881
rect -12544 3779 -12510 3813
rect -12544 3711 -12510 3745
rect -12544 3643 -12510 3677
rect -12544 3575 -12510 3609
rect -12544 3507 -12510 3541
rect -12448 4391 -12414 4425
rect -12448 4323 -12414 4357
rect -12448 4255 -12414 4289
rect -12448 4187 -12414 4221
rect -12448 4119 -12414 4153
rect -12448 4051 -12414 4085
rect -12448 3983 -12414 4017
rect -12448 3915 -12414 3949
rect -12448 3847 -12414 3881
rect -12448 3779 -12414 3813
rect -12448 3711 -12414 3745
rect -12448 3643 -12414 3677
rect -12448 3575 -12414 3609
rect -12448 3507 -12414 3541
rect -12352 4391 -12318 4425
rect -12352 4323 -12318 4357
rect -12352 4255 -12318 4289
rect -12352 4187 -12318 4221
rect -12352 4119 -12318 4153
rect -12352 4051 -12318 4085
rect -12352 3983 -12318 4017
rect -12352 3915 -12318 3949
rect -12352 3847 -12318 3881
rect -12352 3779 -12318 3813
rect -12352 3711 -12318 3745
rect -12352 3643 -12318 3677
rect -12352 3575 -12318 3609
rect -12352 3507 -12318 3541
rect -12256 4391 -12222 4425
rect -12256 4323 -12222 4357
rect -12256 4255 -12222 4289
rect -12256 4187 -12222 4221
rect -12256 4119 -12222 4153
rect -12256 4051 -12222 4085
rect -12256 3983 -12222 4017
rect -12256 3915 -12222 3949
rect -12256 3847 -12222 3881
rect -12256 3779 -12222 3813
rect -12256 3711 -12222 3745
rect -12256 3643 -12222 3677
rect -12256 3575 -12222 3609
rect -12256 3507 -12222 3541
rect -12160 4391 -12126 4425
rect -12160 4323 -12126 4357
rect -12160 4255 -12126 4289
rect -12160 4187 -12126 4221
rect -12160 4119 -12126 4153
rect -12160 4051 -12126 4085
rect -12160 3983 -12126 4017
rect -12160 3915 -12126 3949
rect -12160 3847 -12126 3881
rect -12160 3779 -12126 3813
rect -12160 3711 -12126 3745
rect -12160 3643 -12126 3677
rect -12160 3575 -12126 3609
rect -12160 3507 -12126 3541
rect -12064 4391 -12030 4425
rect -12064 4323 -12030 4357
rect -12064 4255 -12030 4289
rect -12064 4187 -12030 4221
rect -12064 4119 -12030 4153
rect -12064 4051 -12030 4085
rect -12064 3983 -12030 4017
rect -12064 3915 -12030 3949
rect -12064 3847 -12030 3881
rect -12064 3779 -12030 3813
rect -12064 3711 -12030 3745
rect -12064 3643 -12030 3677
rect -12064 3575 -12030 3609
rect -12064 3507 -12030 3541
rect -11968 4391 -11934 4425
rect -11968 4323 -11934 4357
rect -11968 4255 -11934 4289
rect -11968 4187 -11934 4221
rect -11968 4119 -11934 4153
rect -11968 4051 -11934 4085
rect -11968 3983 -11934 4017
rect -11968 3915 -11934 3949
rect -11968 3847 -11934 3881
rect -11968 3779 -11934 3813
rect -11968 3711 -11934 3745
rect -11968 3643 -11934 3677
rect -11968 3575 -11934 3609
rect -11968 3507 -11934 3541
rect -11760 4393 -11726 4427
rect -11760 4325 -11726 4359
rect -11760 4257 -11726 4291
rect -11760 4189 -11726 4223
rect -11760 4121 -11726 4155
rect -11760 4053 -11726 4087
rect -11760 3985 -11726 4019
rect -11760 3917 -11726 3951
rect -11760 3849 -11726 3883
rect -11760 3781 -11726 3815
rect -11760 3713 -11726 3747
rect -11760 3645 -11726 3679
rect -11760 3577 -11726 3611
rect -11760 3509 -11726 3543
rect -11664 4393 -11630 4427
rect -11664 4325 -11630 4359
rect -11664 4257 -11630 4291
rect -11664 4189 -11630 4223
rect -11664 4121 -11630 4155
rect -11664 4053 -11630 4087
rect -11664 3985 -11630 4019
rect -11664 3917 -11630 3951
rect -11664 3849 -11630 3883
rect -11664 3781 -11630 3815
rect -11664 3713 -11630 3747
rect -11664 3645 -11630 3679
rect -11664 3577 -11630 3611
rect -11664 3509 -11630 3543
rect -11568 4393 -11534 4427
rect -11568 4325 -11534 4359
rect -11568 4257 -11534 4291
rect -11568 4189 -11534 4223
rect -11568 4121 -11534 4155
rect -11568 4053 -11534 4087
rect -11568 3985 -11534 4019
rect -11568 3917 -11534 3951
rect -11568 3849 -11534 3883
rect -11568 3781 -11534 3815
rect -11568 3713 -11534 3747
rect -11568 3645 -11534 3679
rect -11568 3577 -11534 3611
rect -11568 3509 -11534 3543
rect -11472 4393 -11438 4427
rect -11472 4325 -11438 4359
rect -11472 4257 -11438 4291
rect -11472 4189 -11438 4223
rect -11472 4121 -11438 4155
rect -11472 4053 -11438 4087
rect -11472 3985 -11438 4019
rect -11472 3917 -11438 3951
rect -11472 3849 -11438 3883
rect -11472 3781 -11438 3815
rect -11472 3713 -11438 3747
rect -11472 3645 -11438 3679
rect -11472 3577 -11438 3611
rect -11472 3509 -11438 3543
rect -11376 4393 -11342 4427
rect -11376 4325 -11342 4359
rect -11376 4257 -11342 4291
rect -11376 4189 -11342 4223
rect -11376 4121 -11342 4155
rect -11376 4053 -11342 4087
rect -11376 3985 -11342 4019
rect -11376 3917 -11342 3951
rect -11376 3849 -11342 3883
rect -11376 3781 -11342 3815
rect -11376 3713 -11342 3747
rect -11376 3645 -11342 3679
rect -11376 3577 -11342 3611
rect -11376 3509 -11342 3543
rect -11280 4393 -11246 4427
rect -11280 4325 -11246 4359
rect -11280 4257 -11246 4291
rect -11280 4189 -11246 4223
rect -11280 4121 -11246 4155
rect -11280 4053 -11246 4087
rect -11280 3985 -11246 4019
rect -11280 3917 -11246 3951
rect -11280 3849 -11246 3883
rect -11280 3781 -11246 3815
rect -11280 3713 -11246 3747
rect -11280 3645 -11246 3679
rect -11280 3577 -11246 3611
rect -11280 3509 -11246 3543
rect -10290 4377 -10256 4411
rect -10290 4309 -10256 4343
rect -10290 4241 -10256 4275
rect -10290 4173 -10256 4207
rect -10290 4105 -10256 4139
rect -10290 4037 -10256 4071
rect -10290 3969 -10256 4003
rect -10290 3901 -10256 3935
rect -10290 3833 -10256 3867
rect -10290 3765 -10256 3799
rect -10290 3697 -10256 3731
rect -10290 3629 -10256 3663
rect -10290 3561 -10256 3595
rect -10290 3493 -10256 3527
rect -10194 4377 -10160 4411
rect -10194 4309 -10160 4343
rect -10194 4241 -10160 4275
rect -10194 4173 -10160 4207
rect -10194 4105 -10160 4139
rect -10194 4037 -10160 4071
rect -10194 3969 -10160 4003
rect -10194 3901 -10160 3935
rect -10194 3833 -10160 3867
rect -10194 3765 -10160 3799
rect -10194 3697 -10160 3731
rect -10194 3629 -10160 3663
rect -10194 3561 -10160 3595
rect -10194 3493 -10160 3527
rect -10098 4377 -10064 4411
rect -10098 4309 -10064 4343
rect -10098 4241 -10064 4275
rect -10098 4173 -10064 4207
rect -10098 4105 -10064 4139
rect -10098 4037 -10064 4071
rect -10098 3969 -10064 4003
rect -10098 3901 -10064 3935
rect -10098 3833 -10064 3867
rect -10098 3765 -10064 3799
rect -10098 3697 -10064 3731
rect -10098 3629 -10064 3663
rect -10098 3561 -10064 3595
rect -10098 3493 -10064 3527
rect -10002 4377 -9968 4411
rect -10002 4309 -9968 4343
rect -10002 4241 -9968 4275
rect -10002 4173 -9968 4207
rect -10002 4105 -9968 4139
rect -10002 4037 -9968 4071
rect -10002 3969 -9968 4003
rect -10002 3901 -9968 3935
rect -10002 3833 -9968 3867
rect -10002 3765 -9968 3799
rect -10002 3697 -9968 3731
rect -10002 3629 -9968 3663
rect -10002 3561 -9968 3595
rect -10002 3493 -9968 3527
rect -9906 4377 -9872 4411
rect -9906 4309 -9872 4343
rect -9906 4241 -9872 4275
rect -9906 4173 -9872 4207
rect -9906 4105 -9872 4139
rect -9906 4037 -9872 4071
rect -9906 3969 -9872 4003
rect -9906 3901 -9872 3935
rect -9906 3833 -9872 3867
rect -9906 3765 -9872 3799
rect -9906 3697 -9872 3731
rect -9906 3629 -9872 3663
rect -9906 3561 -9872 3595
rect -9906 3493 -9872 3527
rect -9810 4377 -9776 4411
rect -9810 4309 -9776 4343
rect -9810 4241 -9776 4275
rect -9810 4173 -9776 4207
rect -9810 4105 -9776 4139
rect -9810 4037 -9776 4071
rect -9810 3969 -9776 4003
rect -9810 3901 -9776 3935
rect -9810 3833 -9776 3867
rect -9810 3765 -9776 3799
rect -9810 3697 -9776 3731
rect -9810 3629 -9776 3663
rect -9810 3561 -9776 3595
rect -9810 3493 -9776 3527
rect -9714 4377 -9680 4411
rect -9714 4309 -9680 4343
rect -9714 4241 -9680 4275
rect -9714 4173 -9680 4207
rect -9714 4105 -9680 4139
rect -9714 4037 -9680 4071
rect -9714 3969 -9680 4003
rect -9714 3901 -9680 3935
rect -9714 3833 -9680 3867
rect -9714 3765 -9680 3799
rect -9714 3697 -9680 3731
rect -9714 3629 -9680 3663
rect -9714 3561 -9680 3595
rect -9714 3493 -9680 3527
rect -9618 4377 -9584 4411
rect -9618 4309 -9584 4343
rect -9618 4241 -9584 4275
rect -9618 4173 -9584 4207
rect -9618 4105 -9584 4139
rect -9618 4037 -9584 4071
rect -9618 3969 -9584 4003
rect -9618 3901 -9584 3935
rect -9618 3833 -9584 3867
rect -9618 3765 -9584 3799
rect -9618 3697 -9584 3731
rect -9618 3629 -9584 3663
rect -9618 3561 -9584 3595
rect -9618 3493 -9584 3527
rect -9522 4377 -9488 4411
rect -9522 4309 -9488 4343
rect -9522 4241 -9488 4275
rect -9522 4173 -9488 4207
rect -9522 4105 -9488 4139
rect -9522 4037 -9488 4071
rect -9522 3969 -9488 4003
rect -9522 3901 -9488 3935
rect -9522 3833 -9488 3867
rect -9522 3765 -9488 3799
rect -9522 3697 -9488 3731
rect -9522 3629 -9488 3663
rect -9522 3561 -9488 3595
rect -9522 3493 -9488 3527
rect -9426 4377 -9392 4411
rect -9426 4309 -9392 4343
rect -9426 4241 -9392 4275
rect -9426 4173 -9392 4207
rect -9426 4105 -9392 4139
rect -9426 4037 -9392 4071
rect -9426 3969 -9392 4003
rect -9426 3901 -9392 3935
rect -9426 3833 -9392 3867
rect -9426 3765 -9392 3799
rect -9426 3697 -9392 3731
rect -9426 3629 -9392 3663
rect -9426 3561 -9392 3595
rect -9426 3493 -9392 3527
rect -9330 4377 -9296 4411
rect -9330 4309 -9296 4343
rect -9330 4241 -9296 4275
rect -9330 4173 -9296 4207
rect -9330 4105 -9296 4139
rect -9330 4037 -9296 4071
rect -9330 3969 -9296 4003
rect -9330 3901 -9296 3935
rect -9330 3833 -9296 3867
rect -9330 3765 -9296 3799
rect -9330 3697 -9296 3731
rect -9330 3629 -9296 3663
rect -9330 3561 -9296 3595
rect -9330 3493 -9296 3527
rect -9234 4377 -9200 4411
rect -9234 4309 -9200 4343
rect -9234 4241 -9200 4275
rect -9234 4173 -9200 4207
rect -9234 4105 -9200 4139
rect -9234 4037 -9200 4071
rect -9234 3969 -9200 4003
rect -9234 3901 -9200 3935
rect -9234 3833 -9200 3867
rect -9234 3765 -9200 3799
rect -9234 3697 -9200 3731
rect -9234 3629 -9200 3663
rect -9234 3561 -9200 3595
rect -9234 3493 -9200 3527
rect -9138 4377 -9104 4411
rect -9138 4309 -9104 4343
rect -9138 4241 -9104 4275
rect -9138 4173 -9104 4207
rect -9138 4105 -9104 4139
rect -9138 4037 -9104 4071
rect -9138 3969 -9104 4003
rect -9138 3901 -9104 3935
rect -9138 3833 -9104 3867
rect -9138 3765 -9104 3799
rect -9138 3697 -9104 3731
rect -9138 3629 -9104 3663
rect -9138 3561 -9104 3595
rect -9138 3493 -9104 3527
rect -9042 4377 -9008 4411
rect -9042 4309 -9008 4343
rect -9042 4241 -9008 4275
rect -9042 4173 -9008 4207
rect -9042 4105 -9008 4139
rect -9042 4037 -9008 4071
rect -9042 3969 -9008 4003
rect -9042 3901 -9008 3935
rect -9042 3833 -9008 3867
rect -9042 3765 -9008 3799
rect -9042 3697 -9008 3731
rect -9042 3629 -9008 3663
rect -9042 3561 -9008 3595
rect -9042 3493 -9008 3527
rect -8946 4377 -8912 4411
rect -8946 4309 -8912 4343
rect -8946 4241 -8912 4275
rect -8946 4173 -8912 4207
rect -8946 4105 -8912 4139
rect -8946 4037 -8912 4071
rect -8946 3969 -8912 4003
rect -8946 3901 -8912 3935
rect -8946 3833 -8912 3867
rect -8946 3765 -8912 3799
rect -8946 3697 -8912 3731
rect -8946 3629 -8912 3663
rect -8946 3561 -8912 3595
rect -8946 3493 -8912 3527
rect -8850 4377 -8816 4411
rect -8850 4309 -8816 4343
rect -8850 4241 -8816 4275
rect -8850 4173 -8816 4207
rect -8850 4105 -8816 4139
rect -8850 4037 -8816 4071
rect -8850 3969 -8816 4003
rect -8850 3901 -8816 3935
rect -8850 3833 -8816 3867
rect -8850 3765 -8816 3799
rect -8850 3697 -8816 3731
rect -8850 3629 -8816 3663
rect -8850 3561 -8816 3595
rect -8850 3493 -8816 3527
rect -8754 4377 -8720 4411
rect -8754 4309 -8720 4343
rect -8754 4241 -8720 4275
rect -8754 4173 -8720 4207
rect -8754 4105 -8720 4139
rect -8754 4037 -8720 4071
rect -8754 3969 -8720 4003
rect -8754 3901 -8720 3935
rect -8754 3833 -8720 3867
rect -8754 3765 -8720 3799
rect -8754 3697 -8720 3731
rect -8754 3629 -8720 3663
rect -8754 3561 -8720 3595
rect -8754 3493 -8720 3527
rect -8658 4377 -8624 4411
rect -8658 4309 -8624 4343
rect -8658 4241 -8624 4275
rect -8658 4173 -8624 4207
rect -8658 4105 -8624 4139
rect -8658 4037 -8624 4071
rect -8658 3969 -8624 4003
rect -8658 3901 -8624 3935
rect -8658 3833 -8624 3867
rect -8658 3765 -8624 3799
rect -8658 3697 -8624 3731
rect -8658 3629 -8624 3663
rect -8658 3561 -8624 3595
rect -8658 3493 -8624 3527
rect -8562 4377 -8528 4411
rect -8562 4309 -8528 4343
rect -8562 4241 -8528 4275
rect -8562 4173 -8528 4207
rect -8562 4105 -8528 4139
rect -8562 4037 -8528 4071
rect -8562 3969 -8528 4003
rect -8562 3901 -8528 3935
rect -8562 3833 -8528 3867
rect -8562 3765 -8528 3799
rect -8562 3697 -8528 3731
rect -8562 3629 -8528 3663
rect -8562 3561 -8528 3595
rect -8562 3493 -8528 3527
rect -8466 4377 -8432 4411
rect -8466 4309 -8432 4343
rect -8466 4241 -8432 4275
rect -8466 4173 -8432 4207
rect -8466 4105 -8432 4139
rect -8466 4037 -8432 4071
rect -8466 3969 -8432 4003
rect -8466 3901 -8432 3935
rect -8466 3833 -8432 3867
rect -8466 3765 -8432 3799
rect -8466 3697 -8432 3731
rect -8466 3629 -8432 3663
rect -8466 3561 -8432 3595
rect -8466 3493 -8432 3527
rect -8370 4377 -8336 4411
rect -8370 4309 -8336 4343
rect -8370 4241 -8336 4275
rect -8370 4173 -8336 4207
rect -8370 4105 -8336 4139
rect -8370 4037 -8336 4071
rect -8370 3969 -8336 4003
rect -8370 3901 -8336 3935
rect -8370 3833 -8336 3867
rect -8370 3765 -8336 3799
rect -8370 3697 -8336 3731
rect -8370 3629 -8336 3663
rect -8370 3561 -8336 3595
rect -8370 3493 -8336 3527
rect -8146 4383 -8112 4417
rect -8146 4315 -8112 4349
rect -8146 4247 -8112 4281
rect -8146 4179 -8112 4213
rect -8146 4111 -8112 4145
rect -8146 4043 -8112 4077
rect -8146 3975 -8112 4009
rect -8146 3907 -8112 3941
rect -8146 3839 -8112 3873
rect -8146 3771 -8112 3805
rect -8146 3703 -8112 3737
rect -8146 3635 -8112 3669
rect -8146 3567 -8112 3601
rect -8146 3499 -8112 3533
rect -8050 4383 -8016 4417
rect -8050 4315 -8016 4349
rect -8050 4247 -8016 4281
rect -8050 4179 -8016 4213
rect -8050 4111 -8016 4145
rect -8050 4043 -8016 4077
rect -8050 3975 -8016 4009
rect -8050 3907 -8016 3941
rect -8050 3839 -8016 3873
rect -8050 3771 -8016 3805
rect -8050 3703 -8016 3737
rect -8050 3635 -8016 3669
rect -8050 3567 -8016 3601
rect -8050 3499 -8016 3533
rect -7954 4383 -7920 4417
rect -7954 4315 -7920 4349
rect -7954 4247 -7920 4281
rect -7954 4179 -7920 4213
rect -7954 4111 -7920 4145
rect -7954 4043 -7920 4077
rect -7954 3975 -7920 4009
rect -7954 3907 -7920 3941
rect -7954 3839 -7920 3873
rect -7954 3771 -7920 3805
rect -7954 3703 -7920 3737
rect -7954 3635 -7920 3669
rect -7954 3567 -7920 3601
rect -7954 3499 -7920 3533
rect -7858 4383 -7824 4417
rect -7858 4315 -7824 4349
rect -7858 4247 -7824 4281
rect -7858 4179 -7824 4213
rect -7858 4111 -7824 4145
rect -7858 4043 -7824 4077
rect -7858 3975 -7824 4009
rect -7858 3907 -7824 3941
rect -7858 3839 -7824 3873
rect -7858 3771 -7824 3805
rect -7858 3703 -7824 3737
rect -7858 3635 -7824 3669
rect -7858 3567 -7824 3601
rect -7858 3499 -7824 3533
rect -7762 4383 -7728 4417
rect -7762 4315 -7728 4349
rect -7762 4247 -7728 4281
rect -7762 4179 -7728 4213
rect -7762 4111 -7728 4145
rect -7762 4043 -7728 4077
rect -7762 3975 -7728 4009
rect -7762 3907 -7728 3941
rect -7762 3839 -7728 3873
rect -7762 3771 -7728 3805
rect -7762 3703 -7728 3737
rect -7762 3635 -7728 3669
rect -7762 3567 -7728 3601
rect -7762 3499 -7728 3533
rect -7666 4383 -7632 4417
rect -7666 4315 -7632 4349
rect -7666 4247 -7632 4281
rect -7666 4179 -7632 4213
rect -7666 4111 -7632 4145
rect -7666 4043 -7632 4077
rect -7666 3975 -7632 4009
rect -7666 3907 -7632 3941
rect -7666 3839 -7632 3873
rect -7666 3771 -7632 3805
rect -7666 3703 -7632 3737
rect -7666 3635 -7632 3669
rect -7666 3567 -7632 3601
rect -7666 3499 -7632 3533
rect -7570 4383 -7536 4417
rect -7570 4315 -7536 4349
rect -7570 4247 -7536 4281
rect -7570 4179 -7536 4213
rect -7570 4111 -7536 4145
rect -7570 4043 -7536 4077
rect -7570 3975 -7536 4009
rect -7570 3907 -7536 3941
rect -7570 3839 -7536 3873
rect -7570 3771 -7536 3805
rect -7570 3703 -7536 3737
rect -7570 3635 -7536 3669
rect -7570 3567 -7536 3601
rect -7570 3499 -7536 3533
rect -7474 4383 -7440 4417
rect -7474 4315 -7440 4349
rect -7474 4247 -7440 4281
rect -7474 4179 -7440 4213
rect -7474 4111 -7440 4145
rect -7474 4043 -7440 4077
rect -7474 3975 -7440 4009
rect -7474 3907 -7440 3941
rect -7474 3839 -7440 3873
rect -7474 3771 -7440 3805
rect -7474 3703 -7440 3737
rect -7474 3635 -7440 3669
rect -7474 3567 -7440 3601
rect -7474 3499 -7440 3533
rect -7378 4383 -7344 4417
rect -7378 4315 -7344 4349
rect -7378 4247 -7344 4281
rect -7378 4179 -7344 4213
rect -7378 4111 -7344 4145
rect -7378 4043 -7344 4077
rect -7378 3975 -7344 4009
rect -7378 3907 -7344 3941
rect -7378 3839 -7344 3873
rect -7378 3771 -7344 3805
rect -7378 3703 -7344 3737
rect -7378 3635 -7344 3669
rect -7378 3567 -7344 3601
rect -7378 3499 -7344 3533
rect -7282 4383 -7248 4417
rect -7282 4315 -7248 4349
rect -7282 4247 -7248 4281
rect -7282 4179 -7248 4213
rect -7282 4111 -7248 4145
rect -7282 4043 -7248 4077
rect -7282 3975 -7248 4009
rect -7282 3907 -7248 3941
rect -7282 3839 -7248 3873
rect -7282 3771 -7248 3805
rect -7282 3703 -7248 3737
rect -7282 3635 -7248 3669
rect -7282 3567 -7248 3601
rect -7282 3499 -7248 3533
rect -7186 4383 -7152 4417
rect -7186 4315 -7152 4349
rect -7186 4247 -7152 4281
rect -7186 4179 -7152 4213
rect -7186 4111 -7152 4145
rect -7186 4043 -7152 4077
rect -7186 3975 -7152 4009
rect -7186 3907 -7152 3941
rect -7186 3839 -7152 3873
rect -7186 3771 -7152 3805
rect -7186 3703 -7152 3737
rect -7186 3635 -7152 3669
rect -7186 3567 -7152 3601
rect -7186 3499 -7152 3533
rect -7090 4383 -7056 4417
rect -7090 4315 -7056 4349
rect -7090 4247 -7056 4281
rect -7090 4179 -7056 4213
rect -7090 4111 -7056 4145
rect -7090 4043 -7056 4077
rect -7090 3975 -7056 4009
rect -7090 3907 -7056 3941
rect -7090 3839 -7056 3873
rect -7090 3771 -7056 3805
rect -7090 3703 -7056 3737
rect -7090 3635 -7056 3669
rect -7090 3567 -7056 3601
rect -7090 3499 -7056 3533
rect -6994 4383 -6960 4417
rect -6994 4315 -6960 4349
rect -6994 4247 -6960 4281
rect -6994 4179 -6960 4213
rect -6994 4111 -6960 4145
rect -6994 4043 -6960 4077
rect -6994 3975 -6960 4009
rect -6994 3907 -6960 3941
rect -6994 3839 -6960 3873
rect -6994 3771 -6960 3805
rect -6994 3703 -6960 3737
rect -6994 3635 -6960 3669
rect -6994 3567 -6960 3601
rect -6994 3499 -6960 3533
rect -6898 4383 -6864 4417
rect -6898 4315 -6864 4349
rect -6898 4247 -6864 4281
rect -6898 4179 -6864 4213
rect -6898 4111 -6864 4145
rect -6898 4043 -6864 4077
rect -6898 3975 -6864 4009
rect -6898 3907 -6864 3941
rect -6898 3839 -6864 3873
rect -6898 3771 -6864 3805
rect -6898 3703 -6864 3737
rect -6898 3635 -6864 3669
rect -6898 3567 -6864 3601
rect -6898 3499 -6864 3533
rect -6802 4383 -6768 4417
rect -6802 4315 -6768 4349
rect -6802 4247 -6768 4281
rect -6802 4179 -6768 4213
rect -6802 4111 -6768 4145
rect -6802 4043 -6768 4077
rect -6802 3975 -6768 4009
rect -6802 3907 -6768 3941
rect -6802 3839 -6768 3873
rect -6802 3771 -6768 3805
rect -6802 3703 -6768 3737
rect -6802 3635 -6768 3669
rect -6802 3567 -6768 3601
rect -6802 3499 -6768 3533
rect -6706 4383 -6672 4417
rect -6706 4315 -6672 4349
rect -6706 4247 -6672 4281
rect -6706 4179 -6672 4213
rect -6706 4111 -6672 4145
rect -6706 4043 -6672 4077
rect -6706 3975 -6672 4009
rect -6706 3907 -6672 3941
rect -6706 3839 -6672 3873
rect -6706 3771 -6672 3805
rect -6706 3703 -6672 3737
rect -6706 3635 -6672 3669
rect -6706 3567 -6672 3601
rect -6706 3499 -6672 3533
rect -6462 4389 -6428 4423
rect -6462 4321 -6428 4355
rect -6462 4253 -6428 4287
rect -6462 4185 -6428 4219
rect -6462 4117 -6428 4151
rect -6462 4049 -6428 4083
rect -6462 3981 -6428 4015
rect -6462 3913 -6428 3947
rect -6462 3845 -6428 3879
rect -6462 3777 -6428 3811
rect -6462 3709 -6428 3743
rect -6462 3641 -6428 3675
rect -6462 3573 -6428 3607
rect -6462 3505 -6428 3539
rect -6366 4389 -6332 4423
rect -6366 4321 -6332 4355
rect -6366 4253 -6332 4287
rect -6366 4185 -6332 4219
rect -6366 4117 -6332 4151
rect -6366 4049 -6332 4083
rect -6366 3981 -6332 4015
rect -6366 3913 -6332 3947
rect -6366 3845 -6332 3879
rect -6366 3777 -6332 3811
rect -6366 3709 -6332 3743
rect -6366 3641 -6332 3675
rect -6366 3573 -6332 3607
rect -6366 3505 -6332 3539
rect -6270 4389 -6236 4423
rect -6270 4321 -6236 4355
rect -6270 4253 -6236 4287
rect -6270 4185 -6236 4219
rect -6270 4117 -6236 4151
rect -6270 4049 -6236 4083
rect -6270 3981 -6236 4015
rect -6270 3913 -6236 3947
rect -6270 3845 -6236 3879
rect -6270 3777 -6236 3811
rect -6270 3709 -6236 3743
rect -6270 3641 -6236 3675
rect -6270 3573 -6236 3607
rect -6270 3505 -6236 3539
rect -6174 4389 -6140 4423
rect -6174 4321 -6140 4355
rect -6174 4253 -6140 4287
rect -6174 4185 -6140 4219
rect -6174 4117 -6140 4151
rect -6174 4049 -6140 4083
rect -6174 3981 -6140 4015
rect -6174 3913 -6140 3947
rect -6174 3845 -6140 3879
rect -6174 3777 -6140 3811
rect -6174 3709 -6140 3743
rect -6174 3641 -6140 3675
rect -6174 3573 -6140 3607
rect -6174 3505 -6140 3539
rect -6078 4389 -6044 4423
rect -6078 4321 -6044 4355
rect -6078 4253 -6044 4287
rect -6078 4185 -6044 4219
rect -6078 4117 -6044 4151
rect -6078 4049 -6044 4083
rect -6078 3981 -6044 4015
rect -6078 3913 -6044 3947
rect -6078 3845 -6044 3879
rect -6078 3777 -6044 3811
rect -6078 3709 -6044 3743
rect -6078 3641 -6044 3675
rect -6078 3573 -6044 3607
rect -6078 3505 -6044 3539
rect -5982 4389 -5948 4423
rect -5982 4321 -5948 4355
rect -5982 4253 -5948 4287
rect -5982 4185 -5948 4219
rect -5982 4117 -5948 4151
rect -5982 4049 -5948 4083
rect -5982 3981 -5948 4015
rect -5982 3913 -5948 3947
rect -5982 3845 -5948 3879
rect -5982 3777 -5948 3811
rect -5982 3709 -5948 3743
rect -5982 3641 -5948 3675
rect -5982 3573 -5948 3607
rect -5982 3505 -5948 3539
rect -5886 4389 -5852 4423
rect -5886 4321 -5852 4355
rect -5886 4253 -5852 4287
rect -5886 4185 -5852 4219
rect -5886 4117 -5852 4151
rect -5886 4049 -5852 4083
rect -5886 3981 -5852 4015
rect -5886 3913 -5852 3947
rect -5886 3845 -5852 3879
rect -5886 3777 -5852 3811
rect -5886 3709 -5852 3743
rect -5886 3641 -5852 3675
rect -5886 3573 -5852 3607
rect -5886 3505 -5852 3539
rect -5790 4389 -5756 4423
rect -5790 4321 -5756 4355
rect -5790 4253 -5756 4287
rect -5790 4185 -5756 4219
rect -5790 4117 -5756 4151
rect -5790 4049 -5756 4083
rect -5790 3981 -5756 4015
rect -5790 3913 -5756 3947
rect -5790 3845 -5756 3879
rect -5790 3777 -5756 3811
rect -5790 3709 -5756 3743
rect -5790 3641 -5756 3675
rect -5790 3573 -5756 3607
rect -5790 3505 -5756 3539
rect -5694 4389 -5660 4423
rect -5694 4321 -5660 4355
rect -5694 4253 -5660 4287
rect -5694 4185 -5660 4219
rect -5694 4117 -5660 4151
rect -5694 4049 -5660 4083
rect -5694 3981 -5660 4015
rect -5694 3913 -5660 3947
rect -5694 3845 -5660 3879
rect -5694 3777 -5660 3811
rect -5694 3709 -5660 3743
rect -5694 3641 -5660 3675
rect -5694 3573 -5660 3607
rect -5694 3505 -5660 3539
rect -5598 4389 -5564 4423
rect -5598 4321 -5564 4355
rect -5598 4253 -5564 4287
rect -5598 4185 -5564 4219
rect -5598 4117 -5564 4151
rect -5598 4049 -5564 4083
rect -5598 3981 -5564 4015
rect -5598 3913 -5564 3947
rect -5598 3845 -5564 3879
rect -5598 3777 -5564 3811
rect -5598 3709 -5564 3743
rect -5598 3641 -5564 3675
rect -5598 3573 -5564 3607
rect -5598 3505 -5564 3539
rect -5502 4389 -5468 4423
rect -5502 4321 -5468 4355
rect -5502 4253 -5468 4287
rect -5502 4185 -5468 4219
rect -5502 4117 -5468 4151
rect -5502 4049 -5468 4083
rect -5502 3981 -5468 4015
rect -5502 3913 -5468 3947
rect -5502 3845 -5468 3879
rect -5502 3777 -5468 3811
rect -5502 3709 -5468 3743
rect -5502 3641 -5468 3675
rect -5502 3573 -5468 3607
rect -5502 3505 -5468 3539
rect -5294 4391 -5260 4425
rect -5294 4323 -5260 4357
rect -5294 4255 -5260 4289
rect -5294 4187 -5260 4221
rect -5294 4119 -5260 4153
rect -5294 4051 -5260 4085
rect -5294 3983 -5260 4017
rect -5294 3915 -5260 3949
rect -5294 3847 -5260 3881
rect -5294 3779 -5260 3813
rect -5294 3711 -5260 3745
rect -5294 3643 -5260 3677
rect -5294 3575 -5260 3609
rect -5294 3507 -5260 3541
rect -5198 4391 -5164 4425
rect -5198 4323 -5164 4357
rect -5198 4255 -5164 4289
rect -5198 4187 -5164 4221
rect -5198 4119 -5164 4153
rect -5198 4051 -5164 4085
rect -5198 3983 -5164 4017
rect -5198 3915 -5164 3949
rect -5198 3847 -5164 3881
rect -5198 3779 -5164 3813
rect -5198 3711 -5164 3745
rect -5198 3643 -5164 3677
rect -5198 3575 -5164 3609
rect -5198 3507 -5164 3541
rect -5102 4391 -5068 4425
rect -5102 4323 -5068 4357
rect -5102 4255 -5068 4289
rect -5102 4187 -5068 4221
rect -5102 4119 -5068 4153
rect -5102 4051 -5068 4085
rect -5102 3983 -5068 4017
rect -5102 3915 -5068 3949
rect -5102 3847 -5068 3881
rect -5102 3779 -5068 3813
rect -5102 3711 -5068 3745
rect -5102 3643 -5068 3677
rect -5102 3575 -5068 3609
rect -5102 3507 -5068 3541
rect -5006 4391 -4972 4425
rect -5006 4323 -4972 4357
rect -5006 4255 -4972 4289
rect -5006 4187 -4972 4221
rect -5006 4119 -4972 4153
rect -5006 4051 -4972 4085
rect -5006 3983 -4972 4017
rect -5006 3915 -4972 3949
rect -5006 3847 -4972 3881
rect -5006 3779 -4972 3813
rect -5006 3711 -4972 3745
rect -5006 3643 -4972 3677
rect -5006 3575 -4972 3609
rect -5006 3507 -4972 3541
rect -4910 4391 -4876 4425
rect -4910 4323 -4876 4357
rect -4910 4255 -4876 4289
rect -4910 4187 -4876 4221
rect -4910 4119 -4876 4153
rect -4910 4051 -4876 4085
rect -4910 3983 -4876 4017
rect -4910 3915 -4876 3949
rect -4910 3847 -4876 3881
rect -4910 3779 -4876 3813
rect -4910 3711 -4876 3745
rect -4910 3643 -4876 3677
rect -4910 3575 -4876 3609
rect -4910 3507 -4876 3541
rect -4814 4391 -4780 4425
rect -4814 4323 -4780 4357
rect -4814 4255 -4780 4289
rect -4814 4187 -4780 4221
rect -4814 4119 -4780 4153
rect -4814 4051 -4780 4085
rect -4814 3983 -4780 4017
rect -4814 3915 -4780 3949
rect 1484 4461 1518 4495
rect 1484 4393 1518 4427
rect 1484 4325 1518 4359
rect 1484 4257 1518 4291
rect 1484 4189 1518 4223
rect 1484 4121 1518 4155
rect 1484 4053 1518 4087
rect 1484 3985 1518 4019
rect 1580 4869 1614 4903
rect 1580 4801 1614 4835
rect 1580 4733 1614 4767
rect 1580 4665 1614 4699
rect 1580 4597 1614 4631
rect 1580 4529 1614 4563
rect 1580 4461 1614 4495
rect 1580 4393 1614 4427
rect 1580 4325 1614 4359
rect 1580 4257 1614 4291
rect 1580 4189 1614 4223
rect 1580 4121 1614 4155
rect 1580 4053 1614 4087
rect 1580 3985 1614 4019
rect 1676 4869 1710 4903
rect 1676 4801 1710 4835
rect 1676 4733 1710 4767
rect 1676 4665 1710 4699
rect 1676 4597 1710 4631
rect 1676 4529 1710 4563
rect 1676 4461 1710 4495
rect 1676 4393 1710 4427
rect 1676 4325 1710 4359
rect 1676 4257 1710 4291
rect 1676 4189 1710 4223
rect 1676 4121 1710 4155
rect 1676 4053 1710 4087
rect 1676 3985 1710 4019
rect 1772 4869 1806 4903
rect 1772 4801 1806 4835
rect 1772 4733 1806 4767
rect 1772 4665 1806 4699
rect 1772 4597 1806 4631
rect 1772 4529 1806 4563
rect 1772 4461 1806 4495
rect 1772 4393 1806 4427
rect 1772 4325 1806 4359
rect 1772 4257 1806 4291
rect 1772 4189 1806 4223
rect 1772 4121 1806 4155
rect 1772 4053 1806 4087
rect 1772 3985 1806 4019
rect 15518 4977 15552 5011
rect 1868 4869 1902 4903
rect 1868 4801 1902 4835
rect 1868 4733 1902 4767
rect 1868 4665 1902 4699
rect 1868 4597 1902 4631
rect 1868 4529 1902 4563
rect 1868 4461 1902 4495
rect 1868 4393 1902 4427
rect 1868 4325 1902 4359
rect 1868 4257 1902 4291
rect 1868 4189 1902 4223
rect 1868 4121 1902 4155
rect 1868 4053 1902 4087
rect 1868 3985 1902 4019
rect 4440 4853 4474 4887
rect 4440 4785 4474 4819
rect 4440 4717 4474 4751
rect 4440 4649 4474 4683
rect 4440 4581 4474 4615
rect 4440 4513 4474 4547
rect 4440 4445 4474 4479
rect 4440 4377 4474 4411
rect 4440 4309 4474 4343
rect 4440 4241 4474 4275
rect 4440 4173 4474 4207
rect 4440 4105 4474 4139
rect 4440 4037 4474 4071
rect 4440 3969 4474 4003
rect -4814 3847 -4780 3881
rect 4536 4853 4570 4887
rect 4536 4785 4570 4819
rect 4536 4717 4570 4751
rect 4536 4649 4570 4683
rect 4536 4581 4570 4615
rect 4536 4513 4570 4547
rect 4536 4445 4570 4479
rect 4536 4377 4570 4411
rect 4536 4309 4570 4343
rect 4536 4241 4570 4275
rect 4536 4173 4570 4207
rect 4536 4105 4570 4139
rect 4536 4037 4570 4071
rect 4536 3969 4570 4003
rect 4632 4853 4666 4887
rect 4632 4785 4666 4819
rect 4632 4717 4666 4751
rect 4632 4649 4666 4683
rect 4632 4581 4666 4615
rect 4632 4513 4666 4547
rect 4632 4445 4666 4479
rect 4632 4377 4666 4411
rect 4632 4309 4666 4343
rect 4632 4241 4666 4275
rect 4632 4173 4666 4207
rect 4632 4105 4666 4139
rect 4632 4037 4666 4071
rect 4632 3969 4666 4003
rect 4728 4853 4762 4887
rect 4728 4785 4762 4819
rect 4728 4717 4762 4751
rect 4728 4649 4762 4683
rect 4728 4581 4762 4615
rect 4728 4513 4762 4547
rect 4728 4445 4762 4479
rect 4728 4377 4762 4411
rect 4728 4309 4762 4343
rect 4728 4241 4762 4275
rect 4728 4173 4762 4207
rect 4728 4105 4762 4139
rect 4728 4037 4762 4071
rect 4728 3969 4762 4003
rect 4824 4853 4858 4887
rect 4824 4785 4858 4819
rect 4824 4717 4858 4751
rect 4824 4649 4858 4683
rect 4824 4581 4858 4615
rect 4824 4513 4858 4547
rect 4824 4445 4858 4479
rect 4824 4377 4858 4411
rect 4824 4309 4858 4343
rect 4824 4241 4858 4275
rect 4824 4173 4858 4207
rect 4824 4105 4858 4139
rect 4824 4037 4858 4071
rect 4824 3969 4858 4003
rect 7470 4853 7504 4887
rect 7470 4785 7504 4819
rect 7470 4717 7504 4751
rect 7470 4649 7504 4683
rect 7470 4581 7504 4615
rect 7470 4513 7504 4547
rect 7470 4445 7504 4479
rect 7470 4377 7504 4411
rect 7470 4309 7504 4343
rect 7470 4241 7504 4275
rect 7470 4173 7504 4207
rect 7470 4105 7504 4139
rect 7470 4037 7504 4071
rect 7470 3969 7504 4003
rect 7566 4853 7600 4887
rect 7566 4785 7600 4819
rect 7566 4717 7600 4751
rect 7566 4649 7600 4683
rect 7566 4581 7600 4615
rect 7566 4513 7600 4547
rect 7566 4445 7600 4479
rect 7566 4377 7600 4411
rect 7566 4309 7600 4343
rect 7566 4241 7600 4275
rect 7566 4173 7600 4207
rect 7566 4105 7600 4139
rect 7566 4037 7600 4071
rect 7566 3969 7600 4003
rect 7662 4853 7696 4887
rect 7662 4785 7696 4819
rect 7662 4717 7696 4751
rect 7662 4649 7696 4683
rect 7662 4581 7696 4615
rect 7662 4513 7696 4547
rect 7662 4445 7696 4479
rect 7662 4377 7696 4411
rect 7662 4309 7696 4343
rect 7662 4241 7696 4275
rect 7662 4173 7696 4207
rect 7662 4105 7696 4139
rect 7662 4037 7696 4071
rect 7662 3969 7696 4003
rect 7758 4853 7792 4887
rect 7758 4785 7792 4819
rect 7758 4717 7792 4751
rect 7758 4649 7792 4683
rect 7758 4581 7792 4615
rect 7758 4513 7792 4547
rect 7758 4445 7792 4479
rect 7758 4377 7792 4411
rect 7758 4309 7792 4343
rect 7758 4241 7792 4275
rect 7758 4173 7792 4207
rect 7758 4105 7792 4139
rect 7758 4037 7792 4071
rect 7758 3969 7792 4003
rect 7854 4853 7888 4887
rect 7854 4785 7888 4819
rect 7854 4717 7888 4751
rect 7854 4649 7888 4683
rect 7854 4581 7888 4615
rect 7854 4513 7888 4547
rect 7854 4445 7888 4479
rect 7854 4377 7888 4411
rect 7854 4309 7888 4343
rect 7854 4241 7888 4275
rect 7854 4173 7888 4207
rect 7854 4105 7888 4139
rect 7854 4037 7888 4071
rect 7854 3969 7888 4003
rect 10558 4851 10592 4885
rect 10558 4783 10592 4817
rect 10558 4715 10592 4749
rect 10558 4647 10592 4681
rect 10558 4579 10592 4613
rect 10558 4511 10592 4545
rect 10558 4443 10592 4477
rect 10558 4375 10592 4409
rect 10558 4307 10592 4341
rect 10558 4239 10592 4273
rect 10558 4171 10592 4205
rect 10558 4103 10592 4137
rect 10558 4035 10592 4069
rect 10558 3967 10592 4001
rect -4814 3779 -4780 3813
rect 10654 4851 10688 4885
rect 10654 4783 10688 4817
rect 10654 4715 10688 4749
rect 10654 4647 10688 4681
rect 10654 4579 10688 4613
rect 10654 4511 10688 4545
rect 10654 4443 10688 4477
rect 10654 4375 10688 4409
rect 10654 4307 10688 4341
rect 10654 4239 10688 4273
rect 10654 4171 10688 4205
rect 10654 4103 10688 4137
rect 10654 4035 10688 4069
rect 10654 3967 10688 4001
rect 10750 4851 10784 4885
rect 10750 4783 10784 4817
rect 10750 4715 10784 4749
rect 10750 4647 10784 4681
rect 10750 4579 10784 4613
rect 10750 4511 10784 4545
rect 10750 4443 10784 4477
rect 10750 4375 10784 4409
rect 10750 4307 10784 4341
rect 10750 4239 10784 4273
rect 10750 4171 10784 4205
rect 10750 4103 10784 4137
rect 10750 4035 10784 4069
rect 10750 3967 10784 4001
rect 10846 4851 10880 4885
rect 10846 4783 10880 4817
rect 10846 4715 10880 4749
rect 10846 4647 10880 4681
rect 10846 4579 10880 4613
rect 10846 4511 10880 4545
rect 10846 4443 10880 4477
rect 10846 4375 10880 4409
rect 10846 4307 10880 4341
rect 10846 4239 10880 4273
rect 10846 4171 10880 4205
rect 10846 4103 10880 4137
rect 10846 4035 10880 4069
rect 10846 3967 10880 4001
rect 15518 4909 15552 4943
rect 10942 4851 10976 4885
rect 10942 4783 10976 4817
rect 10942 4715 10976 4749
rect 10942 4647 10976 4681
rect 10942 4579 10976 4613
rect 10942 4511 10976 4545
rect 10942 4443 10976 4477
rect 10942 4375 10976 4409
rect 10942 4307 10976 4341
rect 10942 4239 10976 4273
rect 10942 4171 10976 4205
rect 10942 4103 10976 4137
rect 10942 4035 10976 4069
rect 10942 3967 10976 4001
rect 13714 4825 13748 4859
rect 13714 4757 13748 4791
rect 13714 4689 13748 4723
rect 13714 4621 13748 4655
rect 13714 4553 13748 4587
rect 13714 4485 13748 4519
rect 13714 4417 13748 4451
rect 13714 4349 13748 4383
rect 13714 4281 13748 4315
rect 13714 4213 13748 4247
rect 13714 4145 13748 4179
rect 13714 4077 13748 4111
rect 13714 4009 13748 4043
rect 13714 3941 13748 3975
rect -4814 3711 -4780 3745
rect 13810 4825 13844 4859
rect 13810 4757 13844 4791
rect 13810 4689 13844 4723
rect 13810 4621 13844 4655
rect 13810 4553 13844 4587
rect 13810 4485 13844 4519
rect 13810 4417 13844 4451
rect 13810 4349 13844 4383
rect 13810 4281 13844 4315
rect 13810 4213 13844 4247
rect 13810 4145 13844 4179
rect 13810 4077 13844 4111
rect 13810 4009 13844 4043
rect 13810 3941 13844 3975
rect 13906 4825 13940 4859
rect 13906 4757 13940 4791
rect 13906 4689 13940 4723
rect 13906 4621 13940 4655
rect 13906 4553 13940 4587
rect 13906 4485 13940 4519
rect 13906 4417 13940 4451
rect 13906 4349 13940 4383
rect 13906 4281 13940 4315
rect 13906 4213 13940 4247
rect 13906 4145 13940 4179
rect 13906 4077 13940 4111
rect 13906 4009 13940 4043
rect 13906 3941 13940 3975
rect 14002 4825 14036 4859
rect 14002 4757 14036 4791
rect 14002 4689 14036 4723
rect 14002 4621 14036 4655
rect 14002 4553 14036 4587
rect 14002 4485 14036 4519
rect 14002 4417 14036 4451
rect 14002 4349 14036 4383
rect 14002 4281 14036 4315
rect 14002 4213 14036 4247
rect 14002 4145 14036 4179
rect 14002 4077 14036 4111
rect 14002 4009 14036 4043
rect 14002 3941 14036 3975
rect 14098 4825 14132 4859
rect 14098 4757 14132 4791
rect 14098 4689 14132 4723
rect 14098 4621 14132 4655
rect 14098 4553 14132 4587
rect 14098 4485 14132 4519
rect 14098 4417 14132 4451
rect 14098 4349 14132 4383
rect 14098 4281 14132 4315
rect 14098 4213 14132 4247
rect 14098 4145 14132 4179
rect 14098 4077 14132 4111
rect 14098 4009 14132 4043
rect 14098 3941 14132 3975
rect 15518 4841 15552 4875
rect 15518 4773 15552 4807
rect 15518 4705 15552 4739
rect 15518 4637 15552 4671
rect 15518 4569 15552 4603
rect 15518 4501 15552 4535
rect 15518 4433 15552 4467
rect 15518 4365 15552 4399
rect 15518 4297 15552 4331
rect 15518 4229 15552 4263
rect 15518 4161 15552 4195
rect 15518 4093 15552 4127
rect 15518 4025 15552 4059
rect 15518 3957 15552 3991
rect 15614 5861 15648 5895
rect 15614 5793 15648 5827
rect 15614 5725 15648 5759
rect 15614 5657 15648 5691
rect 15614 5589 15648 5623
rect 15614 5521 15648 5555
rect 15614 5453 15648 5487
rect 15614 5385 15648 5419
rect 15614 5317 15648 5351
rect 15614 5249 15648 5283
rect 15614 5181 15648 5215
rect 15614 5113 15648 5147
rect 15614 5045 15648 5079
rect 15614 4977 15648 5011
rect 15614 4909 15648 4943
rect 15614 4841 15648 4875
rect 15614 4773 15648 4807
rect 15614 4705 15648 4739
rect 15614 4637 15648 4671
rect 15614 4569 15648 4603
rect 15614 4501 15648 4535
rect 15614 4433 15648 4467
rect 15614 4365 15648 4399
rect 15614 4297 15648 4331
rect 15614 4229 15648 4263
rect 15614 4161 15648 4195
rect 15614 4093 15648 4127
rect 15614 4025 15648 4059
rect 15614 3957 15648 3991
rect 15710 5861 15744 5895
rect 15710 5793 15744 5827
rect 15710 5725 15744 5759
rect 15710 5657 15744 5691
rect 15710 5589 15744 5623
rect 15710 5521 15744 5555
rect 15710 5453 15744 5487
rect 15710 5385 15744 5419
rect 15710 5317 15744 5351
rect 15710 5249 15744 5283
rect 15710 5181 15744 5215
rect 15710 5113 15744 5147
rect 15710 5045 15744 5079
rect 15710 4977 15744 5011
rect 15710 4909 15744 4943
rect 15710 4841 15744 4875
rect 15710 4773 15744 4807
rect 15710 4705 15744 4739
rect 15710 4637 15744 4671
rect 15710 4569 15744 4603
rect 15710 4501 15744 4535
rect 15710 4433 15744 4467
rect 15710 4365 15744 4399
rect 15710 4297 15744 4331
rect 15710 4229 15744 4263
rect 15710 4161 15744 4195
rect 16782 5055 16816 5089
rect 16782 4987 16816 5021
rect 16782 4919 16816 4953
rect 16782 4851 16816 4885
rect 16782 4783 16816 4817
rect 16782 4715 16816 4749
rect 16782 4647 16816 4681
rect 16782 4579 16816 4613
rect 16782 4511 16816 4545
rect 16782 4443 16816 4477
rect 16782 4375 16816 4409
rect 16782 4307 16816 4341
rect 16782 4239 16816 4273
rect 16782 4171 16816 4205
rect 16878 5055 16912 5089
rect 16878 4987 16912 5021
rect 16878 4919 16912 4953
rect 16878 4851 16912 4885
rect 16878 4783 16912 4817
rect 16878 4715 16912 4749
rect 16878 4647 16912 4681
rect 16878 4579 16912 4613
rect 16878 4511 16912 4545
rect 16878 4443 16912 4477
rect 16878 4375 16912 4409
rect 16878 4307 16912 4341
rect 16878 4239 16912 4273
rect 16878 4171 16912 4205
rect 16974 5055 17008 5089
rect 16974 4987 17008 5021
rect 16974 4919 17008 4953
rect 16974 4851 17008 4885
rect 16974 4783 17008 4817
rect 16974 4715 17008 4749
rect 16974 4647 17008 4681
rect 16974 4579 17008 4613
rect 16974 4511 17008 4545
rect 16974 4443 17008 4477
rect 16974 4375 17008 4409
rect 16974 4307 17008 4341
rect 16974 4239 17008 4273
rect 16974 4171 17008 4205
rect 17070 5055 17104 5089
rect 17070 4987 17104 5021
rect 17070 4919 17104 4953
rect 17070 4851 17104 4885
rect 17070 4783 17104 4817
rect 17070 4715 17104 4749
rect 17070 4647 17104 4681
rect 17070 4579 17104 4613
rect 17070 4511 17104 4545
rect 17070 4443 17104 4477
rect 17070 4375 17104 4409
rect 17070 4307 17104 4341
rect 17070 4239 17104 4273
rect 17070 4171 17104 4205
rect 17166 5055 17200 5089
rect 17166 4987 17200 5021
rect 17166 4919 17200 4953
rect 17166 4851 17200 4885
rect 17166 4783 17200 4817
rect 17166 4715 17200 4749
rect 17166 4647 17200 4681
rect 17166 4579 17200 4613
rect 17166 4511 17200 4545
rect 17166 4443 17200 4477
rect 17166 4375 17200 4409
rect 17166 4307 17200 4341
rect 17166 4239 17200 4273
rect 17166 4171 17200 4205
rect 17262 5055 17296 5089
rect 17262 4987 17296 5021
rect 17262 4919 17296 4953
rect 17262 4851 17296 4885
rect 17262 4783 17296 4817
rect 17262 4715 17296 4749
rect 17262 4647 17296 4681
rect 17262 4579 17296 4613
rect 17262 4511 17296 4545
rect 17262 4443 17296 4477
rect 17262 4375 17296 4409
rect 17262 4307 17296 4341
rect 17262 4239 17296 4273
rect 17262 4171 17296 4205
rect 17470 5053 17504 5087
rect 17470 4985 17504 5019
rect 17470 4917 17504 4951
rect 17470 4849 17504 4883
rect 17470 4781 17504 4815
rect 17470 4713 17504 4747
rect 17470 4645 17504 4679
rect 17470 4577 17504 4611
rect 17470 4509 17504 4543
rect 17470 4441 17504 4475
rect 17470 4373 17504 4407
rect 17470 4305 17504 4339
rect 17470 4237 17504 4271
rect 17470 4169 17504 4203
rect 15710 4093 15744 4127
rect 15710 4025 15744 4059
rect 15710 3957 15744 3991
rect 17566 5053 17600 5087
rect 17566 4985 17600 5019
rect 17566 4917 17600 4951
rect 17566 4849 17600 4883
rect 17566 4781 17600 4815
rect 17566 4713 17600 4747
rect 17566 4645 17600 4679
rect 17566 4577 17600 4611
rect 17566 4509 17600 4543
rect 17566 4441 17600 4475
rect 17566 4373 17600 4407
rect 17566 4305 17600 4339
rect 17566 4237 17600 4271
rect 17566 4169 17600 4203
rect 17662 5053 17696 5087
rect 17662 4985 17696 5019
rect 17662 4917 17696 4951
rect 17662 4849 17696 4883
rect 17662 4781 17696 4815
rect 17662 4713 17696 4747
rect 17662 4645 17696 4679
rect 17662 4577 17696 4611
rect 17662 4509 17696 4543
rect 17662 4441 17696 4475
rect 17662 4373 17696 4407
rect 17662 4305 17696 4339
rect 17662 4237 17696 4271
rect 17662 4169 17696 4203
rect 17758 5053 17792 5087
rect 17758 4985 17792 5019
rect 17758 4917 17792 4951
rect 17758 4849 17792 4883
rect 17758 4781 17792 4815
rect 17758 4713 17792 4747
rect 17758 4645 17792 4679
rect 17758 4577 17792 4611
rect 17758 4509 17792 4543
rect 17758 4441 17792 4475
rect 17758 4373 17792 4407
rect 17758 4305 17792 4339
rect 17758 4237 17792 4271
rect 17758 4169 17792 4203
rect 17854 5053 17888 5087
rect 17854 4985 17888 5019
rect 17854 4917 17888 4951
rect 17854 4849 17888 4883
rect 17854 4781 17888 4815
rect 17854 4713 17888 4747
rect 17854 4645 17888 4679
rect 17854 4577 17888 4611
rect 17854 4509 17888 4543
rect 17854 4441 17888 4475
rect 17854 4373 17888 4407
rect 17854 4305 17888 4339
rect 17854 4237 17888 4271
rect 17854 4169 17888 4203
rect 17950 5053 17984 5087
rect 17950 4985 17984 5019
rect 17950 4917 17984 4951
rect 17950 4849 17984 4883
rect 17950 4781 17984 4815
rect 17950 4713 17984 4747
rect 17950 4645 17984 4679
rect 17950 4577 17984 4611
rect 17950 4509 17984 4543
rect 17950 4441 17984 4475
rect 17950 4373 17984 4407
rect 17950 4305 17984 4339
rect 17950 4237 17984 4271
rect 17950 4169 17984 4203
rect 18046 5053 18080 5087
rect 18046 4985 18080 5019
rect 18046 4917 18080 4951
rect 18046 4849 18080 4883
rect 18046 4781 18080 4815
rect 18046 4713 18080 4747
rect 18046 4645 18080 4679
rect 18046 4577 18080 4611
rect 18046 4509 18080 4543
rect 18046 4441 18080 4475
rect 18046 4373 18080 4407
rect 18046 4305 18080 4339
rect 18046 4237 18080 4271
rect 18046 4169 18080 4203
rect 18142 5053 18176 5087
rect 18142 4985 18176 5019
rect 18142 4917 18176 4951
rect 18142 4849 18176 4883
rect 18142 4781 18176 4815
rect 18142 4713 18176 4747
rect 18142 4645 18176 4679
rect 18142 4577 18176 4611
rect 18142 4509 18176 4543
rect 18142 4441 18176 4475
rect 18142 4373 18176 4407
rect 18142 4305 18176 4339
rect 18142 4237 18176 4271
rect 18142 4169 18176 4203
rect 18238 5053 18272 5087
rect 18238 4985 18272 5019
rect 18238 4917 18272 4951
rect 18238 4849 18272 4883
rect 18238 4781 18272 4815
rect 18238 4713 18272 4747
rect 18238 4645 18272 4679
rect 18238 4577 18272 4611
rect 18238 4509 18272 4543
rect 18238 4441 18272 4475
rect 18238 4373 18272 4407
rect 18238 4305 18272 4339
rect 18238 4237 18272 4271
rect 18238 4169 18272 4203
rect 18334 5053 18368 5087
rect 18334 4985 18368 5019
rect 18334 4917 18368 4951
rect 18334 4849 18368 4883
rect 18334 4781 18368 4815
rect 18334 4713 18368 4747
rect 18334 4645 18368 4679
rect 18334 4577 18368 4611
rect 18334 4509 18368 4543
rect 18334 4441 18368 4475
rect 18334 4373 18368 4407
rect 18334 4305 18368 4339
rect 18334 4237 18368 4271
rect 18334 4169 18368 4203
rect 18430 5053 18464 5087
rect 18430 4985 18464 5019
rect 18430 4917 18464 4951
rect 18430 4849 18464 4883
rect 18430 4781 18464 4815
rect 18430 4713 18464 4747
rect 18430 4645 18464 4679
rect 18430 4577 18464 4611
rect 18430 4509 18464 4543
rect 18430 4441 18464 4475
rect 18430 4373 18464 4407
rect 18430 4305 18464 4339
rect 18430 4237 18464 4271
rect 18430 4169 18464 4203
rect 18674 5047 18708 5081
rect 18674 4979 18708 5013
rect 18674 4911 18708 4945
rect 18674 4843 18708 4877
rect 18674 4775 18708 4809
rect 18674 4707 18708 4741
rect 18674 4639 18708 4673
rect 18674 4571 18708 4605
rect 18674 4503 18708 4537
rect 18674 4435 18708 4469
rect 18674 4367 18708 4401
rect 18674 4299 18708 4333
rect 18674 4231 18708 4265
rect 18674 4163 18708 4197
rect 18770 5047 18804 5081
rect 18770 4979 18804 5013
rect 18770 4911 18804 4945
rect 18770 4843 18804 4877
rect 18770 4775 18804 4809
rect 18770 4707 18804 4741
rect 18770 4639 18804 4673
rect 18770 4571 18804 4605
rect 18770 4503 18804 4537
rect 18770 4435 18804 4469
rect 18770 4367 18804 4401
rect 18770 4299 18804 4333
rect 18770 4231 18804 4265
rect 18770 4163 18804 4197
rect 18866 5047 18900 5081
rect 18866 4979 18900 5013
rect 18866 4911 18900 4945
rect 18866 4843 18900 4877
rect 18866 4775 18900 4809
rect 18866 4707 18900 4741
rect 18866 4639 18900 4673
rect 18866 4571 18900 4605
rect 18866 4503 18900 4537
rect 18866 4435 18900 4469
rect 18866 4367 18900 4401
rect 18866 4299 18900 4333
rect 18866 4231 18900 4265
rect 18866 4163 18900 4197
rect 18962 5047 18996 5081
rect 18962 4979 18996 5013
rect 18962 4911 18996 4945
rect 18962 4843 18996 4877
rect 18962 4775 18996 4809
rect 18962 4707 18996 4741
rect 18962 4639 18996 4673
rect 18962 4571 18996 4605
rect 18962 4503 18996 4537
rect 18962 4435 18996 4469
rect 18962 4367 18996 4401
rect 18962 4299 18996 4333
rect 18962 4231 18996 4265
rect 18962 4163 18996 4197
rect 19058 5047 19092 5081
rect 19058 4979 19092 5013
rect 19058 4911 19092 4945
rect 19058 4843 19092 4877
rect 19058 4775 19092 4809
rect 19058 4707 19092 4741
rect 19058 4639 19092 4673
rect 19058 4571 19092 4605
rect 19058 4503 19092 4537
rect 19058 4435 19092 4469
rect 19058 4367 19092 4401
rect 19058 4299 19092 4333
rect 19058 4231 19092 4265
rect 19058 4163 19092 4197
rect 19154 5047 19188 5081
rect 19154 4979 19188 5013
rect 19154 4911 19188 4945
rect 19154 4843 19188 4877
rect 19154 4775 19188 4809
rect 19154 4707 19188 4741
rect 19154 4639 19188 4673
rect 19154 4571 19188 4605
rect 19154 4503 19188 4537
rect 19154 4435 19188 4469
rect 19154 4367 19188 4401
rect 19154 4299 19188 4333
rect 19154 4231 19188 4265
rect 19154 4163 19188 4197
rect 19250 5047 19284 5081
rect 19250 4979 19284 5013
rect 19250 4911 19284 4945
rect 19250 4843 19284 4877
rect 19250 4775 19284 4809
rect 19250 4707 19284 4741
rect 19250 4639 19284 4673
rect 19250 4571 19284 4605
rect 19250 4503 19284 4537
rect 19250 4435 19284 4469
rect 19250 4367 19284 4401
rect 19250 4299 19284 4333
rect 19250 4231 19284 4265
rect 19250 4163 19284 4197
rect 19346 5047 19380 5081
rect 19346 4979 19380 5013
rect 19346 4911 19380 4945
rect 19346 4843 19380 4877
rect 19346 4775 19380 4809
rect 19346 4707 19380 4741
rect 19346 4639 19380 4673
rect 19346 4571 19380 4605
rect 19346 4503 19380 4537
rect 19346 4435 19380 4469
rect 19346 4367 19380 4401
rect 19346 4299 19380 4333
rect 19346 4231 19380 4265
rect 19346 4163 19380 4197
rect 19442 5047 19476 5081
rect 19442 4979 19476 5013
rect 19442 4911 19476 4945
rect 19442 4843 19476 4877
rect 19442 4775 19476 4809
rect 19442 4707 19476 4741
rect 19442 4639 19476 4673
rect 19442 4571 19476 4605
rect 19442 4503 19476 4537
rect 19442 4435 19476 4469
rect 19442 4367 19476 4401
rect 19442 4299 19476 4333
rect 19442 4231 19476 4265
rect 19442 4163 19476 4197
rect 19538 5047 19572 5081
rect 19538 4979 19572 5013
rect 19538 4911 19572 4945
rect 19538 4843 19572 4877
rect 19538 4775 19572 4809
rect 19538 4707 19572 4741
rect 19538 4639 19572 4673
rect 19538 4571 19572 4605
rect 19538 4503 19572 4537
rect 19538 4435 19572 4469
rect 19538 4367 19572 4401
rect 19538 4299 19572 4333
rect 19538 4231 19572 4265
rect 19538 4163 19572 4197
rect 19634 5047 19668 5081
rect 19634 4979 19668 5013
rect 19634 4911 19668 4945
rect 19634 4843 19668 4877
rect 19634 4775 19668 4809
rect 19634 4707 19668 4741
rect 19634 4639 19668 4673
rect 19634 4571 19668 4605
rect 19634 4503 19668 4537
rect 19634 4435 19668 4469
rect 19634 4367 19668 4401
rect 19634 4299 19668 4333
rect 19634 4231 19668 4265
rect 19634 4163 19668 4197
rect 19730 5047 19764 5081
rect 19730 4979 19764 5013
rect 19730 4911 19764 4945
rect 19730 4843 19764 4877
rect 19730 4775 19764 4809
rect 19730 4707 19764 4741
rect 19730 4639 19764 4673
rect 19730 4571 19764 4605
rect 19730 4503 19764 4537
rect 19730 4435 19764 4469
rect 19730 4367 19764 4401
rect 19730 4299 19764 4333
rect 19730 4231 19764 4265
rect 19730 4163 19764 4197
rect 19826 5047 19860 5081
rect 19826 4979 19860 5013
rect 19826 4911 19860 4945
rect 19826 4843 19860 4877
rect 19826 4775 19860 4809
rect 19826 4707 19860 4741
rect 19826 4639 19860 4673
rect 19826 4571 19860 4605
rect 19826 4503 19860 4537
rect 19826 4435 19860 4469
rect 19826 4367 19860 4401
rect 19826 4299 19860 4333
rect 19826 4231 19860 4265
rect 19826 4163 19860 4197
rect 19922 5047 19956 5081
rect 19922 4979 19956 5013
rect 19922 4911 19956 4945
rect 19922 4843 19956 4877
rect 19922 4775 19956 4809
rect 19922 4707 19956 4741
rect 19922 4639 19956 4673
rect 19922 4571 19956 4605
rect 19922 4503 19956 4537
rect 19922 4435 19956 4469
rect 19922 4367 19956 4401
rect 19922 4299 19956 4333
rect 19922 4231 19956 4265
rect 19922 4163 19956 4197
rect 20018 5047 20052 5081
rect 20018 4979 20052 5013
rect 20018 4911 20052 4945
rect 20018 4843 20052 4877
rect 20018 4775 20052 4809
rect 20018 4707 20052 4741
rect 20018 4639 20052 4673
rect 20018 4571 20052 4605
rect 20018 4503 20052 4537
rect 20018 4435 20052 4469
rect 20018 4367 20052 4401
rect 20018 4299 20052 4333
rect 20018 4231 20052 4265
rect 20018 4163 20052 4197
rect 20114 5047 20148 5081
rect 20114 4979 20148 5013
rect 20114 4911 20148 4945
rect 20114 4843 20148 4877
rect 20114 4775 20148 4809
rect 20114 4707 20148 4741
rect 20114 4639 20148 4673
rect 20114 4571 20148 4605
rect 20114 4503 20148 4537
rect 20114 4435 20148 4469
rect 20114 4367 20148 4401
rect 20114 4299 20148 4333
rect 20114 4231 20148 4265
rect 20114 4163 20148 4197
rect 20338 5041 20372 5075
rect 20338 4973 20372 5007
rect 20338 4905 20372 4939
rect 20338 4837 20372 4871
rect 20338 4769 20372 4803
rect 20338 4701 20372 4735
rect 20338 4633 20372 4667
rect 20338 4565 20372 4599
rect 20338 4497 20372 4531
rect 20338 4429 20372 4463
rect 20338 4361 20372 4395
rect 20338 4293 20372 4327
rect 20338 4225 20372 4259
rect 20338 4157 20372 4191
rect 20434 5041 20468 5075
rect 20434 4973 20468 5007
rect 20434 4905 20468 4939
rect 20434 4837 20468 4871
rect 20434 4769 20468 4803
rect 20434 4701 20468 4735
rect 20434 4633 20468 4667
rect 20434 4565 20468 4599
rect 20434 4497 20468 4531
rect 20434 4429 20468 4463
rect 20434 4361 20468 4395
rect 20434 4293 20468 4327
rect 20434 4225 20468 4259
rect 20434 4157 20468 4191
rect 20530 5041 20564 5075
rect 20530 4973 20564 5007
rect 20530 4905 20564 4939
rect 20530 4837 20564 4871
rect 20530 4769 20564 4803
rect 20530 4701 20564 4735
rect 20530 4633 20564 4667
rect 20530 4565 20564 4599
rect 20530 4497 20564 4531
rect 20530 4429 20564 4463
rect 20530 4361 20564 4395
rect 20530 4293 20564 4327
rect 20530 4225 20564 4259
rect 20530 4157 20564 4191
rect 20626 5041 20660 5075
rect 20626 4973 20660 5007
rect 20626 4905 20660 4939
rect 20626 4837 20660 4871
rect 20626 4769 20660 4803
rect 20626 4701 20660 4735
rect 20626 4633 20660 4667
rect 20626 4565 20660 4599
rect 20626 4497 20660 4531
rect 20626 4429 20660 4463
rect 20626 4361 20660 4395
rect 20626 4293 20660 4327
rect 20626 4225 20660 4259
rect 20626 4157 20660 4191
rect 20722 5041 20756 5075
rect 20722 4973 20756 5007
rect 20722 4905 20756 4939
rect 20722 4837 20756 4871
rect 20722 4769 20756 4803
rect 20722 4701 20756 4735
rect 20722 4633 20756 4667
rect 20722 4565 20756 4599
rect 20722 4497 20756 4531
rect 20722 4429 20756 4463
rect 20722 4361 20756 4395
rect 20722 4293 20756 4327
rect 20722 4225 20756 4259
rect 20722 4157 20756 4191
rect 20818 5041 20852 5075
rect 20818 4973 20852 5007
rect 20818 4905 20852 4939
rect 20818 4837 20852 4871
rect 20818 4769 20852 4803
rect 20818 4701 20852 4735
rect 20818 4633 20852 4667
rect 20818 4565 20852 4599
rect 20818 4497 20852 4531
rect 20818 4429 20852 4463
rect 20818 4361 20852 4395
rect 20818 4293 20852 4327
rect 20818 4225 20852 4259
rect 20818 4157 20852 4191
rect 20914 5041 20948 5075
rect 20914 4973 20948 5007
rect 20914 4905 20948 4939
rect 20914 4837 20948 4871
rect 20914 4769 20948 4803
rect 20914 4701 20948 4735
rect 20914 4633 20948 4667
rect 20914 4565 20948 4599
rect 20914 4497 20948 4531
rect 20914 4429 20948 4463
rect 20914 4361 20948 4395
rect 20914 4293 20948 4327
rect 20914 4225 20948 4259
rect 20914 4157 20948 4191
rect 21010 5041 21044 5075
rect 21010 4973 21044 5007
rect 21010 4905 21044 4939
rect 21010 4837 21044 4871
rect 21010 4769 21044 4803
rect 21010 4701 21044 4735
rect 21010 4633 21044 4667
rect 21010 4565 21044 4599
rect 21010 4497 21044 4531
rect 21010 4429 21044 4463
rect 21010 4361 21044 4395
rect 21010 4293 21044 4327
rect 21010 4225 21044 4259
rect 21010 4157 21044 4191
rect 21106 5041 21140 5075
rect 21106 4973 21140 5007
rect 21106 4905 21140 4939
rect 21106 4837 21140 4871
rect 21106 4769 21140 4803
rect 21106 4701 21140 4735
rect 21106 4633 21140 4667
rect 21106 4565 21140 4599
rect 21106 4497 21140 4531
rect 21106 4429 21140 4463
rect 21106 4361 21140 4395
rect 21106 4293 21140 4327
rect 21106 4225 21140 4259
rect 21106 4157 21140 4191
rect 21202 5041 21236 5075
rect 21202 4973 21236 5007
rect 21202 4905 21236 4939
rect 21202 4837 21236 4871
rect 21202 4769 21236 4803
rect 21202 4701 21236 4735
rect 21202 4633 21236 4667
rect 21202 4565 21236 4599
rect 21202 4497 21236 4531
rect 21202 4429 21236 4463
rect 21202 4361 21236 4395
rect 21202 4293 21236 4327
rect 21202 4225 21236 4259
rect 21202 4157 21236 4191
rect 21298 5041 21332 5075
rect 21298 4973 21332 5007
rect 21298 4905 21332 4939
rect 21298 4837 21332 4871
rect 21298 4769 21332 4803
rect 21298 4701 21332 4735
rect 21298 4633 21332 4667
rect 21298 4565 21332 4599
rect 21298 4497 21332 4531
rect 21298 4429 21332 4463
rect 21298 4361 21332 4395
rect 21298 4293 21332 4327
rect 21298 4225 21332 4259
rect 21298 4157 21332 4191
rect 21394 5041 21428 5075
rect 21394 4973 21428 5007
rect 21394 4905 21428 4939
rect 21394 4837 21428 4871
rect 21394 4769 21428 4803
rect 21394 4701 21428 4735
rect 21394 4633 21428 4667
rect 21394 4565 21428 4599
rect 21394 4497 21428 4531
rect 21394 4429 21428 4463
rect 21394 4361 21428 4395
rect 21394 4293 21428 4327
rect 21394 4225 21428 4259
rect 21394 4157 21428 4191
rect 21490 5041 21524 5075
rect 21490 4973 21524 5007
rect 21490 4905 21524 4939
rect 21490 4837 21524 4871
rect 21490 4769 21524 4803
rect 21490 4701 21524 4735
rect 21490 4633 21524 4667
rect 21490 4565 21524 4599
rect 21490 4497 21524 4531
rect 21490 4429 21524 4463
rect 21490 4361 21524 4395
rect 21490 4293 21524 4327
rect 21490 4225 21524 4259
rect 21490 4157 21524 4191
rect 21586 5041 21620 5075
rect 21586 4973 21620 5007
rect 21586 4905 21620 4939
rect 21586 4837 21620 4871
rect 21586 4769 21620 4803
rect 21586 4701 21620 4735
rect 21586 4633 21620 4667
rect 21586 4565 21620 4599
rect 21586 4497 21620 4531
rect 21586 4429 21620 4463
rect 21586 4361 21620 4395
rect 21586 4293 21620 4327
rect 21586 4225 21620 4259
rect 21586 4157 21620 4191
rect 21682 5041 21716 5075
rect 21682 4973 21716 5007
rect 21682 4905 21716 4939
rect 21682 4837 21716 4871
rect 21682 4769 21716 4803
rect 21682 4701 21716 4735
rect 21682 4633 21716 4667
rect 21682 4565 21716 4599
rect 21682 4497 21716 4531
rect 21682 4429 21716 4463
rect 21682 4361 21716 4395
rect 21682 4293 21716 4327
rect 21682 4225 21716 4259
rect 21682 4157 21716 4191
rect 21778 5041 21812 5075
rect 21778 4973 21812 5007
rect 21778 4905 21812 4939
rect 21778 4837 21812 4871
rect 21778 4769 21812 4803
rect 21778 4701 21812 4735
rect 21778 4633 21812 4667
rect 21778 4565 21812 4599
rect 21778 4497 21812 4531
rect 21778 4429 21812 4463
rect 21778 4361 21812 4395
rect 21778 4293 21812 4327
rect 21778 4225 21812 4259
rect 21778 4157 21812 4191
rect 21874 5041 21908 5075
rect 21874 4973 21908 5007
rect 21874 4905 21908 4939
rect 21874 4837 21908 4871
rect 21874 4769 21908 4803
rect 21874 4701 21908 4735
rect 21874 4633 21908 4667
rect 21874 4565 21908 4599
rect 21874 4497 21908 4531
rect 21874 4429 21908 4463
rect 21874 4361 21908 4395
rect 21874 4293 21908 4327
rect 21874 4225 21908 4259
rect 21874 4157 21908 4191
rect 21970 5041 22004 5075
rect 21970 4973 22004 5007
rect 21970 4905 22004 4939
rect 21970 4837 22004 4871
rect 21970 4769 22004 4803
rect 21970 4701 22004 4735
rect 21970 4633 22004 4667
rect 21970 4565 22004 4599
rect 21970 4497 22004 4531
rect 21970 4429 22004 4463
rect 21970 4361 22004 4395
rect 21970 4293 22004 4327
rect 21970 4225 22004 4259
rect 21970 4157 22004 4191
rect 22066 5041 22100 5075
rect 22066 4973 22100 5007
rect 22066 4905 22100 4939
rect 22066 4837 22100 4871
rect 22066 4769 22100 4803
rect 22066 4701 22100 4735
rect 22066 4633 22100 4667
rect 22066 4565 22100 4599
rect 22066 4497 22100 4531
rect 22066 4429 22100 4463
rect 22066 4361 22100 4395
rect 22066 4293 22100 4327
rect 22066 4225 22100 4259
rect 22066 4157 22100 4191
rect 22162 5041 22196 5075
rect 22162 4973 22196 5007
rect 22162 4905 22196 4939
rect 22162 4837 22196 4871
rect 22162 4769 22196 4803
rect 22162 4701 22196 4735
rect 22162 4633 22196 4667
rect 22162 4565 22196 4599
rect 22162 4497 22196 4531
rect 22162 4429 22196 4463
rect 22162 4361 22196 4395
rect 22162 4293 22196 4327
rect 22162 4225 22196 4259
rect 22162 4157 22196 4191
rect 22258 5041 22292 5075
rect 22258 4973 22292 5007
rect 22258 4905 22292 4939
rect 22258 4837 22292 4871
rect 22258 4769 22292 4803
rect 22258 4701 22292 4735
rect 22258 4633 22292 4667
rect 22258 4565 22292 4599
rect 22258 4497 22292 4531
rect 22258 4429 22292 4463
rect 22258 4361 22292 4395
rect 22258 4293 22292 4327
rect 22258 4225 22292 4259
rect 22258 4157 22292 4191
rect 23270 5053 23304 5087
rect 23270 4985 23304 5019
rect 23270 4917 23304 4951
rect 23270 4849 23304 4883
rect 23270 4781 23304 4815
rect 23270 4713 23304 4747
rect 23270 4645 23304 4679
rect 23270 4577 23304 4611
rect 23270 4509 23304 4543
rect 23270 4441 23304 4475
rect 23270 4373 23304 4407
rect 23270 4305 23304 4339
rect 23270 4237 23304 4271
rect 23270 4169 23304 4203
rect 23366 5053 23400 5087
rect 23366 4985 23400 5019
rect 23366 4917 23400 4951
rect 23366 4849 23400 4883
rect 23366 4781 23400 4815
rect 23366 4713 23400 4747
rect 23366 4645 23400 4679
rect 23366 4577 23400 4611
rect 23366 4509 23400 4543
rect 23366 4441 23400 4475
rect 23366 4373 23400 4407
rect 23366 4305 23400 4339
rect 23366 4237 23400 4271
rect 23366 4169 23400 4203
rect 23462 5053 23496 5087
rect 23462 4985 23496 5019
rect 23462 4917 23496 4951
rect 23462 4849 23496 4883
rect 23462 4781 23496 4815
rect 23462 4713 23496 4747
rect 23462 4645 23496 4679
rect 23462 4577 23496 4611
rect 23462 4509 23496 4543
rect 23462 4441 23496 4475
rect 23462 4373 23496 4407
rect 23462 4305 23496 4339
rect 23462 4237 23496 4271
rect 23462 4169 23496 4203
rect 23558 5053 23592 5087
rect 23558 4985 23592 5019
rect 23558 4917 23592 4951
rect 23558 4849 23592 4883
rect 23558 4781 23592 4815
rect 23558 4713 23592 4747
rect 23558 4645 23592 4679
rect 23558 4577 23592 4611
rect 23558 4509 23592 4543
rect 23558 4441 23592 4475
rect 23558 4373 23592 4407
rect 23558 4305 23592 4339
rect 23558 4237 23592 4271
rect 23558 4169 23592 4203
rect 23654 5053 23688 5087
rect 23654 4985 23688 5019
rect 23654 4917 23688 4951
rect 23654 4849 23688 4883
rect 23654 4781 23688 4815
rect 23654 4713 23688 4747
rect 23654 4645 23688 4679
rect 23654 4577 23688 4611
rect 23654 4509 23688 4543
rect 23654 4441 23688 4475
rect 23654 4373 23688 4407
rect 23654 4305 23688 4339
rect 23654 4237 23688 4271
rect 23654 4169 23688 4203
rect 23750 5053 23784 5087
rect 23750 4985 23784 5019
rect 23750 4917 23784 4951
rect 23750 4849 23784 4883
rect 23750 4781 23784 4815
rect 23750 4713 23784 4747
rect 23750 4645 23784 4679
rect 23750 4577 23784 4611
rect 23750 4509 23784 4543
rect 23750 4441 23784 4475
rect 23750 4373 23784 4407
rect 23750 4305 23784 4339
rect 23750 4237 23784 4271
rect 23750 4169 23784 4203
rect 23958 5051 23992 5085
rect 23958 4983 23992 5017
rect 23958 4915 23992 4949
rect 23958 4847 23992 4881
rect 23958 4779 23992 4813
rect 23958 4711 23992 4745
rect 23958 4643 23992 4677
rect 23958 4575 23992 4609
rect 23958 4507 23992 4541
rect 23958 4439 23992 4473
rect 23958 4371 23992 4405
rect 23958 4303 23992 4337
rect 23958 4235 23992 4269
rect 23958 4167 23992 4201
rect 24054 5051 24088 5085
rect 24054 4983 24088 5017
rect 24054 4915 24088 4949
rect 24054 4847 24088 4881
rect 24054 4779 24088 4813
rect 24054 4711 24088 4745
rect 24054 4643 24088 4677
rect 24054 4575 24088 4609
rect 24054 4507 24088 4541
rect 24054 4439 24088 4473
rect 24054 4371 24088 4405
rect 24054 4303 24088 4337
rect 24054 4235 24088 4269
rect 24054 4167 24088 4201
rect 24150 5051 24184 5085
rect 24150 4983 24184 5017
rect 24150 4915 24184 4949
rect 24150 4847 24184 4881
rect 24150 4779 24184 4813
rect 24150 4711 24184 4745
rect 24150 4643 24184 4677
rect 24150 4575 24184 4609
rect 24150 4507 24184 4541
rect 24150 4439 24184 4473
rect 24150 4371 24184 4405
rect 24150 4303 24184 4337
rect 24150 4235 24184 4269
rect 24150 4167 24184 4201
rect 24246 5051 24280 5085
rect 24246 4983 24280 5017
rect 24246 4915 24280 4949
rect 24246 4847 24280 4881
rect 24246 4779 24280 4813
rect 24246 4711 24280 4745
rect 24246 4643 24280 4677
rect 24246 4575 24280 4609
rect 24246 4507 24280 4541
rect 24246 4439 24280 4473
rect 24246 4371 24280 4405
rect 24246 4303 24280 4337
rect 24246 4235 24280 4269
rect 24246 4167 24280 4201
rect 24342 5051 24376 5085
rect 24342 4983 24376 5017
rect 24342 4915 24376 4949
rect 24342 4847 24376 4881
rect 24342 4779 24376 4813
rect 24342 4711 24376 4745
rect 24342 4643 24376 4677
rect 24342 4575 24376 4609
rect 24342 4507 24376 4541
rect 24342 4439 24376 4473
rect 24342 4371 24376 4405
rect 24342 4303 24376 4337
rect 24342 4235 24376 4269
rect 24342 4167 24376 4201
rect 24438 5051 24472 5085
rect 24438 4983 24472 5017
rect 24438 4915 24472 4949
rect 24438 4847 24472 4881
rect 24438 4779 24472 4813
rect 24438 4711 24472 4745
rect 24438 4643 24472 4677
rect 24438 4575 24472 4609
rect 24438 4507 24472 4541
rect 24438 4439 24472 4473
rect 24438 4371 24472 4405
rect 24438 4303 24472 4337
rect 24438 4235 24472 4269
rect 24438 4167 24472 4201
rect 24534 5051 24568 5085
rect 24534 4983 24568 5017
rect 24534 4915 24568 4949
rect 24534 4847 24568 4881
rect 24534 4779 24568 4813
rect 24534 4711 24568 4745
rect 24534 4643 24568 4677
rect 24534 4575 24568 4609
rect 24534 4507 24568 4541
rect 24534 4439 24568 4473
rect 24534 4371 24568 4405
rect 24534 4303 24568 4337
rect 24534 4235 24568 4269
rect 24534 4167 24568 4201
rect 24630 5051 24664 5085
rect 24630 4983 24664 5017
rect 24630 4915 24664 4949
rect 24630 4847 24664 4881
rect 24630 4779 24664 4813
rect 24630 4711 24664 4745
rect 24630 4643 24664 4677
rect 24630 4575 24664 4609
rect 24630 4507 24664 4541
rect 24630 4439 24664 4473
rect 24630 4371 24664 4405
rect 24630 4303 24664 4337
rect 24630 4235 24664 4269
rect 24630 4167 24664 4201
rect 24726 5051 24760 5085
rect 24726 4983 24760 5017
rect 24726 4915 24760 4949
rect 24726 4847 24760 4881
rect 24726 4779 24760 4813
rect 24726 4711 24760 4745
rect 24726 4643 24760 4677
rect 24726 4575 24760 4609
rect 24726 4507 24760 4541
rect 24726 4439 24760 4473
rect 24726 4371 24760 4405
rect 24726 4303 24760 4337
rect 24726 4235 24760 4269
rect 24726 4167 24760 4201
rect 24822 5051 24856 5085
rect 24822 4983 24856 5017
rect 24822 4915 24856 4949
rect 24822 4847 24856 4881
rect 24822 4779 24856 4813
rect 24822 4711 24856 4745
rect 24822 4643 24856 4677
rect 24822 4575 24856 4609
rect 24822 4507 24856 4541
rect 24822 4439 24856 4473
rect 24822 4371 24856 4405
rect 24822 4303 24856 4337
rect 24822 4235 24856 4269
rect 24822 4167 24856 4201
rect 24918 5051 24952 5085
rect 24918 4983 24952 5017
rect 24918 4915 24952 4949
rect 24918 4847 24952 4881
rect 24918 4779 24952 4813
rect 24918 4711 24952 4745
rect 24918 4643 24952 4677
rect 24918 4575 24952 4609
rect 24918 4507 24952 4541
rect 24918 4439 24952 4473
rect 24918 4371 24952 4405
rect 24918 4303 24952 4337
rect 24918 4235 24952 4269
rect 24918 4167 24952 4201
rect 25162 5045 25196 5079
rect 25162 4977 25196 5011
rect 25162 4909 25196 4943
rect 25162 4841 25196 4875
rect 25162 4773 25196 4807
rect 25162 4705 25196 4739
rect 25162 4637 25196 4671
rect 25162 4569 25196 4603
rect 25162 4501 25196 4535
rect 25162 4433 25196 4467
rect 25162 4365 25196 4399
rect 25162 4297 25196 4331
rect 25162 4229 25196 4263
rect 25162 4161 25196 4195
rect 25258 5045 25292 5079
rect 25258 4977 25292 5011
rect 25258 4909 25292 4943
rect 25258 4841 25292 4875
rect 25258 4773 25292 4807
rect 25258 4705 25292 4739
rect 25258 4637 25292 4671
rect 25258 4569 25292 4603
rect 25258 4501 25292 4535
rect 25258 4433 25292 4467
rect 25258 4365 25292 4399
rect 25258 4297 25292 4331
rect 25258 4229 25292 4263
rect 25258 4161 25292 4195
rect 25354 5045 25388 5079
rect 25354 4977 25388 5011
rect 25354 4909 25388 4943
rect 25354 4841 25388 4875
rect 25354 4773 25388 4807
rect 25354 4705 25388 4739
rect 25354 4637 25388 4671
rect 25354 4569 25388 4603
rect 25354 4501 25388 4535
rect 25354 4433 25388 4467
rect 25354 4365 25388 4399
rect 25354 4297 25388 4331
rect 25354 4229 25388 4263
rect 25354 4161 25388 4195
rect 25450 5045 25484 5079
rect 25450 4977 25484 5011
rect 25450 4909 25484 4943
rect 25450 4841 25484 4875
rect 25450 4773 25484 4807
rect 25450 4705 25484 4739
rect 25450 4637 25484 4671
rect 25450 4569 25484 4603
rect 25450 4501 25484 4535
rect 25450 4433 25484 4467
rect 25450 4365 25484 4399
rect 25450 4297 25484 4331
rect 25450 4229 25484 4263
rect 25450 4161 25484 4195
rect 25546 5045 25580 5079
rect 25546 4977 25580 5011
rect 25546 4909 25580 4943
rect 25546 4841 25580 4875
rect 25546 4773 25580 4807
rect 25546 4705 25580 4739
rect 25546 4637 25580 4671
rect 25546 4569 25580 4603
rect 25546 4501 25580 4535
rect 25546 4433 25580 4467
rect 25546 4365 25580 4399
rect 25546 4297 25580 4331
rect 25546 4229 25580 4263
rect 25546 4161 25580 4195
rect 25642 5045 25676 5079
rect 25642 4977 25676 5011
rect 25642 4909 25676 4943
rect 25642 4841 25676 4875
rect 25642 4773 25676 4807
rect 25642 4705 25676 4739
rect 25642 4637 25676 4671
rect 25642 4569 25676 4603
rect 25642 4501 25676 4535
rect 25642 4433 25676 4467
rect 25642 4365 25676 4399
rect 25642 4297 25676 4331
rect 25642 4229 25676 4263
rect 25642 4161 25676 4195
rect 25738 5045 25772 5079
rect 25738 4977 25772 5011
rect 25738 4909 25772 4943
rect 25738 4841 25772 4875
rect 25738 4773 25772 4807
rect 25738 4705 25772 4739
rect 25738 4637 25772 4671
rect 25738 4569 25772 4603
rect 25738 4501 25772 4535
rect 25738 4433 25772 4467
rect 25738 4365 25772 4399
rect 25738 4297 25772 4331
rect 25738 4229 25772 4263
rect 25738 4161 25772 4195
rect 25834 5045 25868 5079
rect 25834 4977 25868 5011
rect 25834 4909 25868 4943
rect 25834 4841 25868 4875
rect 25834 4773 25868 4807
rect 25834 4705 25868 4739
rect 25834 4637 25868 4671
rect 25834 4569 25868 4603
rect 25834 4501 25868 4535
rect 25834 4433 25868 4467
rect 25834 4365 25868 4399
rect 25834 4297 25868 4331
rect 25834 4229 25868 4263
rect 25834 4161 25868 4195
rect 25930 5045 25964 5079
rect 25930 4977 25964 5011
rect 25930 4909 25964 4943
rect 25930 4841 25964 4875
rect 25930 4773 25964 4807
rect 25930 4705 25964 4739
rect 25930 4637 25964 4671
rect 25930 4569 25964 4603
rect 25930 4501 25964 4535
rect 25930 4433 25964 4467
rect 25930 4365 25964 4399
rect 25930 4297 25964 4331
rect 25930 4229 25964 4263
rect 25930 4161 25964 4195
rect 26026 5045 26060 5079
rect 26026 4977 26060 5011
rect 26026 4909 26060 4943
rect 26026 4841 26060 4875
rect 26026 4773 26060 4807
rect 26026 4705 26060 4739
rect 26026 4637 26060 4671
rect 26026 4569 26060 4603
rect 26026 4501 26060 4535
rect 26026 4433 26060 4467
rect 26026 4365 26060 4399
rect 26026 4297 26060 4331
rect 26026 4229 26060 4263
rect 26026 4161 26060 4195
rect 26122 5045 26156 5079
rect 26122 4977 26156 5011
rect 26122 4909 26156 4943
rect 26122 4841 26156 4875
rect 26122 4773 26156 4807
rect 26122 4705 26156 4739
rect 26122 4637 26156 4671
rect 26122 4569 26156 4603
rect 26122 4501 26156 4535
rect 26122 4433 26156 4467
rect 26122 4365 26156 4399
rect 26122 4297 26156 4331
rect 26122 4229 26156 4263
rect 26122 4161 26156 4195
rect 26218 5045 26252 5079
rect 26218 4977 26252 5011
rect 26218 4909 26252 4943
rect 26218 4841 26252 4875
rect 26218 4773 26252 4807
rect 26218 4705 26252 4739
rect 26218 4637 26252 4671
rect 26218 4569 26252 4603
rect 26218 4501 26252 4535
rect 26218 4433 26252 4467
rect 26218 4365 26252 4399
rect 26218 4297 26252 4331
rect 26218 4229 26252 4263
rect 26218 4161 26252 4195
rect 26314 5045 26348 5079
rect 26314 4977 26348 5011
rect 26314 4909 26348 4943
rect 26314 4841 26348 4875
rect 26314 4773 26348 4807
rect 26314 4705 26348 4739
rect 26314 4637 26348 4671
rect 26314 4569 26348 4603
rect 26314 4501 26348 4535
rect 26314 4433 26348 4467
rect 26314 4365 26348 4399
rect 26314 4297 26348 4331
rect 26314 4229 26348 4263
rect 26314 4161 26348 4195
rect 26410 5045 26444 5079
rect 26410 4977 26444 5011
rect 26410 4909 26444 4943
rect 26410 4841 26444 4875
rect 26410 4773 26444 4807
rect 26410 4705 26444 4739
rect 26410 4637 26444 4671
rect 26410 4569 26444 4603
rect 26410 4501 26444 4535
rect 26410 4433 26444 4467
rect 26410 4365 26444 4399
rect 26410 4297 26444 4331
rect 26410 4229 26444 4263
rect 26410 4161 26444 4195
rect 26506 5045 26540 5079
rect 26506 4977 26540 5011
rect 26506 4909 26540 4943
rect 26506 4841 26540 4875
rect 26506 4773 26540 4807
rect 26506 4705 26540 4739
rect 26506 4637 26540 4671
rect 26506 4569 26540 4603
rect 26506 4501 26540 4535
rect 26506 4433 26540 4467
rect 26506 4365 26540 4399
rect 26506 4297 26540 4331
rect 26506 4229 26540 4263
rect 26506 4161 26540 4195
rect 26602 5045 26636 5079
rect 26602 4977 26636 5011
rect 26602 4909 26636 4943
rect 26602 4841 26636 4875
rect 26602 4773 26636 4807
rect 26602 4705 26636 4739
rect 26602 4637 26636 4671
rect 26602 4569 26636 4603
rect 26602 4501 26636 4535
rect 26602 4433 26636 4467
rect 26602 4365 26636 4399
rect 26602 4297 26636 4331
rect 26602 4229 26636 4263
rect 26602 4161 26636 4195
rect 26826 5039 26860 5073
rect 26826 4971 26860 5005
rect 26826 4903 26860 4937
rect 26826 4835 26860 4869
rect 26826 4767 26860 4801
rect 26826 4699 26860 4733
rect 26826 4631 26860 4665
rect 26826 4563 26860 4597
rect 26826 4495 26860 4529
rect 26826 4427 26860 4461
rect 26826 4359 26860 4393
rect 26826 4291 26860 4325
rect 26826 4223 26860 4257
rect 26826 4155 26860 4189
rect 26922 5039 26956 5073
rect 26922 4971 26956 5005
rect 26922 4903 26956 4937
rect 26922 4835 26956 4869
rect 26922 4767 26956 4801
rect 26922 4699 26956 4733
rect 26922 4631 26956 4665
rect 26922 4563 26956 4597
rect 26922 4495 26956 4529
rect 26922 4427 26956 4461
rect 26922 4359 26956 4393
rect 26922 4291 26956 4325
rect 26922 4223 26956 4257
rect 26922 4155 26956 4189
rect 27018 5039 27052 5073
rect 27018 4971 27052 5005
rect 27018 4903 27052 4937
rect 27018 4835 27052 4869
rect 27018 4767 27052 4801
rect 27018 4699 27052 4733
rect 27018 4631 27052 4665
rect 27018 4563 27052 4597
rect 27018 4495 27052 4529
rect 27018 4427 27052 4461
rect 27018 4359 27052 4393
rect 27018 4291 27052 4325
rect 27018 4223 27052 4257
rect 27018 4155 27052 4189
rect 27114 5039 27148 5073
rect 27114 4971 27148 5005
rect 27114 4903 27148 4937
rect 27114 4835 27148 4869
rect 27114 4767 27148 4801
rect 27114 4699 27148 4733
rect 27114 4631 27148 4665
rect 27114 4563 27148 4597
rect 27114 4495 27148 4529
rect 27114 4427 27148 4461
rect 27114 4359 27148 4393
rect 27114 4291 27148 4325
rect 27114 4223 27148 4257
rect 27114 4155 27148 4189
rect 27210 5039 27244 5073
rect 27210 4971 27244 5005
rect 27210 4903 27244 4937
rect 27210 4835 27244 4869
rect 27210 4767 27244 4801
rect 27210 4699 27244 4733
rect 27210 4631 27244 4665
rect 27210 4563 27244 4597
rect 27210 4495 27244 4529
rect 27210 4427 27244 4461
rect 27210 4359 27244 4393
rect 27210 4291 27244 4325
rect 27210 4223 27244 4257
rect 27210 4155 27244 4189
rect 27306 5039 27340 5073
rect 27306 4971 27340 5005
rect 27306 4903 27340 4937
rect 27306 4835 27340 4869
rect 27306 4767 27340 4801
rect 27306 4699 27340 4733
rect 27306 4631 27340 4665
rect 27306 4563 27340 4597
rect 27306 4495 27340 4529
rect 27306 4427 27340 4461
rect 27306 4359 27340 4393
rect 27306 4291 27340 4325
rect 27306 4223 27340 4257
rect 27306 4155 27340 4189
rect 27402 5039 27436 5073
rect 27402 4971 27436 5005
rect 27402 4903 27436 4937
rect 27402 4835 27436 4869
rect 27402 4767 27436 4801
rect 27402 4699 27436 4733
rect 27402 4631 27436 4665
rect 27402 4563 27436 4597
rect 27402 4495 27436 4529
rect 27402 4427 27436 4461
rect 27402 4359 27436 4393
rect 27402 4291 27436 4325
rect 27402 4223 27436 4257
rect 27402 4155 27436 4189
rect 27498 5039 27532 5073
rect 27498 4971 27532 5005
rect 27498 4903 27532 4937
rect 27498 4835 27532 4869
rect 27498 4767 27532 4801
rect 27498 4699 27532 4733
rect 27498 4631 27532 4665
rect 27498 4563 27532 4597
rect 27498 4495 27532 4529
rect 27498 4427 27532 4461
rect 27498 4359 27532 4393
rect 27498 4291 27532 4325
rect 27498 4223 27532 4257
rect 27498 4155 27532 4189
rect 27594 5039 27628 5073
rect 27594 4971 27628 5005
rect 27594 4903 27628 4937
rect 27594 4835 27628 4869
rect 27594 4767 27628 4801
rect 27594 4699 27628 4733
rect 27594 4631 27628 4665
rect 27594 4563 27628 4597
rect 27594 4495 27628 4529
rect 27594 4427 27628 4461
rect 27594 4359 27628 4393
rect 27594 4291 27628 4325
rect 27594 4223 27628 4257
rect 27594 4155 27628 4189
rect 27690 5039 27724 5073
rect 27690 4971 27724 5005
rect 27690 4903 27724 4937
rect 27690 4835 27724 4869
rect 27690 4767 27724 4801
rect 27690 4699 27724 4733
rect 27690 4631 27724 4665
rect 27690 4563 27724 4597
rect 27690 4495 27724 4529
rect 27690 4427 27724 4461
rect 27690 4359 27724 4393
rect 27690 4291 27724 4325
rect 27690 4223 27724 4257
rect 27690 4155 27724 4189
rect 27786 5039 27820 5073
rect 27786 4971 27820 5005
rect 27786 4903 27820 4937
rect 27786 4835 27820 4869
rect 27786 4767 27820 4801
rect 27786 4699 27820 4733
rect 27786 4631 27820 4665
rect 27786 4563 27820 4597
rect 27786 4495 27820 4529
rect 27786 4427 27820 4461
rect 27786 4359 27820 4393
rect 27786 4291 27820 4325
rect 27786 4223 27820 4257
rect 27786 4155 27820 4189
rect 27882 5039 27916 5073
rect 27882 4971 27916 5005
rect 27882 4903 27916 4937
rect 27882 4835 27916 4869
rect 27882 4767 27916 4801
rect 27882 4699 27916 4733
rect 27882 4631 27916 4665
rect 27882 4563 27916 4597
rect 27882 4495 27916 4529
rect 27882 4427 27916 4461
rect 27882 4359 27916 4393
rect 27882 4291 27916 4325
rect 27882 4223 27916 4257
rect 27882 4155 27916 4189
rect 27978 5039 28012 5073
rect 27978 4971 28012 5005
rect 27978 4903 28012 4937
rect 27978 4835 28012 4869
rect 27978 4767 28012 4801
rect 27978 4699 28012 4733
rect 27978 4631 28012 4665
rect 27978 4563 28012 4597
rect 27978 4495 28012 4529
rect 27978 4427 28012 4461
rect 27978 4359 28012 4393
rect 27978 4291 28012 4325
rect 27978 4223 28012 4257
rect 27978 4155 28012 4189
rect 28074 5039 28108 5073
rect 28074 4971 28108 5005
rect 28074 4903 28108 4937
rect 28074 4835 28108 4869
rect 28074 4767 28108 4801
rect 28074 4699 28108 4733
rect 28074 4631 28108 4665
rect 28074 4563 28108 4597
rect 28074 4495 28108 4529
rect 28074 4427 28108 4461
rect 28074 4359 28108 4393
rect 28074 4291 28108 4325
rect 28074 4223 28108 4257
rect 28074 4155 28108 4189
rect 28170 5039 28204 5073
rect 28170 4971 28204 5005
rect 28170 4903 28204 4937
rect 28170 4835 28204 4869
rect 28170 4767 28204 4801
rect 28170 4699 28204 4733
rect 28170 4631 28204 4665
rect 28170 4563 28204 4597
rect 28170 4495 28204 4529
rect 28170 4427 28204 4461
rect 28170 4359 28204 4393
rect 28170 4291 28204 4325
rect 28170 4223 28204 4257
rect 28170 4155 28204 4189
rect 28266 5039 28300 5073
rect 28266 4971 28300 5005
rect 28266 4903 28300 4937
rect 28266 4835 28300 4869
rect 28266 4767 28300 4801
rect 28266 4699 28300 4733
rect 28266 4631 28300 4665
rect 28266 4563 28300 4597
rect 28266 4495 28300 4529
rect 28266 4427 28300 4461
rect 28266 4359 28300 4393
rect 28266 4291 28300 4325
rect 28266 4223 28300 4257
rect 28266 4155 28300 4189
rect 28362 5039 28396 5073
rect 28362 4971 28396 5005
rect 28362 4903 28396 4937
rect 28362 4835 28396 4869
rect 28362 4767 28396 4801
rect 28362 4699 28396 4733
rect 28362 4631 28396 4665
rect 28362 4563 28396 4597
rect 28362 4495 28396 4529
rect 28362 4427 28396 4461
rect 28362 4359 28396 4393
rect 28362 4291 28396 4325
rect 28362 4223 28396 4257
rect 28362 4155 28396 4189
rect 28458 5039 28492 5073
rect 28458 4971 28492 5005
rect 28458 4903 28492 4937
rect 28458 4835 28492 4869
rect 28458 4767 28492 4801
rect 28458 4699 28492 4733
rect 28458 4631 28492 4665
rect 28458 4563 28492 4597
rect 28458 4495 28492 4529
rect 28458 4427 28492 4461
rect 28458 4359 28492 4393
rect 28458 4291 28492 4325
rect 28458 4223 28492 4257
rect 28458 4155 28492 4189
rect 28554 5039 28588 5073
rect 28554 4971 28588 5005
rect 28554 4903 28588 4937
rect 28554 4835 28588 4869
rect 28554 4767 28588 4801
rect 28554 4699 28588 4733
rect 28554 4631 28588 4665
rect 28554 4563 28588 4597
rect 28554 4495 28588 4529
rect 28554 4427 28588 4461
rect 28554 4359 28588 4393
rect 28554 4291 28588 4325
rect 28554 4223 28588 4257
rect 28554 4155 28588 4189
rect 28650 5039 28684 5073
rect 28650 4971 28684 5005
rect 28650 4903 28684 4937
rect 28650 4835 28684 4869
rect 28650 4767 28684 4801
rect 28650 4699 28684 4733
rect 28650 4631 28684 4665
rect 28650 4563 28684 4597
rect 28650 4495 28684 4529
rect 28650 4427 28684 4461
rect 28650 4359 28684 4393
rect 28650 4291 28684 4325
rect 28650 4223 28684 4257
rect 28650 4155 28684 4189
rect 28746 5039 28780 5073
rect 28746 4971 28780 5005
rect 28746 4903 28780 4937
rect 28746 4835 28780 4869
rect 28746 4767 28780 4801
rect 28746 4699 28780 4733
rect 28746 4631 28780 4665
rect 28746 4563 28780 4597
rect 28746 4495 28780 4529
rect 28746 4427 28780 4461
rect 28746 4359 28780 4393
rect 28746 4291 28780 4325
rect 28746 4223 28780 4257
rect 28746 4155 28780 4189
rect -4814 3643 -4780 3677
rect -4814 3575 -4780 3609
rect -4814 3507 -4780 3541
<< psubdiff >>
rect 16642 2334 22276 2342
rect 16642 2164 16688 2334
rect 22230 2164 22276 2334
rect 16642 2156 22276 2164
rect 23130 2332 28764 2340
rect 23130 2162 23176 2332
rect 28718 2162 28764 2332
rect 23130 2154 28764 2162
rect -16740 1672 -11106 1680
rect -23570 1660 -17936 1668
rect -23570 1490 -23524 1660
rect -17982 1490 -17936 1660
rect -16740 1502 -16694 1672
rect -11152 1502 -11106 1672
rect -16740 1494 -11106 1502
rect -10274 1670 -4640 1678
rect -10274 1500 -10228 1670
rect -4686 1500 -4640 1670
rect -10274 1492 -4640 1500
rect -23570 1482 -17936 1490
rect 250 -963 15780 -948
rect 250 -1269 280 -963
rect 15750 -1269 15780 -963
rect 250 -1284 15780 -1269
<< nsubdiff >>
rect -1372 8157 15840 8180
rect -1372 7851 -1317 8157
rect 15785 7851 15840 8157
rect -1372 7828 15840 7851
rect -23604 4805 -18086 4826
rect -23604 4635 -23548 4805
rect -18142 4635 -18086 4805
rect -23604 4614 -18086 4635
rect -16774 4817 -11256 4838
rect -16774 4647 -16718 4817
rect -11312 4647 -11256 4817
rect -16774 4626 -11256 4647
rect -10308 4815 -4790 4836
rect -10308 4645 -10252 4815
rect -4846 4645 -4790 4815
rect -10308 4624 -4790 4645
rect 16792 5479 22310 5500
rect 16792 5309 16848 5479
rect 22254 5309 22310 5479
rect 16792 5288 22310 5309
rect 23280 5477 28798 5498
rect 23280 5307 23336 5477
rect 28742 5307 28798 5477
rect 23280 5286 28798 5307
<< psubdiffcont >>
rect 16688 2164 22230 2334
rect 23176 2162 28718 2332
rect -23524 1490 -17982 1660
rect -16694 1502 -11152 1672
rect -10228 1500 -4686 1670
rect 280 -1269 15750 -963
<< nsubdiffcont >>
rect -1317 7851 15785 8157
rect -23548 4635 -18142 4805
rect -16718 4647 -11312 4817
rect -10252 4645 -4846 4815
rect 16848 5309 22254 5479
rect 23336 5307 28742 5477
<< poly >>
rect 272 6807 338 6823
rect 272 6773 288 6807
rect 322 6773 338 6807
rect 272 6757 338 6773
rect 2712 6803 2778 6819
rect 2712 6769 2728 6803
rect 2762 6769 2778 6803
rect 290 6702 320 6757
rect 2712 6753 2778 6769
rect 3228 6791 3294 6807
rect 3228 6757 3244 6791
rect 3278 6757 3294 6791
rect 2730 6706 2760 6753
rect 3228 6741 3294 6757
rect 5668 6787 5734 6803
rect 5668 6753 5684 6787
rect 5718 6753 5734 6787
rect 290 6674 370 6702
rect 2682 6696 2760 6706
rect 244 6644 1330 6674
rect 244 6606 274 6644
rect 340 6606 370 6644
rect 436 6606 466 6644
rect 532 6606 562 6644
rect 628 6606 658 6644
rect 724 6606 754 6644
rect 820 6606 850 6644
rect 916 6606 946 6644
rect 1012 6606 1042 6644
rect 1108 6606 1138 6644
rect 1204 6606 1234 6644
rect 1300 6606 1330 6644
rect 2010 6666 2760 6696
rect 3246 6686 3276 6741
rect 5668 6737 5734 6753
rect 6258 6791 6324 6807
rect 6258 6757 6274 6791
rect 6308 6757 6324 6791
rect 6258 6741 6324 6757
rect 8698 6787 8764 6803
rect 8698 6753 8714 6787
rect 8748 6753 8764 6787
rect 5686 6690 5716 6737
rect -1606 5936 -1566 5962
rect -1508 5936 -1468 5962
rect -1410 5936 -1370 5962
rect -1312 5936 -1272 5962
rect -1214 5936 -1174 5962
rect -1116 5936 -1076 5962
rect -1018 5936 -978 5962
rect -920 5936 -880 5962
rect 2010 6602 2040 6666
rect 2106 6602 2136 6666
rect 2202 6602 2232 6666
rect 2298 6602 2328 6666
rect 2394 6602 2424 6666
rect 2490 6602 2520 6666
rect 2586 6602 2616 6666
rect 2682 6602 2712 6666
rect 3246 6658 3326 6686
rect 5638 6680 5716 6690
rect 3200 6628 4286 6658
rect 244 5580 274 5606
rect 340 5580 370 5606
rect 436 5580 466 5606
rect 532 5580 562 5606
rect 628 5580 658 5606
rect 724 5580 754 5606
rect 820 5580 850 5606
rect 916 5580 946 5606
rect 1012 5580 1042 5606
rect 1108 5580 1138 5606
rect 1204 5580 1234 5606
rect 1300 5580 1330 5606
rect 3200 6590 3230 6628
rect 3296 6590 3326 6628
rect 3392 6590 3422 6628
rect 3488 6590 3518 6628
rect 3584 6590 3614 6628
rect 3680 6590 3710 6628
rect 3776 6590 3806 6628
rect 3872 6590 3902 6628
rect 3968 6590 3998 6628
rect 4064 6590 4094 6628
rect 4160 6590 4190 6628
rect 4256 6590 4286 6628
rect 4966 6650 5716 6680
rect 6276 6686 6306 6741
rect 8698 6737 8764 6753
rect 9346 6789 9412 6805
rect 9346 6755 9362 6789
rect 9396 6755 9412 6789
rect 9346 6739 9412 6755
rect 11786 6785 11852 6801
rect 11786 6751 11802 6785
rect 11836 6751 11852 6785
rect 8716 6690 8746 6737
rect 6276 6658 6356 6686
rect 8668 6680 8746 6690
rect 2010 5576 2040 5602
rect 2106 5576 2136 5602
rect 2202 5576 2232 5602
rect 2298 5576 2328 5602
rect 2394 5576 2424 5602
rect 2490 5576 2520 5602
rect 2586 5576 2616 5602
rect 2682 5576 2712 5602
rect 4966 6586 4996 6650
rect 5062 6586 5092 6650
rect 5158 6586 5188 6650
rect 5254 6586 5284 6650
rect 5350 6586 5380 6650
rect 5446 6586 5476 6650
rect 5542 6586 5572 6650
rect 5638 6586 5668 6650
rect 6230 6628 7316 6658
rect 6230 6590 6260 6628
rect 6326 6590 6356 6628
rect 6422 6590 6452 6628
rect 6518 6590 6548 6628
rect 6614 6590 6644 6628
rect 6710 6590 6740 6628
rect 6806 6590 6836 6628
rect 6902 6590 6932 6628
rect 6998 6590 7028 6628
rect 7094 6590 7124 6628
rect 7190 6590 7220 6628
rect 7286 6590 7316 6628
rect 7996 6650 8746 6680
rect 9364 6684 9394 6739
rect 11786 6735 11852 6751
rect 12502 6763 12568 6779
rect 11804 6688 11834 6735
rect 12502 6729 12518 6763
rect 12552 6729 12568 6763
rect 12502 6713 12568 6729
rect 14942 6759 15008 6775
rect 14942 6725 14958 6759
rect 14992 6725 15008 6759
rect 9364 6656 9444 6684
rect 11756 6678 11834 6688
rect 3200 5564 3230 5590
rect 3296 5564 3326 5590
rect 3392 5564 3422 5590
rect 3488 5564 3518 5590
rect 3584 5564 3614 5590
rect 3680 5564 3710 5590
rect 3776 5564 3806 5590
rect 3872 5564 3902 5590
rect 3968 5564 3998 5590
rect 4064 5564 4094 5590
rect 4160 5564 4190 5590
rect 4256 5564 4286 5590
rect 7996 6586 8026 6650
rect 8092 6586 8122 6650
rect 8188 6586 8218 6650
rect 8284 6586 8314 6650
rect 8380 6586 8410 6650
rect 8476 6586 8506 6650
rect 8572 6586 8602 6650
rect 8668 6586 8698 6650
rect 9318 6626 10404 6656
rect 9318 6588 9348 6626
rect 9414 6588 9444 6626
rect 9510 6588 9540 6626
rect 9606 6588 9636 6626
rect 9702 6588 9732 6626
rect 9798 6588 9828 6626
rect 9894 6588 9924 6626
rect 9990 6588 10020 6626
rect 10086 6588 10116 6626
rect 10182 6588 10212 6626
rect 10278 6588 10308 6626
rect 10374 6588 10404 6626
rect 11084 6648 11834 6678
rect 12520 6658 12550 6713
rect 14942 6709 15008 6725
rect 14960 6662 14990 6709
rect 4966 5560 4996 5586
rect 5062 5560 5092 5586
rect 5158 5560 5188 5586
rect 5254 5560 5284 5586
rect 5350 5560 5380 5586
rect 5446 5560 5476 5586
rect 5542 5560 5572 5586
rect 5638 5560 5668 5586
rect 6230 5564 6260 5590
rect 6326 5564 6356 5590
rect 6422 5564 6452 5590
rect 6518 5564 6548 5590
rect 6614 5564 6644 5590
rect 6710 5564 6740 5590
rect 6806 5564 6836 5590
rect 6902 5564 6932 5590
rect 6998 5564 7028 5590
rect 7094 5564 7124 5590
rect 7190 5564 7220 5590
rect 7286 5564 7316 5590
rect 11084 6584 11114 6648
rect 11180 6584 11210 6648
rect 11276 6584 11306 6648
rect 11372 6584 11402 6648
rect 11468 6584 11498 6648
rect 11564 6584 11594 6648
rect 11660 6584 11690 6648
rect 11756 6584 11786 6648
rect 12520 6630 12600 6658
rect 14912 6652 14990 6662
rect 12474 6600 13560 6630
rect 7996 5560 8026 5586
rect 8092 5560 8122 5586
rect 8188 5560 8218 5586
rect 8284 5560 8314 5586
rect 8380 5560 8410 5586
rect 8476 5560 8506 5586
rect 8572 5560 8602 5586
rect 8668 5560 8698 5586
rect 9318 5562 9348 5588
rect 9414 5562 9444 5588
rect 9510 5562 9540 5588
rect 9606 5562 9636 5588
rect 9702 5562 9732 5588
rect 9798 5562 9828 5588
rect 9894 5562 9924 5588
rect 9990 5562 10020 5588
rect 10086 5562 10116 5588
rect 10182 5562 10212 5588
rect 10278 5562 10308 5588
rect 10374 5562 10404 5588
rect 12474 6562 12504 6600
rect 12570 6562 12600 6600
rect 12666 6562 12696 6600
rect 12762 6562 12792 6600
rect 12858 6562 12888 6600
rect 12954 6562 12984 6600
rect 13050 6562 13080 6600
rect 13146 6562 13176 6600
rect 13242 6562 13272 6600
rect 13338 6562 13368 6600
rect 13434 6562 13464 6600
rect 13530 6562 13560 6600
rect 14240 6622 14990 6652
rect 11084 5558 11114 5584
rect 11180 5558 11210 5584
rect 11276 5558 11306 5584
rect 11372 5558 11402 5584
rect 11468 5558 11498 5584
rect 11564 5558 11594 5584
rect 11660 5558 11690 5584
rect 11756 5558 11786 5584
rect 14240 6558 14270 6622
rect 14336 6558 14366 6622
rect 14432 6558 14462 6622
rect 14528 6558 14558 6622
rect 14624 6558 14654 6622
rect 14720 6558 14750 6622
rect 14816 6558 14846 6622
rect 14912 6558 14942 6622
rect 12474 5536 12504 5562
rect 12570 5536 12600 5562
rect 12666 5536 12696 5562
rect 12762 5536 12792 5562
rect 12858 5536 12888 5562
rect 12954 5536 12984 5562
rect 13050 5536 13080 5562
rect 13146 5536 13176 5562
rect 13242 5536 13272 5562
rect 13338 5536 13368 5562
rect 13434 5536 13464 5562
rect 13530 5536 13560 5562
rect 15568 5926 15598 5952
rect 15664 5926 15694 5952
rect 14240 5532 14270 5558
rect 14336 5532 14366 5558
rect 14432 5532 14462 5558
rect 14528 5532 14558 5558
rect 14624 5532 14654 5558
rect 14720 5532 14750 5558
rect 14816 5532 14846 5558
rect 14912 5532 14942 5558
rect 1534 4990 1852 5020
rect 1534 4944 1564 4990
rect 1630 4944 1660 4990
rect 1726 4944 1756 4990
rect 1822 4944 1852 4990
rect 4490 4974 4808 5004
rect -1606 4866 -1566 4936
rect -1508 4866 -1468 4936
rect -1410 4868 -1370 4936
rect -1412 4866 -1370 4868
rect -1312 4866 -1272 4936
rect -1214 4866 -1174 4936
rect -1116 4866 -1076 4936
rect -1018 4866 -978 4936
rect -920 4866 -880 4936
rect -1606 4828 -880 4866
rect -1070 4785 -1030 4828
rect -1083 4769 -1017 4785
rect -1083 4735 -1067 4769
rect -1033 4735 -1017 4769
rect -1083 4719 -1017 4735
rect -23536 4442 -23506 4472
rect -23440 4442 -23410 4468
rect -23344 4442 -23314 4472
rect -23248 4442 -23218 4468
rect -23152 4442 -23122 4472
rect -23056 4442 -23026 4468
rect -22960 4442 -22930 4472
rect -22864 4442 -22834 4468
rect -22768 4442 -22738 4472
rect -22672 4442 -22642 4468
rect -22576 4442 -22546 4472
rect -22480 4442 -22450 4468
rect -22384 4442 -22354 4472
rect -22288 4442 -22258 4468
rect -22192 4442 -22162 4472
rect -22096 4442 -22066 4468
rect -22000 4442 -21970 4472
rect -21904 4442 -21874 4468
rect -21808 4442 -21778 4472
rect -21712 4442 -21682 4468
rect -21392 4448 -21362 4474
rect -21296 4448 -21266 4476
rect -21200 4448 -21170 4474
rect -21104 4448 -21074 4476
rect -21008 4448 -20978 4474
rect -20912 4448 -20882 4476
rect -20816 4448 -20786 4474
rect -20720 4448 -20690 4476
rect -20624 4448 -20594 4474
rect -20528 4448 -20498 4476
rect -20432 4448 -20402 4474
rect -20336 4448 -20306 4476
rect -20240 4448 -20210 4474
rect -20144 4448 -20114 4476
rect -20048 4448 -20018 4474
rect -19708 4454 -19678 4480
rect -19612 4454 -19582 4480
rect -19516 4454 -19486 4480
rect -19420 4454 -19390 4480
rect -19324 4454 -19294 4480
rect -19228 4454 -19198 4480
rect -19132 4454 -19102 4480
rect -19036 4454 -19006 4480
rect -18940 4454 -18910 4480
rect -18844 4454 -18814 4480
rect -18540 4456 -18510 4482
rect -18444 4456 -18414 4484
rect -18348 4456 -18318 4482
rect -18252 4456 -18222 4484
rect -18156 4456 -18126 4482
rect -16706 4454 -16676 4484
rect -16610 4454 -16580 4480
rect -16514 4454 -16484 4484
rect -16418 4454 -16388 4480
rect -16322 4454 -16292 4484
rect -16226 4454 -16196 4480
rect -16130 4454 -16100 4484
rect -16034 4454 -16004 4480
rect -15938 4454 -15908 4484
rect -15842 4454 -15812 4480
rect -15746 4454 -15716 4484
rect -15650 4454 -15620 4480
rect -15554 4454 -15524 4484
rect -15458 4454 -15428 4480
rect -15362 4454 -15332 4484
rect -15266 4454 -15236 4480
rect -15170 4454 -15140 4484
rect -15074 4454 -15044 4480
rect -14978 4454 -14948 4484
rect -14882 4454 -14852 4480
rect -14562 4460 -14532 4486
rect -14466 4460 -14436 4488
rect -14370 4460 -14340 4486
rect -14274 4460 -14244 4488
rect -14178 4460 -14148 4486
rect -14082 4460 -14052 4488
rect -13986 4460 -13956 4486
rect -13890 4460 -13860 4488
rect -13794 4460 -13764 4486
rect -13698 4460 -13668 4488
rect -13602 4460 -13572 4486
rect -13506 4460 -13476 4488
rect -13410 4460 -13380 4486
rect -13314 4460 -13284 4488
rect -13218 4460 -13188 4486
rect -12878 4466 -12848 4492
rect -12782 4466 -12752 4492
rect -12686 4466 -12656 4492
rect -12590 4466 -12560 4492
rect -12494 4466 -12464 4492
rect -12398 4466 -12368 4492
rect -12302 4466 -12272 4492
rect -12206 4466 -12176 4492
rect -12110 4466 -12080 4492
rect -12014 4466 -11984 4492
rect -11710 4468 -11680 4494
rect -11614 4468 -11584 4496
rect -11518 4468 -11488 4494
rect -11422 4468 -11392 4496
rect -11326 4468 -11296 4494
rect -23536 3418 -23506 3442
rect -23440 3418 -23410 3442
rect -23344 3418 -23314 3442
rect -23248 3418 -23218 3442
rect -23152 3418 -23122 3442
rect -23056 3418 -23026 3442
rect -22960 3418 -22930 3442
rect -22864 3418 -22834 3442
rect -22768 3418 -22738 3442
rect -22672 3418 -22642 3442
rect -22576 3418 -22546 3442
rect -22480 3418 -22450 3442
rect -22384 3418 -22354 3442
rect -22288 3418 -22258 3442
rect -22192 3418 -22162 3442
rect -22096 3418 -22066 3442
rect -22000 3418 -21970 3442
rect -21904 3418 -21874 3442
rect -21808 3418 -21778 3442
rect -21712 3418 -21682 3442
rect -23536 3388 -21682 3418
rect -21392 3430 -21362 3448
rect -21296 3430 -21266 3448
rect -21200 3430 -21170 3448
rect -21104 3430 -21074 3448
rect -21008 3430 -20978 3448
rect -20912 3430 -20882 3448
rect -20816 3430 -20786 3448
rect -20720 3430 -20690 3448
rect -20624 3430 -20594 3448
rect -20528 3430 -20498 3448
rect -20432 3430 -20402 3448
rect -20336 3430 -20306 3448
rect -20240 3430 -20210 3448
rect -20144 3430 -20114 3448
rect -20048 3430 -20018 3448
rect -21392 3400 -20018 3430
rect -19708 3430 -19678 3454
rect -19612 3430 -19582 3454
rect -19516 3430 -19486 3454
rect -19420 3430 -19390 3454
rect -19324 3430 -19294 3454
rect -19228 3430 -19198 3454
rect -19132 3430 -19102 3454
rect -19036 3430 -19006 3454
rect -18940 3430 -18910 3454
rect -18844 3430 -18814 3454
rect -19708 3400 -18814 3430
rect -18540 3440 -18510 3456
rect -18444 3440 -18414 3456
rect -18348 3440 -18318 3456
rect -18252 3440 -18222 3456
rect -18156 3440 -18126 3456
rect -10240 4452 -10210 4482
rect -10144 4452 -10114 4478
rect -10048 4452 -10018 4482
rect -9952 4452 -9922 4478
rect -9856 4452 -9826 4482
rect -9760 4452 -9730 4478
rect -9664 4452 -9634 4482
rect -9568 4452 -9538 4478
rect -9472 4452 -9442 4482
rect -9376 4452 -9346 4478
rect -9280 4452 -9250 4482
rect -9184 4452 -9154 4478
rect -9088 4452 -9058 4482
rect -8992 4452 -8962 4478
rect -8896 4452 -8866 4482
rect -8800 4452 -8770 4478
rect -8704 4452 -8674 4482
rect -8608 4452 -8578 4478
rect -8512 4452 -8482 4482
rect -8416 4452 -8386 4478
rect -8096 4458 -8066 4484
rect -8000 4458 -7970 4486
rect -7904 4458 -7874 4484
rect -7808 4458 -7778 4486
rect -7712 4458 -7682 4484
rect -7616 4458 -7586 4486
rect -7520 4458 -7490 4484
rect -7424 4458 -7394 4486
rect -7328 4458 -7298 4484
rect -7232 4458 -7202 4486
rect -7136 4458 -7106 4484
rect -7040 4458 -7010 4486
rect -6944 4458 -6914 4484
rect -6848 4458 -6818 4486
rect -6752 4458 -6722 4484
rect -6412 4464 -6382 4490
rect -6316 4464 -6286 4490
rect -6220 4464 -6190 4490
rect -6124 4464 -6094 4490
rect -6028 4464 -5998 4490
rect -5932 4464 -5902 4490
rect -5836 4464 -5806 4490
rect -5740 4464 -5710 4490
rect -5644 4464 -5614 4490
rect -5548 4464 -5518 4490
rect -5244 4466 -5214 4492
rect -5148 4466 -5118 4494
rect -5052 4466 -5022 4492
rect -4956 4466 -4926 4494
rect -4860 4466 -4830 4492
rect -18540 3410 -18126 3440
rect -21712 3291 -21682 3388
rect -20048 3297 -20018 3400
rect -18844 3303 -18814 3400
rect -21730 3275 -21664 3291
rect -21730 3241 -21714 3275
rect -21680 3241 -21664 3275
rect -21730 3225 -21664 3241
rect -20066 3281 -20000 3297
rect -20066 3247 -20050 3281
rect -20016 3247 -20000 3281
rect -20066 3231 -20000 3247
rect -18862 3287 -18796 3303
rect -18862 3253 -18846 3287
rect -18812 3253 -18796 3287
rect -18156 3285 -18126 3410
rect -16706 3434 -16676 3454
rect -16610 3434 -16580 3454
rect -16514 3434 -16484 3454
rect -16418 3434 -16388 3454
rect -16322 3434 -16292 3454
rect -16226 3434 -16196 3454
rect -16130 3434 -16100 3454
rect -16034 3434 -16004 3454
rect -15938 3434 -15908 3454
rect -15842 3434 -15812 3454
rect -15746 3434 -15716 3454
rect -15650 3434 -15620 3454
rect -15554 3434 -15524 3454
rect -15458 3434 -15428 3454
rect -15362 3434 -15332 3454
rect -15266 3434 -15236 3454
rect -15170 3434 -15140 3454
rect -15074 3434 -15044 3454
rect -14978 3434 -14948 3454
rect -14882 3434 -14852 3454
rect -16706 3404 -14852 3434
rect -14562 3442 -14532 3460
rect -14466 3442 -14436 3460
rect -14370 3442 -14340 3460
rect -14274 3442 -14244 3460
rect -14178 3442 -14148 3460
rect -14082 3442 -14052 3460
rect -13986 3442 -13956 3460
rect -13890 3442 -13860 3460
rect -13794 3442 -13764 3460
rect -13698 3442 -13668 3460
rect -13602 3442 -13572 3460
rect -13506 3442 -13476 3460
rect -13410 3442 -13380 3460
rect -13314 3442 -13284 3460
rect -13218 3442 -13188 3460
rect -14562 3412 -13188 3442
rect -12878 3442 -12848 3466
rect -12782 3442 -12752 3466
rect -12686 3442 -12656 3466
rect -12590 3442 -12560 3466
rect -12494 3442 -12464 3466
rect -12398 3442 -12368 3466
rect -12302 3442 -12272 3466
rect -12206 3442 -12176 3466
rect -12110 3442 -12080 3466
rect -12014 3442 -11984 3466
rect -12878 3412 -11984 3442
rect -11710 3452 -11680 3468
rect -11614 3452 -11584 3468
rect -11518 3452 -11488 3468
rect -11422 3452 -11392 3468
rect -11326 3452 -11296 3468
rect 4490 4928 4520 4974
rect 4586 4928 4616 4974
rect 4682 4928 4712 4974
rect 4778 4928 4808 4974
rect 7520 4974 7838 5004
rect 7520 4928 7550 4974
rect 7616 4928 7646 4974
rect 7712 4928 7742 4974
rect 7808 4928 7838 4974
rect 10608 4972 10926 5002
rect 1534 3874 1564 3944
rect 1630 3918 1660 3944
rect 1726 3874 1756 3944
rect 1822 3918 1852 3944
rect 10608 4926 10638 4972
rect 10704 4926 10734 4972
rect 10800 4926 10830 4972
rect 10896 4926 10926 4972
rect 13764 4946 14082 4976
rect 1534 3844 1612 3874
rect 1726 3844 1804 3874
rect 1582 3793 1612 3844
rect 1774 3793 1804 3844
rect 4490 3858 4520 3928
rect 4586 3902 4616 3928
rect 4682 3858 4712 3928
rect 4778 3902 4808 3928
rect 7520 3858 7550 3928
rect 7616 3902 7646 3928
rect 7712 3858 7742 3928
rect 7808 3902 7838 3928
rect 13764 4900 13794 4946
rect 13860 4900 13890 4946
rect 13956 4900 13986 4946
rect 14052 4900 14082 4946
rect 4490 3828 4568 3858
rect 4682 3828 4760 3858
rect 7520 3828 7598 3858
rect 7712 3828 7790 3858
rect 1564 3777 1630 3793
rect 1564 3743 1580 3777
rect 1614 3743 1630 3777
rect 1564 3727 1630 3743
rect 1756 3777 1822 3793
rect 4538 3777 4568 3828
rect 4730 3777 4760 3828
rect 7568 3777 7598 3828
rect 7760 3777 7790 3828
rect 10608 3856 10638 3926
rect 10704 3900 10734 3926
rect 10800 3856 10830 3926
rect 10896 3900 10926 3926
rect 16832 5130 16862 5156
rect 16928 5130 16958 5158
rect 17024 5130 17054 5156
rect 17120 5130 17150 5158
rect 17216 5130 17246 5156
rect 17520 5128 17550 5154
rect 17616 5128 17646 5154
rect 17712 5128 17742 5154
rect 17808 5128 17838 5154
rect 17904 5128 17934 5154
rect 18000 5128 18030 5154
rect 18096 5128 18126 5154
rect 18192 5128 18222 5154
rect 18288 5128 18318 5154
rect 18384 5128 18414 5154
rect 16832 4114 16862 4130
rect 16928 4114 16958 4130
rect 17024 4114 17054 4130
rect 17120 4114 17150 4130
rect 17216 4114 17246 4130
rect 18724 5122 18754 5148
rect 18820 5122 18850 5150
rect 18916 5122 18946 5148
rect 19012 5122 19042 5150
rect 19108 5122 19138 5148
rect 19204 5122 19234 5150
rect 19300 5122 19330 5148
rect 19396 5122 19426 5150
rect 19492 5122 19522 5148
rect 19588 5122 19618 5150
rect 19684 5122 19714 5148
rect 19780 5122 19810 5150
rect 19876 5122 19906 5148
rect 19972 5122 20002 5150
rect 20068 5122 20098 5148
rect 16832 4084 17246 4114
rect 17520 4104 17550 4128
rect 17616 4104 17646 4128
rect 17712 4104 17742 4128
rect 17808 4104 17838 4128
rect 17904 4104 17934 4128
rect 18000 4104 18030 4128
rect 18096 4104 18126 4128
rect 18192 4104 18222 4128
rect 18288 4104 18318 4128
rect 18384 4104 18414 4128
rect 20388 5116 20418 5142
rect 20484 5116 20514 5146
rect 20580 5116 20610 5142
rect 20676 5116 20706 5146
rect 20772 5116 20802 5142
rect 20868 5116 20898 5146
rect 20964 5116 20994 5142
rect 21060 5116 21090 5146
rect 21156 5116 21186 5142
rect 21252 5116 21282 5146
rect 21348 5116 21378 5142
rect 21444 5116 21474 5146
rect 21540 5116 21570 5142
rect 21636 5116 21666 5146
rect 21732 5116 21762 5142
rect 21828 5116 21858 5146
rect 21924 5116 21954 5142
rect 22020 5116 22050 5146
rect 22116 5116 22146 5142
rect 22212 5116 22242 5146
rect 23320 5128 23350 5154
rect 23416 5128 23446 5156
rect 23512 5128 23542 5154
rect 23608 5128 23638 5156
rect 23704 5128 23734 5154
rect 16832 3959 16862 4084
rect 17520 4074 18414 4104
rect 18724 4104 18754 4122
rect 18820 4104 18850 4122
rect 18916 4104 18946 4122
rect 19012 4104 19042 4122
rect 19108 4104 19138 4122
rect 19204 4104 19234 4122
rect 19300 4104 19330 4122
rect 19396 4104 19426 4122
rect 19492 4104 19522 4122
rect 19588 4104 19618 4122
rect 19684 4104 19714 4122
rect 19780 4104 19810 4122
rect 19876 4104 19906 4122
rect 19972 4104 20002 4122
rect 20068 4104 20098 4122
rect 24008 5126 24038 5152
rect 24104 5126 24134 5152
rect 24200 5126 24230 5152
rect 24296 5126 24326 5152
rect 24392 5126 24422 5152
rect 24488 5126 24518 5152
rect 24584 5126 24614 5152
rect 24680 5126 24710 5152
rect 24776 5126 24806 5152
rect 24872 5126 24902 5152
rect 18724 4074 20098 4104
rect 20388 4094 20418 4116
rect 20484 4094 20514 4116
rect 20580 4094 20610 4116
rect 20676 4094 20706 4116
rect 20772 4094 20802 4116
rect 20868 4094 20898 4116
rect 20964 4094 20994 4116
rect 21060 4094 21090 4116
rect 21156 4094 21186 4116
rect 21252 4094 21282 4116
rect 21348 4094 21378 4116
rect 21444 4094 21474 4116
rect 21540 4094 21570 4116
rect 21636 4094 21666 4116
rect 21732 4094 21762 4116
rect 21828 4094 21858 4116
rect 21924 4094 21954 4116
rect 22020 4094 22050 4116
rect 22116 4094 22146 4116
rect 22212 4094 22242 4116
rect 17520 3977 17550 4074
rect 17502 3961 17568 3977
rect 18724 3971 18754 4074
rect 20388 4064 22242 4094
rect 23320 4112 23350 4128
rect 23416 4112 23446 4128
rect 23512 4112 23542 4128
rect 23608 4112 23638 4128
rect 23704 4112 23734 4128
rect 25212 5120 25242 5146
rect 25308 5120 25338 5148
rect 25404 5120 25434 5146
rect 25500 5120 25530 5148
rect 25596 5120 25626 5146
rect 25692 5120 25722 5148
rect 25788 5120 25818 5146
rect 25884 5120 25914 5148
rect 25980 5120 26010 5146
rect 26076 5120 26106 5148
rect 26172 5120 26202 5146
rect 26268 5120 26298 5148
rect 26364 5120 26394 5146
rect 26460 5120 26490 5148
rect 26556 5120 26586 5146
rect 23320 4082 23734 4112
rect 24008 4102 24038 4126
rect 24104 4102 24134 4126
rect 24200 4102 24230 4126
rect 24296 4102 24326 4126
rect 24392 4102 24422 4126
rect 24488 4102 24518 4126
rect 24584 4102 24614 4126
rect 24680 4102 24710 4126
rect 24776 4102 24806 4126
rect 24872 4102 24902 4126
rect 26876 5114 26906 5140
rect 26972 5114 27002 5144
rect 27068 5114 27098 5140
rect 27164 5114 27194 5144
rect 27260 5114 27290 5140
rect 27356 5114 27386 5144
rect 27452 5114 27482 5140
rect 27548 5114 27578 5144
rect 27644 5114 27674 5140
rect 27740 5114 27770 5144
rect 27836 5114 27866 5140
rect 27932 5114 27962 5144
rect 28028 5114 28058 5140
rect 28124 5114 28154 5144
rect 28220 5114 28250 5140
rect 28316 5114 28346 5144
rect 28412 5114 28442 5140
rect 28508 5114 28538 5144
rect 28604 5114 28634 5140
rect 28700 5114 28730 5144
rect 16814 3943 16880 3959
rect 10608 3826 10686 3856
rect 10800 3826 10878 3856
rect 1756 3743 1772 3777
rect 1806 3743 1822 3777
rect 1756 3727 1822 3743
rect 4520 3761 4586 3777
rect 4520 3727 4536 3761
rect 4570 3727 4586 3761
rect 4520 3711 4586 3727
rect 4712 3761 4778 3777
rect 4712 3727 4728 3761
rect 4762 3727 4778 3761
rect 4712 3711 4778 3727
rect 7550 3761 7616 3777
rect 7550 3727 7566 3761
rect 7600 3727 7616 3761
rect 7550 3711 7616 3727
rect 7742 3761 7808 3777
rect 10656 3775 10686 3826
rect 10848 3775 10878 3826
rect 13764 3830 13794 3900
rect 13860 3874 13890 3900
rect 13956 3830 13986 3900
rect 14052 3874 14082 3900
rect 15568 3876 15598 3926
rect 15664 3876 15694 3926
rect 16814 3909 16830 3943
rect 16864 3909 16880 3943
rect 17502 3927 17518 3961
rect 17552 3927 17568 3961
rect 17502 3911 17568 3927
rect 18706 3955 18772 3971
rect 20388 3965 20418 4064
rect 18706 3921 18722 3955
rect 18756 3921 18772 3955
rect 16814 3893 16880 3909
rect 18706 3905 18772 3921
rect 20370 3949 20436 3965
rect 23320 3957 23350 4082
rect 24008 4072 24902 4102
rect 25212 4102 25242 4120
rect 25308 4102 25338 4120
rect 25404 4102 25434 4120
rect 25500 4102 25530 4120
rect 25596 4102 25626 4120
rect 25692 4102 25722 4120
rect 25788 4102 25818 4120
rect 25884 4102 25914 4120
rect 25980 4102 26010 4120
rect 26076 4102 26106 4120
rect 26172 4102 26202 4120
rect 26268 4102 26298 4120
rect 26364 4102 26394 4120
rect 26460 4102 26490 4120
rect 26556 4102 26586 4120
rect 25212 4072 26586 4102
rect 26876 4096 26906 4114
rect 26972 4096 27002 4114
rect 27068 4096 27098 4114
rect 27164 4096 27194 4114
rect 27260 4096 27290 4114
rect 27356 4096 27386 4114
rect 27452 4096 27482 4114
rect 27548 4096 27578 4114
rect 27644 4096 27674 4114
rect 27740 4096 27770 4114
rect 27836 4096 27866 4114
rect 27932 4096 27962 4114
rect 28028 4096 28058 4114
rect 28124 4096 28154 4114
rect 28220 4096 28250 4114
rect 28316 4096 28346 4114
rect 28412 4096 28442 4114
rect 28508 4096 28538 4114
rect 28604 4096 28634 4114
rect 28700 4096 28730 4114
rect 24008 3975 24038 4072
rect 23990 3959 24056 3975
rect 25212 3969 25242 4072
rect 26876 4066 28736 4096
rect 20370 3915 20386 3949
rect 20420 3915 20436 3949
rect 20370 3899 20436 3915
rect 23302 3941 23368 3957
rect 23302 3907 23318 3941
rect 23352 3907 23368 3941
rect 23990 3925 24006 3959
rect 24040 3925 24056 3959
rect 23990 3909 24056 3925
rect 25194 3953 25260 3969
rect 26876 3963 26906 4066
rect 25194 3919 25210 3953
rect 25244 3919 25260 3953
rect 23302 3891 23368 3907
rect 25194 3903 25260 3919
rect 26858 3947 26924 3963
rect 26858 3913 26874 3947
rect 26908 3913 26924 3947
rect 26858 3897 26924 3913
rect 15568 3846 15694 3876
rect 13764 3800 13842 3830
rect 13956 3800 14034 3830
rect 7742 3727 7758 3761
rect 7792 3727 7808 3761
rect 7742 3711 7808 3727
rect 10638 3759 10704 3775
rect 10638 3725 10654 3759
rect 10688 3725 10704 3759
rect 10638 3709 10704 3725
rect 10830 3759 10896 3775
rect 10830 3725 10846 3759
rect 10880 3725 10896 3759
rect 13812 3749 13842 3800
rect 14004 3749 14034 3800
rect 15568 3795 15598 3846
rect 15550 3779 15616 3795
rect 10830 3709 10896 3725
rect 13794 3733 13860 3749
rect 13794 3699 13810 3733
rect 13844 3699 13860 3733
rect 13794 3683 13860 3699
rect 13986 3733 14052 3749
rect 13986 3699 14002 3733
rect 14036 3699 14052 3733
rect 15550 3745 15566 3779
rect 15600 3745 15616 3779
rect 15550 3729 15616 3745
rect 17506 3736 17572 3752
rect 13986 3683 14052 3699
rect 16814 3706 16880 3722
rect 16814 3672 16830 3706
rect 16864 3672 16880 3706
rect 17506 3702 17522 3736
rect 17556 3702 17572 3736
rect 23994 3734 24060 3750
rect 17506 3686 17572 3702
rect 18704 3692 18770 3708
rect 16814 3656 16880 3672
rect 16832 3586 16862 3656
rect 16736 3556 17150 3586
rect 17524 3570 17554 3686
rect 18704 3658 18720 3692
rect 18754 3658 18770 3692
rect 18704 3642 18770 3658
rect 20372 3690 20438 3706
rect 20372 3656 20388 3690
rect 20422 3656 20438 3690
rect 18722 3570 18752 3642
rect 20372 3640 20438 3656
rect 23302 3704 23368 3720
rect 23302 3670 23318 3704
rect 23352 3670 23368 3704
rect 23994 3700 24010 3734
rect 24044 3700 24060 3734
rect 23994 3684 24060 3700
rect 25192 3690 25258 3706
rect 23302 3654 23368 3670
rect 20390 3578 20420 3640
rect 23320 3584 23350 3654
rect 16736 3534 16766 3556
rect 16832 3534 16862 3556
rect 16928 3534 16958 3556
rect 17024 3534 17054 3556
rect 17120 3534 17150 3556
rect 17428 3540 18322 3570
rect -11710 3422 -11296 3452
rect -14882 3303 -14852 3404
rect -13218 3309 -13188 3412
rect -12014 3315 -11984 3412
rect -14900 3287 -14834 3303
rect -18862 3237 -18796 3253
rect -18174 3269 -18108 3285
rect -18174 3235 -18158 3269
rect -18124 3235 -18108 3269
rect -14900 3253 -14884 3287
rect -14850 3253 -14834 3287
rect -14900 3237 -14834 3253
rect -13236 3293 -13170 3309
rect -13236 3259 -13220 3293
rect -13186 3259 -13170 3293
rect -13236 3243 -13170 3259
rect -12032 3299 -11966 3315
rect -12032 3265 -12016 3299
rect -11982 3265 -11966 3299
rect -11326 3297 -11296 3422
rect -10240 3430 -10210 3452
rect -10144 3430 -10114 3452
rect -10048 3430 -10018 3452
rect -9952 3430 -9922 3452
rect -9856 3430 -9826 3452
rect -9760 3430 -9730 3452
rect -9664 3430 -9634 3452
rect -9568 3430 -9538 3452
rect -9472 3430 -9442 3452
rect -9376 3430 -9346 3452
rect -9280 3430 -9250 3452
rect -9184 3430 -9154 3452
rect -9088 3430 -9058 3452
rect -8992 3430 -8962 3452
rect -8896 3430 -8866 3452
rect -8800 3430 -8770 3452
rect -8704 3430 -8674 3452
rect -8608 3430 -8578 3452
rect -8512 3430 -8482 3452
rect -8416 3430 -8386 3452
rect -10240 3400 -8386 3430
rect -8096 3440 -8066 3458
rect -8000 3440 -7970 3458
rect -7904 3440 -7874 3458
rect -7808 3440 -7778 3458
rect -7712 3440 -7682 3458
rect -7616 3440 -7586 3458
rect -7520 3440 -7490 3458
rect -7424 3440 -7394 3458
rect -7328 3440 -7298 3458
rect -7232 3440 -7202 3458
rect -7136 3440 -7106 3458
rect -7040 3440 -7010 3458
rect -6944 3440 -6914 3458
rect -6848 3440 -6818 3458
rect -6752 3440 -6722 3458
rect -8096 3410 -6722 3440
rect -6412 3440 -6382 3464
rect -6316 3440 -6286 3464
rect -6220 3440 -6190 3464
rect -6124 3440 -6094 3464
rect -6028 3440 -5998 3464
rect -5932 3440 -5902 3464
rect -5836 3440 -5806 3464
rect -5740 3440 -5710 3464
rect -5644 3440 -5614 3464
rect -5548 3440 -5518 3464
rect -6412 3410 -5518 3440
rect -5244 3450 -5214 3466
rect -5148 3450 -5118 3466
rect -5052 3450 -5022 3466
rect -4956 3450 -4926 3466
rect -4860 3450 -4830 3466
rect -5244 3420 -4830 3450
rect -8416 3301 -8386 3400
rect -6752 3307 -6722 3410
rect -5548 3313 -5518 3410
rect -12032 3249 -11966 3265
rect -11344 3281 -11278 3297
rect -11344 3247 -11328 3281
rect -11294 3247 -11278 3281
rect -18174 3219 -18108 3235
rect -11344 3231 -11278 3247
rect -8434 3285 -8368 3301
rect -8434 3251 -8418 3285
rect -8384 3251 -8368 3285
rect -8434 3235 -8368 3251
rect -6770 3291 -6704 3307
rect -6770 3257 -6754 3291
rect -6720 3257 -6704 3291
rect -6770 3241 -6704 3257
rect -5566 3297 -5500 3313
rect -5566 3263 -5550 3297
rect -5516 3263 -5500 3297
rect -4860 3295 -4830 3420
rect -1606 3428 -1540 3444
rect -1606 3394 -1590 3428
rect -1556 3394 -1540 3428
rect -1606 3378 -1540 3394
rect -1590 3336 -1560 3378
rect -1636 3300 -934 3336
rect -5566 3247 -5500 3263
rect -4878 3279 -4812 3295
rect -4878 3245 -4862 3279
rect -4828 3245 -4812 3279
rect -4878 3229 -4812 3245
rect -1636 3236 -1606 3300
rect -1540 3236 -1510 3300
rect -1444 3236 -1414 3300
rect -1348 3236 -1318 3300
rect -1252 3236 -1222 3300
rect -1156 3236 -1126 3300
rect -1060 3236 -1030 3300
rect -964 3236 -934 3300
rect -18866 3062 -18800 3078
rect -21732 3016 -21666 3032
rect -21732 2982 -21716 3016
rect -21682 2982 -21666 3016
rect -21732 2966 -21666 2982
rect -20064 3018 -19998 3034
rect -20064 2984 -20048 3018
rect -20014 2984 -19998 3018
rect -18866 3028 -18850 3062
rect -18816 3028 -18800 3062
rect -12036 3074 -11970 3090
rect -18866 3012 -18800 3028
rect -18174 3032 -18108 3048
rect -20064 2968 -19998 2984
rect -21714 2904 -21684 2966
rect -23442 2874 -21588 2904
rect -20046 2896 -20016 2968
rect -18848 2896 -18818 3012
rect -18174 2998 -18158 3032
rect -18124 2998 -18108 3032
rect -18174 2982 -18108 2998
rect -14902 3028 -14836 3044
rect -14902 2994 -14886 3028
rect -14852 2994 -14836 3028
rect -18156 2912 -18126 2982
rect -14902 2978 -14836 2994
rect -13234 3030 -13168 3046
rect -13234 2996 -13218 3030
rect -13184 2996 -13168 3030
rect -12036 3040 -12020 3074
rect -11986 3040 -11970 3074
rect -5570 3072 -5504 3088
rect -12036 3024 -11970 3040
rect -11344 3044 -11278 3060
rect -13234 2980 -13168 2996
rect -14884 2916 -14854 2978
rect -23442 2854 -23412 2874
rect -23346 2854 -23316 2874
rect -23250 2854 -23220 2874
rect -23154 2854 -23124 2874
rect -23058 2854 -23028 2874
rect -22962 2854 -22932 2874
rect -22866 2854 -22836 2874
rect -22770 2854 -22740 2874
rect -22674 2854 -22644 2874
rect -22578 2854 -22548 2874
rect -22482 2854 -22452 2874
rect -22386 2854 -22356 2874
rect -22290 2854 -22260 2874
rect -22194 2854 -22164 2874
rect -22098 2854 -22068 2874
rect -22002 2854 -21972 2874
rect -21906 2854 -21876 2874
rect -21810 2854 -21780 2874
rect -21714 2854 -21684 2874
rect -21618 2854 -21588 2874
rect -21294 2864 -19920 2896
rect -21294 2846 -21264 2864
rect -21198 2846 -21168 2864
rect -21102 2846 -21072 2864
rect -21006 2846 -20976 2864
rect -20910 2846 -20880 2864
rect -20814 2846 -20784 2864
rect -20718 2846 -20688 2864
rect -20622 2846 -20592 2864
rect -20526 2846 -20496 2864
rect -20430 2846 -20400 2864
rect -20334 2846 -20304 2864
rect -20238 2846 -20208 2864
rect -20142 2846 -20112 2864
rect -20046 2846 -20016 2864
rect -19950 2846 -19920 2864
rect -19616 2866 -18722 2896
rect -19616 2850 -19586 2866
rect -19520 2850 -19490 2866
rect -19424 2850 -19394 2866
rect -19328 2850 -19298 2866
rect -19232 2850 -19202 2866
rect -19136 2850 -19106 2866
rect -19040 2850 -19010 2866
rect -18944 2850 -18914 2866
rect -18848 2850 -18818 2866
rect -18752 2850 -18722 2866
rect -18444 2882 -18030 2912
rect -18444 2860 -18414 2882
rect -18348 2860 -18318 2882
rect -18252 2860 -18222 2882
rect -18156 2860 -18126 2882
rect -18060 2860 -18030 2882
rect -16612 2886 -14758 2916
rect -13216 2908 -13186 2980
rect -12018 2908 -11988 3024
rect -11344 3010 -11328 3044
rect -11294 3010 -11278 3044
rect -11344 2994 -11278 3010
rect -8436 3026 -8370 3042
rect -11326 2924 -11296 2994
rect -8436 2992 -8420 3026
rect -8386 2992 -8370 3026
rect -8436 2976 -8370 2992
rect -6768 3028 -6702 3044
rect -6768 2994 -6752 3028
rect -6718 2994 -6702 3028
rect -5570 3038 -5554 3072
rect -5520 3038 -5504 3072
rect -5570 3022 -5504 3038
rect -4878 3042 -4812 3058
rect -6768 2978 -6702 2994
rect -16612 2866 -16582 2886
rect -16516 2866 -16486 2886
rect -16420 2866 -16390 2886
rect -16324 2866 -16294 2886
rect -16228 2866 -16198 2886
rect -16132 2866 -16102 2886
rect -16036 2866 -16006 2886
rect -15940 2866 -15910 2886
rect -15844 2866 -15814 2886
rect -15748 2866 -15718 2886
rect -15652 2866 -15622 2886
rect -15556 2866 -15526 2886
rect -15460 2866 -15430 2886
rect -15364 2866 -15334 2886
rect -15268 2866 -15238 2886
rect -15172 2866 -15142 2886
rect -15076 2866 -15046 2886
rect -14980 2866 -14950 2886
rect -14884 2866 -14854 2886
rect -14788 2866 -14758 2886
rect -14464 2876 -13090 2908
rect -23442 1828 -23412 1854
rect -23346 1828 -23316 1854
rect -23250 1828 -23220 1854
rect -23154 1828 -23124 1854
rect -23058 1828 -23028 1854
rect -22962 1828 -22932 1854
rect -22866 1828 -22836 1854
rect -22770 1828 -22740 1854
rect -22674 1828 -22644 1854
rect -22578 1828 -22548 1854
rect -22482 1828 -22452 1854
rect -22386 1828 -22356 1854
rect -22290 1828 -22260 1854
rect -22194 1828 -22164 1854
rect -22098 1828 -22068 1854
rect -22002 1828 -21972 1854
rect -21906 1828 -21876 1854
rect -21810 1828 -21780 1854
rect -21714 1828 -21684 1854
rect -21618 1828 -21588 1854
rect -14464 2858 -14434 2876
rect -14368 2858 -14338 2876
rect -14272 2858 -14242 2876
rect -14176 2858 -14146 2876
rect -14080 2858 -14050 2876
rect -13984 2858 -13954 2876
rect -13888 2858 -13858 2876
rect -13792 2858 -13762 2876
rect -13696 2858 -13666 2876
rect -13600 2858 -13570 2876
rect -13504 2858 -13474 2876
rect -13408 2858 -13378 2876
rect -13312 2858 -13282 2876
rect -13216 2858 -13186 2876
rect -13120 2858 -13090 2876
rect -12786 2878 -11892 2908
rect -12786 2862 -12756 2878
rect -12690 2862 -12660 2878
rect -12594 2862 -12564 2878
rect -12498 2862 -12468 2878
rect -12402 2862 -12372 2878
rect -12306 2862 -12276 2878
rect -12210 2862 -12180 2878
rect -12114 2862 -12084 2878
rect -12018 2862 -11988 2878
rect -11922 2862 -11892 2878
rect -11614 2894 -11200 2924
rect -8418 2914 -8388 2976
rect -11614 2872 -11584 2894
rect -11518 2872 -11488 2894
rect -11422 2872 -11392 2894
rect -11326 2872 -11296 2894
rect -11230 2872 -11200 2894
rect -10146 2884 -8292 2914
rect -6750 2906 -6720 2978
rect -5552 2906 -5522 3022
rect -4878 3008 -4862 3042
rect -4828 3008 -4812 3042
rect -4878 2992 -4812 3008
rect -4860 2922 -4830 2992
rect -21294 1820 -21264 1846
rect -21198 1820 -21168 1846
rect -21102 1820 -21072 1846
rect -21006 1820 -20976 1846
rect -20910 1820 -20880 1846
rect -20814 1820 -20784 1846
rect -20718 1820 -20688 1846
rect -20622 1820 -20592 1846
rect -20526 1820 -20496 1846
rect -20430 1820 -20400 1846
rect -20334 1820 -20304 1846
rect -20238 1820 -20208 1846
rect -20142 1820 -20112 1846
rect -20046 1820 -20016 1846
rect -19950 1820 -19920 1846
rect -19616 1824 -19586 1850
rect -19520 1824 -19490 1850
rect -19424 1824 -19394 1850
rect -19328 1824 -19298 1850
rect -19232 1824 -19202 1850
rect -19136 1824 -19106 1850
rect -19040 1824 -19010 1850
rect -18944 1824 -18914 1850
rect -18848 1824 -18818 1850
rect -18752 1824 -18722 1850
rect -18444 1834 -18414 1860
rect -18348 1834 -18318 1860
rect -18252 1834 -18222 1860
rect -18156 1834 -18126 1860
rect -18060 1834 -18030 1860
rect -16612 1840 -16582 1866
rect -16516 1840 -16486 1866
rect -16420 1840 -16390 1866
rect -16324 1840 -16294 1866
rect -16228 1840 -16198 1866
rect -16132 1840 -16102 1866
rect -16036 1840 -16006 1866
rect -15940 1840 -15910 1866
rect -15844 1840 -15814 1866
rect -15748 1840 -15718 1866
rect -15652 1840 -15622 1866
rect -15556 1840 -15526 1866
rect -15460 1840 -15430 1866
rect -15364 1840 -15334 1866
rect -15268 1840 -15238 1866
rect -15172 1840 -15142 1866
rect -15076 1840 -15046 1866
rect -14980 1840 -14950 1866
rect -14884 1840 -14854 1866
rect -14788 1840 -14758 1866
rect -10146 2864 -10116 2884
rect -10050 2864 -10020 2884
rect -9954 2864 -9924 2884
rect -9858 2864 -9828 2884
rect -9762 2864 -9732 2884
rect -9666 2864 -9636 2884
rect -9570 2864 -9540 2884
rect -9474 2864 -9444 2884
rect -9378 2864 -9348 2884
rect -9282 2864 -9252 2884
rect -9186 2864 -9156 2884
rect -9090 2864 -9060 2884
rect -8994 2864 -8964 2884
rect -8898 2864 -8868 2884
rect -8802 2864 -8772 2884
rect -8706 2864 -8676 2884
rect -8610 2864 -8580 2884
rect -8514 2864 -8484 2884
rect -8418 2864 -8388 2884
rect -8322 2864 -8292 2884
rect -7998 2874 -6624 2906
rect -14464 1832 -14434 1858
rect -14368 1832 -14338 1858
rect -14272 1832 -14242 1858
rect -14176 1832 -14146 1858
rect -14080 1832 -14050 1858
rect -13984 1832 -13954 1858
rect -13888 1832 -13858 1858
rect -13792 1832 -13762 1858
rect -13696 1832 -13666 1858
rect -13600 1832 -13570 1858
rect -13504 1832 -13474 1858
rect -13408 1832 -13378 1858
rect -13312 1832 -13282 1858
rect -13216 1832 -13186 1858
rect -13120 1832 -13090 1858
rect -12786 1836 -12756 1862
rect -12690 1836 -12660 1862
rect -12594 1836 -12564 1862
rect -12498 1836 -12468 1862
rect -12402 1836 -12372 1862
rect -12306 1836 -12276 1862
rect -12210 1836 -12180 1862
rect -12114 1836 -12084 1862
rect -12018 1836 -11988 1862
rect -11922 1836 -11892 1862
rect -11614 1846 -11584 1872
rect -11518 1846 -11488 1872
rect -11422 1846 -11392 1872
rect -11326 1846 -11296 1872
rect -11230 1846 -11200 1872
rect -7998 2856 -7968 2874
rect -7902 2856 -7872 2874
rect -7806 2856 -7776 2874
rect -7710 2856 -7680 2874
rect -7614 2856 -7584 2874
rect -7518 2856 -7488 2874
rect -7422 2856 -7392 2874
rect -7326 2856 -7296 2874
rect -7230 2856 -7200 2874
rect -7134 2856 -7104 2874
rect -7038 2856 -7008 2874
rect -6942 2856 -6912 2874
rect -6846 2856 -6816 2874
rect -6750 2856 -6720 2874
rect -6654 2856 -6624 2874
rect -6320 2876 -5426 2906
rect -6320 2860 -6290 2876
rect -6224 2860 -6194 2876
rect -6128 2860 -6098 2876
rect -6032 2860 -6002 2876
rect -5936 2860 -5906 2876
rect -5840 2860 -5810 2876
rect -5744 2860 -5714 2876
rect -5648 2860 -5618 2876
rect -5552 2860 -5522 2876
rect -5456 2860 -5426 2876
rect -5148 2892 -4734 2922
rect -5148 2870 -5118 2892
rect -5052 2870 -5022 2892
rect -4956 2870 -4926 2892
rect -4860 2870 -4830 2892
rect -4764 2870 -4734 2892
rect -10146 1838 -10116 1864
rect -10050 1838 -10020 1864
rect -9954 1838 -9924 1864
rect -9858 1838 -9828 1864
rect -9762 1838 -9732 1864
rect -9666 1838 -9636 1864
rect -9570 1838 -9540 1864
rect -9474 1838 -9444 1864
rect -9378 1838 -9348 1864
rect -9282 1838 -9252 1864
rect -9186 1838 -9156 1864
rect -9090 1838 -9060 1864
rect -8994 1838 -8964 1864
rect -8898 1838 -8868 1864
rect -8802 1838 -8772 1864
rect -8706 1838 -8676 1864
rect -8610 1838 -8580 1864
rect -8514 1838 -8484 1864
rect -8418 1838 -8388 1864
rect -8322 1838 -8292 1864
rect 1562 3002 1628 3018
rect 1562 2968 1578 3002
rect 1612 2968 1628 3002
rect 1562 2952 1628 2968
rect 1598 2922 1628 2952
rect 4518 2986 4584 3002
rect 4518 2952 4534 2986
rect 4568 2952 4584 2986
rect 4518 2936 4584 2952
rect 7548 2986 7614 3002
rect 7548 2952 7564 2986
rect 7598 2952 7614 2986
rect 7548 2936 7614 2952
rect 1598 2892 1658 2922
rect 4554 2906 4584 2936
rect 7584 2906 7614 2936
rect 10636 2984 10702 3000
rect 10636 2950 10652 2984
rect 10686 2950 10702 2984
rect 10636 2934 10702 2950
rect 1532 2862 1850 2892
rect 4554 2876 4614 2906
rect 7584 2876 7644 2906
rect 10672 2904 10702 2934
rect 13792 2958 13858 2974
rect 13792 2924 13808 2958
rect 13842 2924 13858 2958
rect 13792 2908 13858 2924
rect 1532 2830 1562 2862
rect 1628 2830 1658 2862
rect 1724 2854 1850 2862
rect 1724 2830 1754 2854
rect 1820 2830 1850 2854
rect 4488 2846 4806 2876
rect -1636 2210 -1606 2236
rect -1540 2210 -1510 2236
rect -1444 2210 -1414 2236
rect -1348 2210 -1318 2236
rect -1252 2210 -1222 2236
rect -1156 2210 -1126 2236
rect -1060 2210 -1030 2236
rect -964 2210 -934 2236
rect -7998 1830 -7968 1856
rect -7902 1830 -7872 1856
rect -7806 1830 -7776 1856
rect -7710 1830 -7680 1856
rect -7614 1830 -7584 1856
rect -7518 1830 -7488 1856
rect -7422 1830 -7392 1856
rect -7326 1830 -7296 1856
rect -7230 1830 -7200 1856
rect -7134 1830 -7104 1856
rect -7038 1830 -7008 1856
rect -6942 1830 -6912 1856
rect -6846 1830 -6816 1856
rect -6750 1830 -6720 1856
rect -6654 1830 -6624 1856
rect -6320 1834 -6290 1860
rect -6224 1834 -6194 1860
rect -6128 1834 -6098 1860
rect -6032 1834 -6002 1860
rect -5936 1834 -5906 1860
rect -5840 1834 -5810 1860
rect -5744 1834 -5714 1860
rect -5648 1834 -5618 1860
rect -5552 1834 -5522 1860
rect -5456 1834 -5426 1860
rect -5148 1844 -5118 1870
rect -5052 1844 -5022 1870
rect -4956 1844 -4926 1870
rect -4860 1844 -4830 1870
rect -4764 1844 -4734 1870
rect 4488 2814 4518 2846
rect 4584 2814 4614 2846
rect 4680 2838 4806 2846
rect 4680 2814 4710 2838
rect 4776 2814 4806 2838
rect 7518 2846 7836 2876
rect 10672 2874 10732 2904
rect 13828 2878 13858 2908
rect 7518 2814 7548 2846
rect 7614 2814 7644 2846
rect 7710 2838 7836 2846
rect 7710 2814 7740 2838
rect 7806 2814 7836 2838
rect 10606 2844 10924 2874
rect 13828 2848 13888 2878
rect 2546 2428 2646 2444
rect 2546 2394 2579 2428
rect 2613 2394 2646 2428
rect 2546 2276 2646 2394
rect 2546 2050 2646 2076
rect 1532 1804 1562 1830
rect 1628 1804 1658 1830
rect 1724 1804 1754 1830
rect 1820 1804 1850 1830
rect 5546 2428 5646 2444
rect 5546 2394 5579 2428
rect 5613 2394 5646 2428
rect 5546 2276 5646 2394
rect 5546 2050 5646 2076
rect 10606 2812 10636 2844
rect 10702 2812 10732 2844
rect 10798 2836 10924 2844
rect 10798 2812 10828 2836
rect 10894 2812 10924 2836
rect 13762 2818 14080 2848
rect 8546 2428 8646 2444
rect 8546 2394 8579 2428
rect 8613 2394 8646 2428
rect 8546 2276 8646 2394
rect 8546 2050 8646 2076
rect 4488 1788 4518 1814
rect 4584 1788 4614 1814
rect 4680 1788 4710 1814
rect 4776 1788 4806 1814
rect 7518 1788 7548 1814
rect 7614 1788 7644 1814
rect 7710 1788 7740 1814
rect 7806 1788 7836 1814
rect 13762 2786 13792 2818
rect 13858 2786 13888 2818
rect 13954 2810 14080 2818
rect 13954 2786 13984 2810
rect 14050 2786 14080 2810
rect 11546 2428 11646 2444
rect 11546 2394 11579 2428
rect 11613 2394 11646 2428
rect 11546 2276 11646 2394
rect 11546 2050 11646 2076
rect 10606 1786 10636 1812
rect 10702 1786 10732 1812
rect 10798 1786 10828 1812
rect 10894 1786 10924 1812
rect 17428 3524 17458 3540
rect 17524 3524 17554 3540
rect 17620 3524 17650 3540
rect 17716 3524 17746 3540
rect 17812 3524 17842 3540
rect 17908 3524 17938 3540
rect 18004 3524 18034 3540
rect 18100 3524 18130 3540
rect 18196 3524 18226 3540
rect 18292 3524 18322 3540
rect 18626 3538 20000 3570
rect 16736 2508 16766 2534
rect 16832 2508 16862 2534
rect 16928 2508 16958 2534
rect 17024 2508 17054 2534
rect 17120 2508 17150 2534
rect 18626 3520 18656 3538
rect 18722 3520 18752 3538
rect 18818 3520 18848 3538
rect 18914 3520 18944 3538
rect 19010 3520 19040 3538
rect 19106 3520 19136 3538
rect 19202 3520 19232 3538
rect 19298 3520 19328 3538
rect 19394 3520 19424 3538
rect 19490 3520 19520 3538
rect 19586 3520 19616 3538
rect 19682 3520 19712 3538
rect 19778 3520 19808 3538
rect 19874 3520 19904 3538
rect 19970 3520 20000 3538
rect 20294 3548 22148 3578
rect 20294 3528 20324 3548
rect 20390 3528 20420 3548
rect 20486 3528 20516 3548
rect 20582 3528 20612 3548
rect 20678 3528 20708 3548
rect 20774 3528 20804 3548
rect 20870 3528 20900 3548
rect 20966 3528 20996 3548
rect 21062 3528 21092 3548
rect 21158 3528 21188 3548
rect 21254 3528 21284 3548
rect 21350 3528 21380 3548
rect 21446 3528 21476 3548
rect 21542 3528 21572 3548
rect 21638 3528 21668 3548
rect 21734 3528 21764 3548
rect 21830 3528 21860 3548
rect 21926 3528 21956 3548
rect 22022 3528 22052 3548
rect 22118 3528 22148 3548
rect 23224 3554 23638 3584
rect 24012 3568 24042 3684
rect 25192 3656 25208 3690
rect 25242 3656 25258 3690
rect 25192 3640 25258 3656
rect 26860 3688 26926 3704
rect 26860 3654 26876 3688
rect 26910 3654 26926 3688
rect 25210 3568 25240 3640
rect 26860 3638 26926 3654
rect 26878 3576 26908 3638
rect 23224 3532 23254 3554
rect 23320 3532 23350 3554
rect 23416 3532 23446 3554
rect 23512 3532 23542 3554
rect 23608 3532 23638 3554
rect 23916 3538 24810 3568
rect 17428 2498 17458 2524
rect 17524 2498 17554 2524
rect 17620 2498 17650 2524
rect 17716 2498 17746 2524
rect 17812 2498 17842 2524
rect 17908 2498 17938 2524
rect 18004 2498 18034 2524
rect 18100 2498 18130 2524
rect 18196 2498 18226 2524
rect 18292 2498 18322 2524
rect 23916 3522 23946 3538
rect 24012 3522 24042 3538
rect 24108 3522 24138 3538
rect 24204 3522 24234 3538
rect 24300 3522 24330 3538
rect 24396 3522 24426 3538
rect 24492 3522 24522 3538
rect 24588 3522 24618 3538
rect 24684 3522 24714 3538
rect 24780 3522 24810 3538
rect 25114 3536 26488 3568
rect 18626 2494 18656 2520
rect 18722 2494 18752 2520
rect 18818 2494 18848 2520
rect 18914 2494 18944 2520
rect 19010 2494 19040 2520
rect 19106 2494 19136 2520
rect 19202 2494 19232 2520
rect 19298 2494 19328 2520
rect 19394 2494 19424 2520
rect 19490 2494 19520 2520
rect 19586 2494 19616 2520
rect 19682 2494 19712 2520
rect 19778 2494 19808 2520
rect 19874 2494 19904 2520
rect 19970 2494 20000 2520
rect 20294 2502 20324 2528
rect 20390 2502 20420 2528
rect 20486 2502 20516 2528
rect 20582 2502 20612 2528
rect 20678 2502 20708 2528
rect 20774 2502 20804 2528
rect 20870 2502 20900 2528
rect 20966 2502 20996 2528
rect 21062 2502 21092 2528
rect 21158 2502 21188 2528
rect 21254 2502 21284 2528
rect 21350 2502 21380 2528
rect 21446 2502 21476 2528
rect 21542 2502 21572 2528
rect 21638 2502 21668 2528
rect 21734 2502 21764 2528
rect 21830 2502 21860 2528
rect 21926 2502 21956 2528
rect 22022 2502 22052 2528
rect 22118 2502 22148 2528
rect 23224 2506 23254 2532
rect 23320 2506 23350 2532
rect 23416 2506 23446 2532
rect 23512 2506 23542 2532
rect 23608 2506 23638 2532
rect 25114 3518 25144 3536
rect 25210 3518 25240 3536
rect 25306 3518 25336 3536
rect 25402 3518 25432 3536
rect 25498 3518 25528 3536
rect 25594 3518 25624 3536
rect 25690 3518 25720 3536
rect 25786 3518 25816 3536
rect 25882 3518 25912 3536
rect 25978 3518 26008 3536
rect 26074 3518 26104 3536
rect 26170 3518 26200 3536
rect 26266 3518 26296 3536
rect 26362 3518 26392 3536
rect 26458 3518 26488 3536
rect 26782 3546 28636 3576
rect 26782 3526 26812 3546
rect 26878 3526 26908 3546
rect 26974 3526 27004 3546
rect 27070 3526 27100 3546
rect 27166 3526 27196 3546
rect 27262 3526 27292 3546
rect 27358 3526 27388 3546
rect 27454 3526 27484 3546
rect 27550 3526 27580 3546
rect 27646 3526 27676 3546
rect 27742 3526 27772 3546
rect 27838 3526 27868 3546
rect 27934 3526 27964 3546
rect 28030 3526 28060 3546
rect 28126 3526 28156 3546
rect 28222 3526 28252 3546
rect 28318 3526 28348 3546
rect 28414 3526 28444 3546
rect 28510 3526 28540 3546
rect 28606 3526 28636 3546
rect 23916 2496 23946 2522
rect 24012 2496 24042 2522
rect 24108 2496 24138 2522
rect 24204 2496 24234 2522
rect 24300 2496 24330 2522
rect 24396 2496 24426 2522
rect 24492 2496 24522 2522
rect 24588 2496 24618 2522
rect 24684 2496 24714 2522
rect 24780 2496 24810 2522
rect 25114 2492 25144 2518
rect 25210 2492 25240 2518
rect 25306 2492 25336 2518
rect 25402 2492 25432 2518
rect 25498 2492 25528 2518
rect 25594 2492 25624 2518
rect 25690 2492 25720 2518
rect 25786 2492 25816 2518
rect 25882 2492 25912 2518
rect 25978 2492 26008 2518
rect 26074 2492 26104 2518
rect 26170 2492 26200 2518
rect 26266 2492 26296 2518
rect 26362 2492 26392 2518
rect 26458 2492 26488 2518
rect 26782 2500 26812 2526
rect 26878 2500 26908 2526
rect 26974 2500 27004 2526
rect 27070 2500 27100 2526
rect 27166 2500 27196 2526
rect 27262 2500 27292 2526
rect 27358 2500 27388 2526
rect 27454 2500 27484 2526
rect 27550 2500 27580 2526
rect 27646 2500 27676 2526
rect 27742 2500 27772 2526
rect 27838 2500 27868 2526
rect 27934 2500 27964 2526
rect 28030 2500 28060 2526
rect 28126 2500 28156 2526
rect 28222 2500 28252 2526
rect 28318 2500 28348 2526
rect 28414 2500 28444 2526
rect 28510 2500 28540 2526
rect 28606 2500 28636 2526
rect 14546 2428 14646 2444
rect 14546 2394 14579 2428
rect 14613 2394 14646 2428
rect 14546 2276 14646 2394
rect 14546 2050 14646 2076
rect 13762 1760 13792 1786
rect 13858 1760 13888 1786
rect 13954 1760 13984 1786
rect 14050 1760 14080 1786
rect 15450 1492 15516 1508
rect 15450 1458 15466 1492
rect 15500 1458 15516 1492
rect 15450 1442 15516 1458
rect -1111 1298 -1045 1314
rect -1111 1264 -1095 1298
rect -1061 1264 -1045 1298
rect -1111 1248 -1045 1264
rect -915 1298 -849 1314
rect -915 1264 -899 1298
rect -865 1264 -849 1298
rect 208 1306 1294 1336
rect 208 1268 238 1306
rect 304 1268 334 1306
rect 400 1268 430 1306
rect 496 1268 526 1306
rect 592 1268 622 1306
rect 688 1268 718 1306
rect 784 1268 814 1306
rect 880 1268 910 1306
rect 976 1268 1006 1306
rect 1072 1268 1102 1306
rect 1168 1268 1198 1306
rect 1264 1268 1294 1306
rect 1976 1310 2966 1340
rect 1976 1268 2006 1310
rect 2072 1268 2102 1310
rect 2168 1268 2198 1310
rect 2264 1268 2294 1310
rect 2360 1268 2390 1310
rect 2456 1268 2486 1310
rect 2552 1268 2582 1310
rect 2648 1268 2678 1310
rect 2744 1268 2774 1310
rect 2840 1268 2870 1310
rect 2936 1268 2966 1310
rect 3164 1290 4250 1320
rect -915 1248 -849 1264
rect -1100 1180 -1060 1248
rect -904 1180 -864 1248
rect -1640 1140 -858 1180
rect -1640 1066 -1600 1140
rect -1542 1066 -1502 1140
rect -1444 1066 -1404 1140
rect -1346 1066 -1306 1140
rect -1248 1066 -1208 1140
rect -1150 1066 -1110 1140
rect -1052 1066 -1012 1140
rect -954 1066 -914 1140
rect 3164 1252 3194 1290
rect 3260 1252 3290 1290
rect 3356 1252 3386 1290
rect 3452 1252 3482 1290
rect 3548 1252 3578 1290
rect 3644 1252 3674 1290
rect 3740 1252 3770 1290
rect 3836 1252 3866 1290
rect 3932 1252 3962 1290
rect 4028 1252 4058 1290
rect 4124 1252 4154 1290
rect 4220 1252 4250 1290
rect 4932 1294 5922 1324
rect 4932 1252 4962 1294
rect 5028 1252 5058 1294
rect 5124 1252 5154 1294
rect 5220 1252 5250 1294
rect 5316 1252 5346 1294
rect 5412 1252 5442 1294
rect 5508 1252 5538 1294
rect 5604 1252 5634 1294
rect 5700 1252 5730 1294
rect 5796 1252 5826 1294
rect 5892 1252 5922 1294
rect 6194 1290 7280 1320
rect 6194 1252 6224 1290
rect 6290 1252 6320 1290
rect 6386 1252 6416 1290
rect 6482 1252 6512 1290
rect 6578 1252 6608 1290
rect 6674 1252 6704 1290
rect 6770 1252 6800 1290
rect 6866 1252 6896 1290
rect 6962 1252 6992 1290
rect 7058 1252 7088 1290
rect 7154 1252 7184 1290
rect 7250 1252 7280 1290
rect 7962 1294 8952 1324
rect 7962 1252 7992 1294
rect 8058 1252 8088 1294
rect 8154 1252 8184 1294
rect 8250 1252 8280 1294
rect 8346 1252 8376 1294
rect 8442 1252 8472 1294
rect 8538 1252 8568 1294
rect 8634 1252 8664 1294
rect 8730 1252 8760 1294
rect 8826 1252 8856 1294
rect 8922 1252 8952 1294
rect 9282 1288 10368 1318
rect 208 214 238 268
rect 304 242 334 268
rect 400 242 430 268
rect 496 242 526 268
rect 592 242 622 268
rect 688 242 718 268
rect 784 242 814 268
rect 880 242 910 268
rect 976 242 1006 268
rect 1072 242 1102 268
rect 1168 242 1198 268
rect 1264 242 1294 268
rect 1976 242 2006 268
rect 2072 242 2102 268
rect 2168 242 2198 268
rect 2264 242 2294 268
rect 2360 242 2390 268
rect 2456 242 2486 268
rect 2552 242 2582 268
rect 2648 242 2678 268
rect 176 184 238 214
rect 2744 208 2774 268
rect 2840 242 2870 268
rect 2936 242 2966 268
rect 9282 1250 9312 1288
rect 9378 1250 9408 1288
rect 9474 1250 9504 1288
rect 9570 1250 9600 1288
rect 9666 1250 9696 1288
rect 9762 1250 9792 1288
rect 9858 1250 9888 1288
rect 9954 1250 9984 1288
rect 10050 1250 10080 1288
rect 10146 1250 10176 1288
rect 10242 1250 10272 1288
rect 10338 1250 10368 1288
rect 11050 1292 12040 1322
rect 15468 1300 15498 1442
rect 11050 1250 11080 1292
rect 11146 1250 11176 1292
rect 11242 1250 11272 1292
rect 11338 1250 11368 1292
rect 11434 1250 11464 1292
rect 11530 1250 11560 1292
rect 11626 1250 11656 1292
rect 11722 1250 11752 1292
rect 11818 1250 11848 1292
rect 11914 1250 11944 1292
rect 12010 1250 12040 1292
rect 12438 1262 13524 1292
rect 176 146 206 184
rect 2744 178 2802 208
rect 3164 198 3194 252
rect 3260 226 3290 252
rect 3356 226 3386 252
rect 3452 226 3482 252
rect 3548 226 3578 252
rect 3644 226 3674 252
rect 3740 226 3770 252
rect 3836 226 3866 252
rect 3932 226 3962 252
rect 4028 226 4058 252
rect 4124 226 4154 252
rect 4220 226 4250 252
rect 4932 226 4962 252
rect 5028 226 5058 252
rect 5124 226 5154 252
rect 5220 226 5250 252
rect 5316 226 5346 252
rect 5412 226 5442 252
rect 5508 226 5538 252
rect 5604 226 5634 252
rect 140 130 206 146
rect 140 96 156 130
rect 190 96 206 130
rect 140 80 206 96
rect 2772 146 2802 178
rect 3132 168 3194 198
rect 5700 192 5730 252
rect 5796 226 5826 252
rect 5892 226 5922 252
rect 6194 198 6224 252
rect 6290 226 6320 252
rect 6386 226 6416 252
rect 6482 226 6512 252
rect 6578 226 6608 252
rect 6674 226 6704 252
rect 6770 226 6800 252
rect 6866 226 6896 252
rect 6962 226 6992 252
rect 7058 226 7088 252
rect 7154 226 7184 252
rect 7250 226 7280 252
rect 7962 226 7992 252
rect 8058 226 8088 252
rect 8154 226 8184 252
rect 8250 226 8280 252
rect 8346 226 8376 252
rect 8442 226 8472 252
rect 8538 226 8568 252
rect 8634 226 8664 252
rect 2772 130 2838 146
rect 3132 130 3162 168
rect 5700 162 5758 192
rect 2772 96 2788 130
rect 2822 96 2838 130
rect 2772 80 2838 96
rect 3096 114 3162 130
rect 3096 80 3112 114
rect 3146 80 3162 114
rect -1640 40 -1600 66
rect -1542 40 -1502 66
rect -1444 40 -1404 66
rect -1346 40 -1306 66
rect -1248 40 -1208 66
rect -1150 40 -1110 66
rect -1052 40 -1012 66
rect -954 40 -914 66
rect 3096 64 3162 80
rect 5728 130 5758 162
rect 6162 168 6224 198
rect 8730 192 8760 252
rect 8826 226 8856 252
rect 8922 226 8952 252
rect 12438 1224 12468 1262
rect 12534 1224 12564 1262
rect 12630 1224 12660 1262
rect 12726 1224 12756 1262
rect 12822 1224 12852 1262
rect 12918 1224 12948 1262
rect 13014 1224 13044 1262
rect 13110 1224 13140 1262
rect 13206 1224 13236 1262
rect 13302 1224 13332 1262
rect 13398 1224 13428 1262
rect 13494 1224 13524 1262
rect 14206 1266 15196 1296
rect 14206 1224 14236 1266
rect 14302 1224 14332 1266
rect 14398 1224 14428 1266
rect 14494 1224 14524 1266
rect 14590 1224 14620 1266
rect 14686 1224 14716 1266
rect 14782 1224 14812 1266
rect 14878 1224 14908 1266
rect 14974 1224 15004 1266
rect 15070 1224 15100 1266
rect 15166 1224 15196 1266
rect 9282 196 9312 250
rect 9378 224 9408 250
rect 9474 224 9504 250
rect 9570 224 9600 250
rect 9666 224 9696 250
rect 9762 224 9792 250
rect 9858 224 9888 250
rect 9954 224 9984 250
rect 10050 224 10080 250
rect 10146 224 10176 250
rect 10242 224 10272 250
rect 10338 224 10368 250
rect 11050 224 11080 250
rect 11146 224 11176 250
rect 11242 224 11272 250
rect 11338 224 11368 250
rect 11434 224 11464 250
rect 11530 224 11560 250
rect 11626 224 11656 250
rect 11722 224 11752 250
rect 6162 130 6192 168
rect 8730 162 8788 192
rect 5728 114 5794 130
rect 5728 80 5744 114
rect 5778 80 5794 114
rect 5728 64 5794 80
rect 6126 114 6192 130
rect 6126 80 6142 114
rect 6176 80 6192 114
rect 6126 64 6192 80
rect 8758 130 8788 162
rect 9250 166 9312 196
rect 11818 190 11848 250
rect 11914 224 11944 250
rect 12010 224 12040 250
rect 8758 114 8824 130
rect 9250 128 9280 166
rect 11818 160 11876 190
rect 12438 170 12468 224
rect 12534 198 12564 224
rect 12630 198 12660 224
rect 12726 198 12756 224
rect 12822 198 12852 224
rect 12918 198 12948 224
rect 13014 198 13044 224
rect 13110 198 13140 224
rect 13206 198 13236 224
rect 13302 198 13332 224
rect 13398 198 13428 224
rect 13494 198 13524 224
rect 14206 198 14236 224
rect 14302 198 14332 224
rect 14398 198 14428 224
rect 14494 198 14524 224
rect 14590 198 14620 224
rect 14686 198 14716 224
rect 14782 198 14812 224
rect 14878 198 14908 224
rect 8758 80 8774 114
rect 8808 80 8824 114
rect 8758 64 8824 80
rect 9214 112 9280 128
rect 9214 78 9230 112
rect 9264 78 9280 112
rect 9214 62 9280 78
rect 11846 128 11876 160
rect 12406 140 12468 170
rect 14974 164 15004 224
rect 15070 198 15100 224
rect 15166 198 15196 224
rect 11846 112 11912 128
rect 11846 78 11862 112
rect 11896 78 11912 112
rect 12406 102 12436 140
rect 14974 134 15032 164
rect 11846 62 11912 78
rect 12370 86 12436 102
rect 12370 52 12386 86
rect 12420 52 12436 86
rect 12370 36 12436 52
rect 15002 102 15032 134
rect 15002 86 15068 102
rect 15002 52 15018 86
rect 15052 52 15068 86
rect 15468 74 15498 100
rect 15002 36 15068 52
<< polycont >>
rect 288 6773 322 6807
rect 2728 6769 2762 6803
rect 3244 6757 3278 6791
rect 5684 6753 5718 6787
rect 6274 6757 6308 6791
rect 8714 6753 8748 6787
rect 9362 6755 9396 6789
rect 11802 6751 11836 6785
rect 12518 6729 12552 6763
rect 14958 6725 14992 6759
rect -1067 4735 -1033 4769
rect -21714 3241 -21680 3275
rect -20050 3247 -20016 3281
rect -18846 3253 -18812 3287
rect 1580 3743 1614 3777
rect 1772 3743 1806 3777
rect 4536 3727 4570 3761
rect 4728 3727 4762 3761
rect 7566 3727 7600 3761
rect 16830 3909 16864 3943
rect 17518 3927 17552 3961
rect 18722 3921 18756 3955
rect 20386 3915 20420 3949
rect 23318 3907 23352 3941
rect 24006 3925 24040 3959
rect 25210 3919 25244 3953
rect 26874 3913 26908 3947
rect 7758 3727 7792 3761
rect 10654 3725 10688 3759
rect 10846 3725 10880 3759
rect 13810 3699 13844 3733
rect 14002 3699 14036 3733
rect 15566 3745 15600 3779
rect 16830 3672 16864 3706
rect 17522 3702 17556 3736
rect 18720 3658 18754 3692
rect 20388 3656 20422 3690
rect 23318 3670 23352 3704
rect 24010 3700 24044 3734
rect -18158 3235 -18124 3269
rect -14884 3253 -14850 3287
rect -13220 3259 -13186 3293
rect -12016 3265 -11982 3299
rect -11328 3247 -11294 3281
rect -8418 3251 -8384 3285
rect -6754 3257 -6720 3291
rect -5550 3263 -5516 3297
rect -1590 3394 -1556 3428
rect -4862 3245 -4828 3279
rect -21716 2982 -21682 3016
rect -20048 2984 -20014 3018
rect -18850 3028 -18816 3062
rect -18158 2998 -18124 3032
rect -14886 2994 -14852 3028
rect -13218 2996 -13184 3030
rect -12020 3040 -11986 3074
rect -11328 3010 -11294 3044
rect -8420 2992 -8386 3026
rect -6752 2994 -6718 3028
rect -5554 3038 -5520 3072
rect -4862 3008 -4828 3042
rect 1578 2968 1612 3002
rect 4534 2952 4568 2986
rect 7564 2952 7598 2986
rect 10652 2950 10686 2984
rect 13808 2924 13842 2958
rect 2579 2394 2613 2428
rect 5579 2394 5613 2428
rect 8579 2394 8613 2428
rect 11579 2394 11613 2428
rect 25208 3656 25242 3690
rect 26876 3654 26910 3688
rect 14579 2394 14613 2428
rect 15466 1458 15500 1492
rect -1095 1264 -1061 1298
rect -899 1264 -865 1298
rect 156 96 190 130
rect 2788 96 2822 130
rect 3112 80 3146 114
rect 5744 80 5778 114
rect 6142 80 6176 114
rect 8774 80 8808 114
rect 9230 78 9264 112
rect 11862 78 11896 112
rect 12386 52 12420 86
rect 15018 52 15052 86
<< locali >>
rect 15414 9057 15674 9088
rect -356 9022 -154 9030
rect -356 8972 -344 9022
rect -380 8844 -344 8972
rect -166 8972 -154 9022
rect 1644 9022 1846 9030
rect 1644 8972 1656 9022
rect -166 8844 -122 8972
rect -380 8180 -122 8844
rect 1620 8844 1656 8972
rect 1834 8972 1846 9022
rect 3644 9022 3846 9030
rect 3644 8972 3656 9022
rect 1834 8844 1878 8972
rect 1620 8180 1878 8844
rect 3620 8844 3656 8972
rect 3834 8972 3846 9022
rect 5644 9022 5846 9030
rect 5644 8972 5656 9022
rect 3834 8844 3878 8972
rect 3620 8180 3878 8844
rect 5620 8844 5656 8972
rect 5834 8972 5846 9022
rect 7644 9022 7846 9030
rect 7644 8972 7656 9022
rect 5834 8844 5878 8972
rect 5620 8180 5878 8844
rect 7620 8844 7656 8972
rect 7834 8972 7846 9022
rect 9644 9022 9846 9030
rect 9644 8972 9656 9022
rect 7834 8844 7878 8972
rect 7620 8180 7878 8844
rect 9620 8844 9656 8972
rect 9834 8972 9846 9022
rect 11644 9022 11846 9030
rect 11644 8972 11656 9022
rect 9834 8844 9878 8972
rect 9620 8180 9878 8844
rect 11620 8844 11656 8972
rect 11834 8972 11846 9022
rect 13644 9022 13846 9030
rect 13644 8972 13656 9022
rect 11834 8844 11878 8972
rect 11620 8180 11878 8844
rect 13620 8844 13656 8972
rect 13834 8972 13846 9022
rect 13834 8844 13878 8972
rect 13620 8180 13878 8844
rect 15414 8879 15454 9057
rect 15632 8879 15674 9057
rect 15414 8842 15674 8879
rect 15414 8180 15672 8842
rect -1364 8157 15832 8180
rect -1364 7851 -1317 8157
rect 15785 7851 15832 8157
rect -1364 7828 15832 7851
rect -262 6728 -142 7828
rect 1662 6896 1912 7828
rect 272 6773 288 6807
rect 322 6773 338 6807
rect 764 6728 798 6858
rect 1662 6792 1694 6896
rect 1888 6792 1912 6896
rect 4522 6880 4772 7828
rect 1662 6758 1912 6792
rect 2712 6769 2728 6803
rect 2762 6769 2778 6803
rect 3228 6757 3244 6791
rect 3278 6757 3294 6791
rect -1190 6644 1392 6728
rect 2440 6702 2474 6754
rect 1960 6668 2768 6702
rect 3720 6684 3754 6842
rect 4522 6776 4552 6880
rect 4746 6776 4772 6880
rect 7456 6878 7706 7828
rect 4522 6762 4772 6776
rect 5668 6753 5684 6787
rect 5718 6753 5734 6787
rect 6258 6757 6274 6791
rect 6308 6757 6324 6791
rect 5396 6686 5430 6738
rect -1188 6042 -1102 6644
rect 194 6591 228 6644
rect 194 6519 228 6531
rect 194 6447 228 6463
rect 194 6375 228 6395
rect 194 6303 228 6327
rect 194 6231 228 6259
rect 194 6159 228 6191
rect 194 6089 228 6123
rect -1652 6006 -834 6042
rect -1652 5921 -1618 6006
rect -1652 5849 -1618 5861
rect -1652 5777 -1618 5793
rect -1652 5705 -1618 5725
rect -1652 5633 -1618 5657
rect -1652 5561 -1618 5589
rect -1652 5489 -1618 5521
rect -1652 5419 -1618 5453
rect -1652 5351 -1618 5383
rect -1652 5283 -1618 5311
rect -1652 5215 -1618 5239
rect -1652 5147 -1618 5167
rect -1652 5079 -1618 5095
rect -1652 5011 -1618 5023
rect -1652 4932 -1618 4951
rect -1554 5921 -1520 5938
rect -1554 5849 -1520 5861
rect -1554 5777 -1520 5793
rect -1554 5705 -1520 5725
rect -1554 5633 -1520 5657
rect -1554 5561 -1520 5589
rect -1554 5489 -1520 5521
rect -1554 5419 -1520 5453
rect -1554 5351 -1520 5383
rect -1554 5283 -1520 5311
rect -1554 5215 -1520 5239
rect -1554 5147 -1520 5167
rect -1554 5079 -1520 5095
rect -1554 5011 -1520 5023
rect -1554 4876 -1520 4951
rect -1456 5921 -1422 6006
rect -1456 5849 -1422 5861
rect -1456 5777 -1422 5793
rect -1456 5705 -1422 5725
rect -1456 5633 -1422 5657
rect -1456 5561 -1422 5589
rect -1456 5489 -1422 5521
rect -1456 5419 -1422 5453
rect -1456 5351 -1422 5383
rect -1456 5283 -1422 5311
rect -1456 5215 -1422 5239
rect -1456 5147 -1422 5167
rect -1456 5079 -1422 5095
rect -1456 5011 -1422 5023
rect -1456 4932 -1422 4951
rect -1358 5921 -1324 5938
rect -1358 5849 -1324 5861
rect -1358 5777 -1324 5793
rect -1358 5705 -1324 5725
rect -1358 5633 -1324 5657
rect -1358 5561 -1324 5589
rect -1358 5489 -1324 5521
rect -1358 5419 -1324 5453
rect -1358 5351 -1324 5383
rect -1358 5283 -1324 5311
rect -1358 5215 -1324 5239
rect -1358 5147 -1324 5167
rect -1358 5079 -1324 5095
rect -1358 5011 -1324 5023
rect -1358 4876 -1324 4951
rect -1260 5921 -1226 6006
rect -1260 5849 -1226 5861
rect -1260 5777 -1226 5793
rect -1260 5705 -1226 5725
rect -1260 5633 -1226 5657
rect -1260 5561 -1226 5589
rect -1260 5489 -1226 5521
rect -1260 5419 -1226 5453
rect -1260 5351 -1226 5383
rect -1260 5283 -1226 5311
rect -1260 5215 -1226 5239
rect -1260 5147 -1226 5167
rect -1260 5079 -1226 5095
rect -1260 5011 -1226 5023
rect -1260 4932 -1226 4951
rect -1162 5921 -1128 5938
rect -1162 5849 -1128 5861
rect -1162 5777 -1128 5793
rect -1162 5705 -1128 5725
rect -1162 5633 -1128 5657
rect -1162 5561 -1128 5589
rect -1162 5489 -1128 5521
rect -1162 5419 -1128 5453
rect -1162 5351 -1128 5383
rect -1162 5283 -1128 5311
rect -1162 5215 -1128 5239
rect -1162 5147 -1128 5167
rect -1162 5079 -1128 5095
rect -1162 5011 -1128 5023
rect -1162 4876 -1128 4951
rect -1064 5921 -1030 6006
rect -1064 5849 -1030 5861
rect -1064 5777 -1030 5793
rect -1064 5705 -1030 5725
rect -1064 5633 -1030 5657
rect -1064 5561 -1030 5589
rect -1064 5489 -1030 5521
rect -1064 5419 -1030 5453
rect -1064 5351 -1030 5383
rect -1064 5283 -1030 5311
rect -1064 5215 -1030 5239
rect -1064 5147 -1030 5167
rect -1064 5079 -1030 5095
rect -1064 5011 -1030 5023
rect -1064 4932 -1030 4951
rect -966 5921 -932 5938
rect -966 5849 -932 5861
rect -966 5777 -932 5793
rect -966 5705 -932 5725
rect -966 5633 -932 5657
rect -966 5561 -932 5589
rect -966 5489 -932 5521
rect -966 5419 -932 5453
rect -966 5351 -932 5383
rect -966 5283 -932 5311
rect -966 5215 -932 5239
rect -966 5147 -932 5167
rect -966 5079 -932 5095
rect -966 5011 -932 5023
rect -966 4876 -932 4951
rect -868 5921 -834 6006
rect -868 5849 -834 5861
rect -868 5777 -834 5793
rect -868 5705 -834 5725
rect -868 5633 -834 5657
rect 194 6021 228 6053
rect 194 5953 228 5981
rect 194 5885 228 5909
rect 194 5817 228 5837
rect 194 5749 228 5765
rect 194 5681 228 5693
rect 194 5602 228 5621
rect 290 6591 324 6608
rect 290 6519 324 6531
rect 290 6447 324 6463
rect 290 6375 324 6395
rect 290 6303 324 6327
rect 290 6231 324 6259
rect 290 6159 324 6191
rect 290 6089 324 6123
rect 290 6021 324 6053
rect 290 5953 324 5981
rect 290 5885 324 5909
rect 290 5817 324 5837
rect 290 5749 324 5765
rect 290 5681 324 5693
rect -868 5561 -834 5589
rect -868 5489 -834 5521
rect 290 5550 324 5621
rect 386 6591 420 6644
rect 386 6519 420 6531
rect 386 6447 420 6463
rect 386 6375 420 6395
rect 386 6303 420 6327
rect 386 6231 420 6259
rect 386 6159 420 6191
rect 386 6089 420 6123
rect 386 6021 420 6053
rect 386 5953 420 5981
rect 386 5885 420 5909
rect 386 5817 420 5837
rect 386 5749 420 5765
rect 386 5681 420 5693
rect 386 5604 420 5621
rect 482 6591 516 6608
rect 482 6519 516 6531
rect 482 6447 516 6463
rect 482 6375 516 6395
rect 482 6303 516 6327
rect 482 6231 516 6259
rect 482 6159 516 6191
rect 482 6089 516 6123
rect 482 6021 516 6053
rect 482 5953 516 5981
rect 482 5885 516 5909
rect 482 5817 516 5837
rect 482 5749 516 5765
rect 482 5681 516 5693
rect 482 5550 516 5621
rect 578 6591 612 6644
rect 578 6519 612 6531
rect 578 6447 612 6463
rect 578 6375 612 6395
rect 578 6303 612 6327
rect 578 6231 612 6259
rect 578 6159 612 6191
rect 578 6089 612 6123
rect 578 6021 612 6053
rect 578 5953 612 5981
rect 578 5885 612 5909
rect 578 5817 612 5837
rect 578 5749 612 5765
rect 578 5681 612 5693
rect 578 5604 612 5621
rect 674 6591 708 6608
rect 674 6519 708 6531
rect 674 6447 708 6463
rect 674 6375 708 6395
rect 674 6303 708 6327
rect 674 6231 708 6259
rect 674 6159 708 6191
rect 674 6089 708 6123
rect 674 6021 708 6053
rect 674 5953 708 5981
rect 674 5885 708 5909
rect 674 5817 708 5837
rect 674 5749 708 5765
rect 674 5681 708 5693
rect 674 5550 708 5621
rect 770 6591 804 6644
rect 770 6519 804 6531
rect 770 6447 804 6463
rect 770 6375 804 6395
rect 770 6303 804 6327
rect 770 6231 804 6259
rect 770 6159 804 6191
rect 770 6089 804 6123
rect 770 6021 804 6053
rect 770 5953 804 5981
rect 770 5885 804 5909
rect 770 5817 804 5837
rect 770 5749 804 5765
rect 770 5681 804 5693
rect 770 5604 804 5621
rect 866 6591 900 6608
rect 866 6519 900 6531
rect 866 6447 900 6463
rect 866 6375 900 6395
rect 866 6303 900 6327
rect 866 6231 900 6259
rect 866 6159 900 6191
rect 866 6089 900 6123
rect 866 6021 900 6053
rect 866 5953 900 5981
rect 866 5885 900 5909
rect 866 5817 900 5837
rect 866 5749 900 5765
rect 866 5681 900 5693
rect 866 5550 900 5621
rect 962 6591 996 6644
rect 962 6519 996 6531
rect 962 6447 996 6463
rect 962 6375 996 6395
rect 962 6303 996 6327
rect 962 6231 996 6259
rect 962 6159 996 6191
rect 962 6089 996 6123
rect 962 6021 996 6053
rect 962 5953 996 5981
rect 962 5885 996 5909
rect 962 5817 996 5837
rect 962 5749 996 5765
rect 962 5681 996 5693
rect 962 5604 996 5621
rect 1058 6591 1092 6608
rect 1058 6519 1092 6531
rect 1058 6447 1092 6463
rect 1058 6375 1092 6395
rect 1058 6303 1092 6327
rect 1058 6231 1092 6259
rect 1058 6159 1092 6191
rect 1058 6089 1092 6123
rect 1058 6021 1092 6053
rect 1058 5953 1092 5981
rect 1058 5885 1092 5909
rect 1058 5817 1092 5837
rect 1058 5749 1092 5765
rect 1058 5681 1092 5693
rect 1058 5550 1092 5621
rect 1154 6591 1188 6644
rect 1154 6519 1188 6531
rect 1154 6447 1188 6463
rect 1154 6375 1188 6395
rect 1154 6303 1188 6327
rect 1154 6231 1188 6259
rect 1154 6159 1188 6191
rect 1154 6089 1188 6123
rect 1154 6021 1188 6053
rect 1154 5953 1188 5981
rect 1154 5885 1188 5909
rect 1154 5817 1188 5837
rect 1154 5749 1188 5765
rect 1154 5681 1188 5693
rect 1154 5604 1188 5621
rect 1250 6591 1284 6608
rect 1250 6519 1284 6531
rect 1250 6447 1284 6463
rect 1250 6375 1284 6395
rect 1250 6303 1284 6327
rect 1250 6231 1284 6259
rect 1250 6159 1284 6191
rect 1250 6089 1284 6123
rect 1250 6021 1284 6053
rect 1250 5953 1284 5981
rect 1250 5885 1284 5909
rect 1250 5817 1284 5837
rect 1250 5749 1284 5765
rect 1250 5681 1284 5693
rect 1250 5550 1284 5621
rect 1346 6591 1380 6644
rect 1346 6519 1380 6531
rect 1346 6447 1380 6463
rect 1346 6375 1380 6395
rect 1346 6303 1380 6327
rect 1346 6231 1380 6259
rect 1346 6159 1380 6191
rect 1346 6089 1380 6123
rect 1346 6021 1380 6053
rect 1346 5953 1380 5981
rect 1346 5885 1380 5909
rect 1346 5817 1380 5837
rect 1346 5749 1380 5765
rect 1346 5681 1380 5693
rect 1346 5604 1380 5621
rect 1960 6587 1994 6668
rect 1960 6515 1994 6527
rect 1960 6443 1994 6459
rect 1960 6371 1994 6391
rect 1960 6299 1994 6323
rect 1960 6227 1994 6255
rect 1960 6155 1994 6187
rect 1960 6085 1994 6119
rect 1960 6017 1994 6049
rect 1960 5949 1994 5977
rect 1960 5881 1994 5905
rect 1960 5813 1994 5833
rect 1960 5745 1994 5761
rect 1960 5677 1994 5689
rect 1960 5598 1994 5617
rect 2056 6587 2090 6604
rect 2056 6515 2090 6527
rect 2056 6443 2090 6459
rect 2056 6371 2090 6391
rect 2056 6299 2090 6323
rect 2056 6227 2090 6255
rect 2056 6155 2090 6187
rect 2056 6085 2090 6119
rect 2056 6017 2090 6049
rect 2056 5949 2090 5977
rect 2056 5881 2090 5905
rect 2056 5813 2090 5833
rect 2056 5745 2090 5761
rect 2056 5677 2090 5689
rect 290 5516 1284 5550
rect 2056 5548 2090 5617
rect 2152 6587 2186 6668
rect 2152 6515 2186 6527
rect 2152 6443 2186 6459
rect 2152 6371 2186 6391
rect 2152 6299 2186 6323
rect 2152 6227 2186 6255
rect 2152 6155 2186 6187
rect 2152 6085 2186 6119
rect 2152 6017 2186 6049
rect 2152 5949 2186 5977
rect 2152 5881 2186 5905
rect 2152 5813 2186 5833
rect 2152 5745 2186 5761
rect 2152 5677 2186 5689
rect 2152 5598 2186 5617
rect 2248 6587 2282 6604
rect 2248 6515 2282 6527
rect 2248 6443 2282 6459
rect 2248 6371 2282 6391
rect 2248 6299 2282 6323
rect 2248 6227 2282 6255
rect 2248 6155 2282 6187
rect 2248 6085 2282 6119
rect 2248 6017 2282 6049
rect 2248 5949 2282 5977
rect 2248 5881 2282 5905
rect 2248 5813 2282 5833
rect 2248 5745 2282 5761
rect 2248 5677 2282 5689
rect 2248 5548 2282 5617
rect 2344 6587 2378 6668
rect 2344 6515 2378 6527
rect 2344 6443 2378 6459
rect 2344 6371 2378 6391
rect 2344 6299 2378 6323
rect 2344 6227 2378 6255
rect 2344 6155 2378 6187
rect 2344 6085 2378 6119
rect 2344 6017 2378 6049
rect 2344 5949 2378 5977
rect 2344 5881 2378 5905
rect 2344 5813 2378 5833
rect 2344 5745 2378 5761
rect 2344 5677 2378 5689
rect 2344 5598 2378 5617
rect 2440 6587 2474 6604
rect 2440 6515 2474 6527
rect 2440 6443 2474 6459
rect 2440 6371 2474 6391
rect 2440 6299 2474 6323
rect 2440 6227 2474 6255
rect 2440 6155 2474 6187
rect 2440 6085 2474 6119
rect 2440 6017 2474 6049
rect 2440 5949 2474 5977
rect 2440 5881 2474 5905
rect 2440 5813 2474 5833
rect 2440 5745 2474 5761
rect 2440 5677 2474 5689
rect 2440 5548 2474 5617
rect 2536 6587 2570 6668
rect 2536 6515 2570 6527
rect 2536 6443 2570 6459
rect 2536 6371 2570 6391
rect 2536 6299 2570 6323
rect 2536 6227 2570 6255
rect 2536 6155 2570 6187
rect 2536 6085 2570 6119
rect 2536 6017 2570 6049
rect 2536 5949 2570 5977
rect 2536 5881 2570 5905
rect 2536 5813 2570 5833
rect 2536 5745 2570 5761
rect 2536 5677 2570 5689
rect 2536 5598 2570 5617
rect 2632 6587 2666 6604
rect 2632 6515 2666 6527
rect 2632 6443 2666 6459
rect 2632 6371 2666 6391
rect 2632 6299 2666 6323
rect 2632 6227 2666 6255
rect 2632 6155 2666 6187
rect 2632 6085 2666 6119
rect 2632 6017 2666 6049
rect 2632 5949 2666 5977
rect 2632 5881 2666 5905
rect 2632 5813 2666 5833
rect 2632 5745 2666 5761
rect 2632 5677 2666 5689
rect 2632 5548 2666 5617
rect 2728 6587 2762 6668
rect 2728 6515 2762 6527
rect 2728 6443 2762 6459
rect 2728 6371 2762 6391
rect 2728 6299 2762 6323
rect 2728 6227 2762 6255
rect 2728 6155 2762 6187
rect 2728 6085 2762 6119
rect 2728 6017 2762 6049
rect 2728 5949 2762 5977
rect 2728 5881 2762 5905
rect 2728 5813 2762 5833
rect 2728 5745 2762 5761
rect 2728 5677 2762 5689
rect 2728 5600 2762 5617
rect 3150 6650 4344 6684
rect 4916 6652 5724 6686
rect 6750 6684 6784 6842
rect 7456 6774 7486 6878
rect 7680 6774 7706 6878
rect 10536 6878 10786 7828
rect 7456 6756 7706 6774
rect 8698 6753 8714 6787
rect 8748 6753 8764 6787
rect 9346 6755 9362 6789
rect 9396 6755 9412 6789
rect 8426 6686 8460 6738
rect 3150 6575 3184 6650
rect 3150 6503 3184 6515
rect 3150 6431 3184 6447
rect 3150 6359 3184 6379
rect 3150 6287 3184 6311
rect 3150 6215 3184 6243
rect 3150 6143 3184 6175
rect 3150 6073 3184 6107
rect 3150 6005 3184 6037
rect 3150 5937 3184 5965
rect 3150 5869 3184 5893
rect 3150 5801 3184 5821
rect 3150 5733 3184 5749
rect 3150 5665 3184 5677
rect 3150 5586 3184 5605
rect 3246 6575 3280 6592
rect 3246 6503 3280 6515
rect 3246 6431 3280 6447
rect 3246 6359 3280 6379
rect 3246 6287 3280 6311
rect 3246 6215 3280 6243
rect 3246 6143 3280 6175
rect 3246 6073 3280 6107
rect 3246 6005 3280 6037
rect 3246 5937 3280 5965
rect 3246 5869 3280 5893
rect 3246 5801 3280 5821
rect 3246 5733 3280 5749
rect 3246 5665 3280 5677
rect -868 5419 -834 5453
rect -868 5351 -834 5383
rect 798 5418 996 5516
rect 2056 5514 2666 5548
rect 3246 5534 3280 5605
rect 3342 6575 3376 6650
rect 3342 6503 3376 6515
rect 3342 6431 3376 6447
rect 3342 6359 3376 6379
rect 3342 6287 3376 6311
rect 3342 6215 3376 6243
rect 3342 6143 3376 6175
rect 3342 6073 3376 6107
rect 3342 6005 3376 6037
rect 3342 5937 3376 5965
rect 3342 5869 3376 5893
rect 3342 5801 3376 5821
rect 3342 5733 3376 5749
rect 3342 5665 3376 5677
rect 3342 5588 3376 5605
rect 3438 6575 3472 6592
rect 3438 6503 3472 6515
rect 3438 6431 3472 6447
rect 3438 6359 3472 6379
rect 3438 6287 3472 6311
rect 3438 6215 3472 6243
rect 3438 6143 3472 6175
rect 3438 6073 3472 6107
rect 3438 6005 3472 6037
rect 3438 5937 3472 5965
rect 3438 5869 3472 5893
rect 3438 5801 3472 5821
rect 3438 5733 3472 5749
rect 3438 5665 3472 5677
rect 3438 5534 3472 5605
rect 3534 6575 3568 6650
rect 3534 6503 3568 6515
rect 3534 6431 3568 6447
rect 3534 6359 3568 6379
rect 3534 6287 3568 6311
rect 3534 6215 3568 6243
rect 3534 6143 3568 6175
rect 3534 6073 3568 6107
rect 3534 6005 3568 6037
rect 3534 5937 3568 5965
rect 3534 5869 3568 5893
rect 3534 5801 3568 5821
rect 3534 5733 3568 5749
rect 3534 5665 3568 5677
rect 3534 5588 3568 5605
rect 3630 6575 3664 6592
rect 3630 6503 3664 6515
rect 3630 6431 3664 6447
rect 3630 6359 3664 6379
rect 3630 6287 3664 6311
rect 3630 6215 3664 6243
rect 3630 6143 3664 6175
rect 3630 6073 3664 6107
rect 3630 6005 3664 6037
rect 3630 5937 3664 5965
rect 3630 5869 3664 5893
rect 3630 5801 3664 5821
rect 3630 5733 3664 5749
rect 3630 5665 3664 5677
rect 3630 5534 3664 5605
rect 3726 6575 3760 6650
rect 3726 6503 3760 6515
rect 3726 6431 3760 6447
rect 3726 6359 3760 6379
rect 3726 6287 3760 6311
rect 3726 6215 3760 6243
rect 3726 6143 3760 6175
rect 3726 6073 3760 6107
rect 3726 6005 3760 6037
rect 3726 5937 3760 5965
rect 3726 5869 3760 5893
rect 3726 5801 3760 5821
rect 3726 5733 3760 5749
rect 3726 5665 3760 5677
rect 3726 5588 3760 5605
rect 3822 6575 3856 6592
rect 3822 6503 3856 6515
rect 3822 6431 3856 6447
rect 3822 6359 3856 6379
rect 3822 6287 3856 6311
rect 3822 6215 3856 6243
rect 3822 6143 3856 6175
rect 3822 6073 3856 6107
rect 3822 6005 3856 6037
rect 3822 5937 3856 5965
rect 3822 5869 3856 5893
rect 3822 5801 3856 5821
rect 3822 5733 3856 5749
rect 3822 5665 3856 5677
rect 3822 5534 3856 5605
rect 3918 6575 3952 6650
rect 3918 6503 3952 6515
rect 3918 6431 3952 6447
rect 3918 6359 3952 6379
rect 3918 6287 3952 6311
rect 3918 6215 3952 6243
rect 3918 6143 3952 6175
rect 3918 6073 3952 6107
rect 3918 6005 3952 6037
rect 3918 5937 3952 5965
rect 3918 5869 3952 5893
rect 3918 5801 3952 5821
rect 3918 5733 3952 5749
rect 3918 5665 3952 5677
rect 3918 5588 3952 5605
rect 4014 6575 4048 6592
rect 4014 6503 4048 6515
rect 4014 6431 4048 6447
rect 4014 6359 4048 6379
rect 4014 6287 4048 6311
rect 4014 6215 4048 6243
rect 4014 6143 4048 6175
rect 4014 6073 4048 6107
rect 4014 6005 4048 6037
rect 4014 5937 4048 5965
rect 4014 5869 4048 5893
rect 4014 5801 4048 5821
rect 4014 5733 4048 5749
rect 4014 5665 4048 5677
rect 4014 5534 4048 5605
rect 4110 6575 4144 6650
rect 4110 6503 4144 6515
rect 4110 6431 4144 6447
rect 4110 6359 4144 6379
rect 4110 6287 4144 6311
rect 4110 6215 4144 6243
rect 4110 6143 4144 6175
rect 4110 6073 4144 6107
rect 4110 6005 4144 6037
rect 4110 5937 4144 5965
rect 4110 5869 4144 5893
rect 4110 5801 4144 5821
rect 4110 5733 4144 5749
rect 4110 5665 4144 5677
rect 4110 5588 4144 5605
rect 4206 6575 4240 6592
rect 4206 6503 4240 6515
rect 4206 6431 4240 6447
rect 4206 6359 4240 6379
rect 4206 6287 4240 6311
rect 4206 6215 4240 6243
rect 4206 6143 4240 6175
rect 4206 6073 4240 6107
rect 4206 6005 4240 6037
rect 4206 5937 4240 5965
rect 4206 5869 4240 5893
rect 4206 5801 4240 5821
rect 4206 5733 4240 5749
rect 4206 5665 4240 5677
rect 4206 5534 4240 5605
rect 4302 6575 4336 6650
rect 4302 6503 4336 6515
rect 4302 6431 4336 6447
rect 4302 6359 4336 6379
rect 4302 6287 4336 6311
rect 4302 6215 4336 6243
rect 4302 6143 4336 6175
rect 4302 6073 4336 6107
rect 4302 6005 4336 6037
rect 4302 5937 4336 5965
rect 4302 5869 4336 5893
rect 4302 5801 4336 5821
rect 4302 5733 4336 5749
rect 4302 5665 4336 5677
rect 4302 5588 4336 5605
rect 4916 6571 4950 6652
rect 4916 6499 4950 6511
rect 4916 6427 4950 6443
rect 4916 6355 4950 6375
rect 4916 6283 4950 6307
rect 4916 6211 4950 6239
rect 4916 6139 4950 6171
rect 4916 6069 4950 6103
rect 4916 6001 4950 6033
rect 4916 5933 4950 5961
rect 4916 5865 4950 5889
rect 4916 5797 4950 5817
rect 4916 5729 4950 5745
rect 4916 5661 4950 5673
rect 4916 5582 4950 5601
rect 5012 6571 5046 6588
rect 5012 6499 5046 6511
rect 5012 6427 5046 6443
rect 5012 6355 5046 6375
rect 5012 6283 5046 6307
rect 5012 6211 5046 6239
rect 5012 6139 5046 6171
rect 5012 6069 5046 6103
rect 5012 6001 5046 6033
rect 5012 5933 5046 5961
rect 5012 5865 5046 5889
rect 5012 5797 5046 5817
rect 5012 5729 5046 5745
rect 5012 5661 5046 5673
rect 798 5372 880 5418
rect 982 5372 996 5418
rect 798 5362 996 5372
rect 2266 5418 2464 5514
rect 3246 5500 4240 5534
rect 5012 5532 5046 5601
rect 5108 6571 5142 6652
rect 5108 6499 5142 6511
rect 5108 6427 5142 6443
rect 5108 6355 5142 6375
rect 5108 6283 5142 6307
rect 5108 6211 5142 6239
rect 5108 6139 5142 6171
rect 5108 6069 5142 6103
rect 5108 6001 5142 6033
rect 5108 5933 5142 5961
rect 5108 5865 5142 5889
rect 5108 5797 5142 5817
rect 5108 5729 5142 5745
rect 5108 5661 5142 5673
rect 5108 5582 5142 5601
rect 5204 6571 5238 6588
rect 5204 6499 5238 6511
rect 5204 6427 5238 6443
rect 5204 6355 5238 6375
rect 5204 6283 5238 6307
rect 5204 6211 5238 6239
rect 5204 6139 5238 6171
rect 5204 6069 5238 6103
rect 5204 6001 5238 6033
rect 5204 5933 5238 5961
rect 5204 5865 5238 5889
rect 5204 5797 5238 5817
rect 5204 5729 5238 5745
rect 5204 5661 5238 5673
rect 5204 5532 5238 5601
rect 5300 6571 5334 6652
rect 5300 6499 5334 6511
rect 5300 6427 5334 6443
rect 5300 6355 5334 6375
rect 5300 6283 5334 6307
rect 5300 6211 5334 6239
rect 5300 6139 5334 6171
rect 5300 6069 5334 6103
rect 5300 6001 5334 6033
rect 5300 5933 5334 5961
rect 5300 5865 5334 5889
rect 5300 5797 5334 5817
rect 5300 5729 5334 5745
rect 5300 5661 5334 5673
rect 5300 5582 5334 5601
rect 5396 6571 5430 6588
rect 5396 6499 5430 6511
rect 5396 6427 5430 6443
rect 5396 6355 5430 6375
rect 5396 6283 5430 6307
rect 5396 6211 5430 6239
rect 5396 6139 5430 6171
rect 5396 6069 5430 6103
rect 5396 6001 5430 6033
rect 5396 5933 5430 5961
rect 5396 5865 5430 5889
rect 5396 5797 5430 5817
rect 5396 5729 5430 5745
rect 5396 5661 5430 5673
rect 5396 5532 5430 5601
rect 5492 6571 5526 6652
rect 5492 6499 5526 6511
rect 5492 6427 5526 6443
rect 5492 6355 5526 6375
rect 5492 6283 5526 6307
rect 5492 6211 5526 6239
rect 5492 6139 5526 6171
rect 5492 6069 5526 6103
rect 5492 6001 5526 6033
rect 5492 5933 5526 5961
rect 5492 5865 5526 5889
rect 5492 5797 5526 5817
rect 5492 5729 5526 5745
rect 5492 5661 5526 5673
rect 5492 5582 5526 5601
rect 5588 6571 5622 6588
rect 5588 6499 5622 6511
rect 5588 6427 5622 6443
rect 5588 6355 5622 6375
rect 5588 6283 5622 6307
rect 5588 6211 5622 6239
rect 5588 6139 5622 6171
rect 5588 6069 5622 6103
rect 5588 6001 5622 6033
rect 5588 5933 5622 5961
rect 5588 5865 5622 5889
rect 5588 5797 5622 5817
rect 5588 5729 5622 5745
rect 5588 5661 5622 5673
rect 5588 5532 5622 5601
rect 5684 6571 5718 6652
rect 5684 6499 5718 6511
rect 5684 6427 5718 6443
rect 5684 6355 5718 6375
rect 5684 6283 5718 6307
rect 5684 6211 5718 6239
rect 5684 6139 5718 6171
rect 5684 6069 5718 6103
rect 5684 6001 5718 6033
rect 5684 5933 5718 5961
rect 5684 5865 5718 5889
rect 5684 5797 5718 5817
rect 5684 5729 5718 5745
rect 5684 5661 5718 5673
rect 5684 5584 5718 5601
rect 6180 6650 7374 6684
rect 7946 6652 8754 6686
rect 9838 6682 9872 6840
rect 10536 6774 10568 6878
rect 10762 6774 10786 6878
rect 13692 6852 13942 7828
rect 10536 6758 10786 6774
rect 11786 6751 11802 6785
rect 11836 6751 11852 6785
rect 11514 6684 11548 6736
rect 12502 6729 12518 6763
rect 12552 6729 12568 6763
rect 6180 6575 6214 6650
rect 6180 6503 6214 6515
rect 6180 6431 6214 6447
rect 6180 6359 6214 6379
rect 6180 6287 6214 6311
rect 6180 6215 6214 6243
rect 6180 6143 6214 6175
rect 6180 6073 6214 6107
rect 6180 6005 6214 6037
rect 6180 5937 6214 5965
rect 6180 5869 6214 5893
rect 6180 5801 6214 5821
rect 6180 5733 6214 5749
rect 6180 5665 6214 5677
rect 6180 5586 6214 5605
rect 6276 6575 6310 6592
rect 6276 6503 6310 6515
rect 6276 6431 6310 6447
rect 6276 6359 6310 6379
rect 6276 6287 6310 6311
rect 6276 6215 6310 6243
rect 6276 6143 6310 6175
rect 6276 6073 6310 6107
rect 6276 6005 6310 6037
rect 6276 5937 6310 5965
rect 6276 5869 6310 5893
rect 6276 5801 6310 5821
rect 6276 5733 6310 5749
rect 6276 5665 6310 5677
rect 2266 5372 2278 5418
rect 2380 5372 2464 5418
rect 2266 5354 2464 5372
rect 3748 5400 3946 5500
rect 5012 5498 5622 5532
rect 6276 5534 6310 5605
rect 6372 6575 6406 6650
rect 6372 6503 6406 6515
rect 6372 6431 6406 6447
rect 6372 6359 6406 6379
rect 6372 6287 6406 6311
rect 6372 6215 6406 6243
rect 6372 6143 6406 6175
rect 6372 6073 6406 6107
rect 6372 6005 6406 6037
rect 6372 5937 6406 5965
rect 6372 5869 6406 5893
rect 6372 5801 6406 5821
rect 6372 5733 6406 5749
rect 6372 5665 6406 5677
rect 6372 5588 6406 5605
rect 6468 6575 6502 6592
rect 6468 6503 6502 6515
rect 6468 6431 6502 6447
rect 6468 6359 6502 6379
rect 6468 6287 6502 6311
rect 6468 6215 6502 6243
rect 6468 6143 6502 6175
rect 6468 6073 6502 6107
rect 6468 6005 6502 6037
rect 6468 5937 6502 5965
rect 6468 5869 6502 5893
rect 6468 5801 6502 5821
rect 6468 5733 6502 5749
rect 6468 5665 6502 5677
rect 6468 5534 6502 5605
rect 6564 6575 6598 6650
rect 6564 6503 6598 6515
rect 6564 6431 6598 6447
rect 6564 6359 6598 6379
rect 6564 6287 6598 6311
rect 6564 6215 6598 6243
rect 6564 6143 6598 6175
rect 6564 6073 6598 6107
rect 6564 6005 6598 6037
rect 6564 5937 6598 5965
rect 6564 5869 6598 5893
rect 6564 5801 6598 5821
rect 6564 5733 6598 5749
rect 6564 5665 6598 5677
rect 6564 5588 6598 5605
rect 6660 6575 6694 6592
rect 6660 6503 6694 6515
rect 6660 6431 6694 6447
rect 6660 6359 6694 6379
rect 6660 6287 6694 6311
rect 6660 6215 6694 6243
rect 6660 6143 6694 6175
rect 6660 6073 6694 6107
rect 6660 6005 6694 6037
rect 6660 5937 6694 5965
rect 6660 5869 6694 5893
rect 6660 5801 6694 5821
rect 6660 5733 6694 5749
rect 6660 5665 6694 5677
rect 6660 5534 6694 5605
rect 6756 6575 6790 6650
rect 6756 6503 6790 6515
rect 6756 6431 6790 6447
rect 6756 6359 6790 6379
rect 6756 6287 6790 6311
rect 6756 6215 6790 6243
rect 6756 6143 6790 6175
rect 6756 6073 6790 6107
rect 6756 6005 6790 6037
rect 6756 5937 6790 5965
rect 6756 5869 6790 5893
rect 6756 5801 6790 5821
rect 6756 5733 6790 5749
rect 6756 5665 6790 5677
rect 6756 5588 6790 5605
rect 6852 6575 6886 6592
rect 6852 6503 6886 6515
rect 6852 6431 6886 6447
rect 6852 6359 6886 6379
rect 6852 6287 6886 6311
rect 6852 6215 6886 6243
rect 6852 6143 6886 6175
rect 6852 6073 6886 6107
rect 6852 6005 6886 6037
rect 6852 5937 6886 5965
rect 6852 5869 6886 5893
rect 6852 5801 6886 5821
rect 6852 5733 6886 5749
rect 6852 5665 6886 5677
rect 6852 5534 6886 5605
rect 6948 6575 6982 6650
rect 6948 6503 6982 6515
rect 6948 6431 6982 6447
rect 6948 6359 6982 6379
rect 6948 6287 6982 6311
rect 6948 6215 6982 6243
rect 6948 6143 6982 6175
rect 6948 6073 6982 6107
rect 6948 6005 6982 6037
rect 6948 5937 6982 5965
rect 6948 5869 6982 5893
rect 6948 5801 6982 5821
rect 6948 5733 6982 5749
rect 6948 5665 6982 5677
rect 6948 5588 6982 5605
rect 7044 6575 7078 6592
rect 7044 6503 7078 6515
rect 7044 6431 7078 6447
rect 7044 6359 7078 6379
rect 7044 6287 7078 6311
rect 7044 6215 7078 6243
rect 7044 6143 7078 6175
rect 7044 6073 7078 6107
rect 7044 6005 7078 6037
rect 7044 5937 7078 5965
rect 7044 5869 7078 5893
rect 7044 5801 7078 5821
rect 7044 5733 7078 5749
rect 7044 5665 7078 5677
rect 7044 5534 7078 5605
rect 7140 6575 7174 6650
rect 7140 6503 7174 6515
rect 7140 6431 7174 6447
rect 7140 6359 7174 6379
rect 7140 6287 7174 6311
rect 7140 6215 7174 6243
rect 7140 6143 7174 6175
rect 7140 6073 7174 6107
rect 7140 6005 7174 6037
rect 7140 5937 7174 5965
rect 7140 5869 7174 5893
rect 7140 5801 7174 5821
rect 7140 5733 7174 5749
rect 7140 5665 7174 5677
rect 7140 5588 7174 5605
rect 7236 6575 7270 6592
rect 7236 6503 7270 6515
rect 7236 6431 7270 6447
rect 7236 6359 7270 6379
rect 7236 6287 7270 6311
rect 7236 6215 7270 6243
rect 7236 6143 7270 6175
rect 7236 6073 7270 6107
rect 7236 6005 7270 6037
rect 7236 5937 7270 5965
rect 7236 5869 7270 5893
rect 7236 5801 7270 5821
rect 7236 5733 7270 5749
rect 7236 5665 7270 5677
rect 7236 5534 7270 5605
rect 7332 6575 7366 6650
rect 7332 6503 7366 6515
rect 7332 6431 7366 6447
rect 7332 6359 7366 6379
rect 7332 6287 7366 6311
rect 7332 6215 7366 6243
rect 7332 6143 7366 6175
rect 7332 6073 7366 6107
rect 7332 6005 7366 6037
rect 7332 5937 7366 5965
rect 7332 5869 7366 5893
rect 7332 5801 7366 5821
rect 7332 5733 7366 5749
rect 7332 5665 7366 5677
rect 7332 5588 7366 5605
rect 7946 6571 7980 6652
rect 7946 6499 7980 6511
rect 7946 6427 7980 6443
rect 7946 6355 7980 6375
rect 7946 6283 7980 6307
rect 7946 6211 7980 6239
rect 7946 6139 7980 6171
rect 7946 6069 7980 6103
rect 7946 6001 7980 6033
rect 7946 5933 7980 5961
rect 7946 5865 7980 5889
rect 7946 5797 7980 5817
rect 7946 5729 7980 5745
rect 7946 5661 7980 5673
rect 7946 5582 7980 5601
rect 8042 6571 8076 6588
rect 8042 6499 8076 6511
rect 8042 6427 8076 6443
rect 8042 6355 8076 6375
rect 8042 6283 8076 6307
rect 8042 6211 8076 6239
rect 8042 6139 8076 6171
rect 8042 6069 8076 6103
rect 8042 6001 8076 6033
rect 8042 5933 8076 5961
rect 8042 5865 8076 5889
rect 8042 5797 8076 5817
rect 8042 5729 8076 5745
rect 8042 5661 8076 5673
rect 6276 5500 7270 5534
rect 8042 5532 8076 5601
rect 8138 6571 8172 6652
rect 8138 6499 8172 6511
rect 8138 6427 8172 6443
rect 8138 6355 8172 6375
rect 8138 6283 8172 6307
rect 8138 6211 8172 6239
rect 8138 6139 8172 6171
rect 8138 6069 8172 6103
rect 8138 6001 8172 6033
rect 8138 5933 8172 5961
rect 8138 5865 8172 5889
rect 8138 5797 8172 5817
rect 8138 5729 8172 5745
rect 8138 5661 8172 5673
rect 8138 5582 8172 5601
rect 8234 6571 8268 6588
rect 8234 6499 8268 6511
rect 8234 6427 8268 6443
rect 8234 6355 8268 6375
rect 8234 6283 8268 6307
rect 8234 6211 8268 6239
rect 8234 6139 8268 6171
rect 8234 6069 8268 6103
rect 8234 6001 8268 6033
rect 8234 5933 8268 5961
rect 8234 5865 8268 5889
rect 8234 5797 8268 5817
rect 8234 5729 8268 5745
rect 8234 5661 8268 5673
rect 8234 5532 8268 5601
rect 8330 6571 8364 6652
rect 8330 6499 8364 6511
rect 8330 6427 8364 6443
rect 8330 6355 8364 6375
rect 8330 6283 8364 6307
rect 8330 6211 8364 6239
rect 8330 6139 8364 6171
rect 8330 6069 8364 6103
rect 8330 6001 8364 6033
rect 8330 5933 8364 5961
rect 8330 5865 8364 5889
rect 8330 5797 8364 5817
rect 8330 5729 8364 5745
rect 8330 5661 8364 5673
rect 8330 5582 8364 5601
rect 8426 6571 8460 6588
rect 8426 6499 8460 6511
rect 8426 6427 8460 6443
rect 8426 6355 8460 6375
rect 8426 6283 8460 6307
rect 8426 6211 8460 6239
rect 8426 6139 8460 6171
rect 8426 6069 8460 6103
rect 8426 6001 8460 6033
rect 8426 5933 8460 5961
rect 8426 5865 8460 5889
rect 8426 5797 8460 5817
rect 8426 5729 8460 5745
rect 8426 5661 8460 5673
rect 8426 5532 8460 5601
rect 8522 6571 8556 6652
rect 8522 6499 8556 6511
rect 8522 6427 8556 6443
rect 8522 6355 8556 6375
rect 8522 6283 8556 6307
rect 8522 6211 8556 6239
rect 8522 6139 8556 6171
rect 8522 6069 8556 6103
rect 8522 6001 8556 6033
rect 8522 5933 8556 5961
rect 8522 5865 8556 5889
rect 8522 5797 8556 5817
rect 8522 5729 8556 5745
rect 8522 5661 8556 5673
rect 8522 5582 8556 5601
rect 8618 6571 8652 6588
rect 8618 6499 8652 6511
rect 8618 6427 8652 6443
rect 8618 6355 8652 6375
rect 8618 6283 8652 6307
rect 8618 6211 8652 6239
rect 8618 6139 8652 6171
rect 8618 6069 8652 6103
rect 8618 6001 8652 6033
rect 8618 5933 8652 5961
rect 8618 5865 8652 5889
rect 8618 5797 8652 5817
rect 8618 5729 8652 5745
rect 8618 5661 8652 5673
rect 8618 5532 8652 5601
rect 8714 6571 8748 6652
rect 8714 6499 8748 6511
rect 8714 6427 8748 6443
rect 8714 6355 8748 6375
rect 8714 6283 8748 6307
rect 8714 6211 8748 6239
rect 8714 6139 8748 6171
rect 8714 6069 8748 6103
rect 8714 6001 8748 6033
rect 8714 5933 8748 5961
rect 8714 5865 8748 5889
rect 8714 5797 8748 5817
rect 8714 5729 8748 5745
rect 8714 5661 8748 5673
rect 8714 5584 8748 5601
rect 9268 6648 10462 6682
rect 11034 6650 11842 6684
rect 12994 6656 13028 6814
rect 13692 6748 13724 6852
rect 13918 6748 13942 6852
rect 13692 6732 13942 6748
rect 14942 6725 14958 6759
rect 14992 6725 15008 6759
rect 14670 6658 14704 6710
rect 9268 6573 9302 6648
rect 9268 6501 9302 6513
rect 9268 6429 9302 6445
rect 9268 6357 9302 6377
rect 9268 6285 9302 6309
rect 9268 6213 9302 6241
rect 9268 6141 9302 6173
rect 9268 6071 9302 6105
rect 9268 6003 9302 6035
rect 9268 5935 9302 5963
rect 9268 5867 9302 5891
rect 9268 5799 9302 5819
rect 9268 5731 9302 5747
rect 9268 5663 9302 5675
rect 9268 5584 9302 5603
rect 9364 6573 9398 6590
rect 9364 6501 9398 6513
rect 9364 6429 9398 6445
rect 9364 6357 9398 6377
rect 9364 6285 9398 6309
rect 9364 6213 9398 6241
rect 9364 6141 9398 6173
rect 9364 6071 9398 6105
rect 9364 6003 9398 6035
rect 9364 5935 9398 5963
rect 9364 5867 9398 5891
rect 9364 5799 9398 5819
rect 9364 5731 9398 5747
rect 9364 5663 9398 5675
rect 3748 5354 3824 5400
rect 3926 5354 3946 5400
rect 3748 5338 3946 5354
rect 5214 5398 5412 5498
rect 5214 5352 5234 5398
rect 5336 5352 5412 5398
rect 5214 5332 5412 5352
rect 6780 5398 6978 5500
rect 8042 5498 8652 5532
rect 9364 5532 9398 5603
rect 9460 6573 9494 6648
rect 9460 6501 9494 6513
rect 9460 6429 9494 6445
rect 9460 6357 9494 6377
rect 9460 6285 9494 6309
rect 9460 6213 9494 6241
rect 9460 6141 9494 6173
rect 9460 6071 9494 6105
rect 9460 6003 9494 6035
rect 9460 5935 9494 5963
rect 9460 5867 9494 5891
rect 9460 5799 9494 5819
rect 9460 5731 9494 5747
rect 9460 5663 9494 5675
rect 9460 5586 9494 5603
rect 9556 6573 9590 6590
rect 9556 6501 9590 6513
rect 9556 6429 9590 6445
rect 9556 6357 9590 6377
rect 9556 6285 9590 6309
rect 9556 6213 9590 6241
rect 9556 6141 9590 6173
rect 9556 6071 9590 6105
rect 9556 6003 9590 6035
rect 9556 5935 9590 5963
rect 9556 5867 9590 5891
rect 9556 5799 9590 5819
rect 9556 5731 9590 5747
rect 9556 5663 9590 5675
rect 9556 5532 9590 5603
rect 9652 6573 9686 6648
rect 9652 6501 9686 6513
rect 9652 6429 9686 6445
rect 9652 6357 9686 6377
rect 9652 6285 9686 6309
rect 9652 6213 9686 6241
rect 9652 6141 9686 6173
rect 9652 6071 9686 6105
rect 9652 6003 9686 6035
rect 9652 5935 9686 5963
rect 9652 5867 9686 5891
rect 9652 5799 9686 5819
rect 9652 5731 9686 5747
rect 9652 5663 9686 5675
rect 9652 5586 9686 5603
rect 9748 6573 9782 6590
rect 9748 6501 9782 6513
rect 9748 6429 9782 6445
rect 9748 6357 9782 6377
rect 9748 6285 9782 6309
rect 9748 6213 9782 6241
rect 9748 6141 9782 6173
rect 9748 6071 9782 6105
rect 9748 6003 9782 6035
rect 9748 5935 9782 5963
rect 9748 5867 9782 5891
rect 9748 5799 9782 5819
rect 9748 5731 9782 5747
rect 9748 5663 9782 5675
rect 9748 5532 9782 5603
rect 9844 6573 9878 6648
rect 9844 6501 9878 6513
rect 9844 6429 9878 6445
rect 9844 6357 9878 6377
rect 9844 6285 9878 6309
rect 9844 6213 9878 6241
rect 9844 6141 9878 6173
rect 9844 6071 9878 6105
rect 9844 6003 9878 6035
rect 9844 5935 9878 5963
rect 9844 5867 9878 5891
rect 9844 5799 9878 5819
rect 9844 5731 9878 5747
rect 9844 5663 9878 5675
rect 9844 5586 9878 5603
rect 9940 6573 9974 6590
rect 9940 6501 9974 6513
rect 9940 6429 9974 6445
rect 9940 6357 9974 6377
rect 9940 6285 9974 6309
rect 9940 6213 9974 6241
rect 9940 6141 9974 6173
rect 9940 6071 9974 6105
rect 9940 6003 9974 6035
rect 9940 5935 9974 5963
rect 9940 5867 9974 5891
rect 9940 5799 9974 5819
rect 9940 5731 9974 5747
rect 9940 5663 9974 5675
rect 9940 5532 9974 5603
rect 10036 6573 10070 6648
rect 10036 6501 10070 6513
rect 10036 6429 10070 6445
rect 10036 6357 10070 6377
rect 10036 6285 10070 6309
rect 10036 6213 10070 6241
rect 10036 6141 10070 6173
rect 10036 6071 10070 6105
rect 10036 6003 10070 6035
rect 10036 5935 10070 5963
rect 10036 5867 10070 5891
rect 10036 5799 10070 5819
rect 10036 5731 10070 5747
rect 10036 5663 10070 5675
rect 10036 5586 10070 5603
rect 10132 6573 10166 6590
rect 10132 6501 10166 6513
rect 10132 6429 10166 6445
rect 10132 6357 10166 6377
rect 10132 6285 10166 6309
rect 10132 6213 10166 6241
rect 10132 6141 10166 6173
rect 10132 6071 10166 6105
rect 10132 6003 10166 6035
rect 10132 5935 10166 5963
rect 10132 5867 10166 5891
rect 10132 5799 10166 5819
rect 10132 5731 10166 5747
rect 10132 5663 10166 5675
rect 10132 5532 10166 5603
rect 10228 6573 10262 6648
rect 10228 6501 10262 6513
rect 10228 6429 10262 6445
rect 10228 6357 10262 6377
rect 10228 6285 10262 6309
rect 10228 6213 10262 6241
rect 10228 6141 10262 6173
rect 10228 6071 10262 6105
rect 10228 6003 10262 6035
rect 10228 5935 10262 5963
rect 10228 5867 10262 5891
rect 10228 5799 10262 5819
rect 10228 5731 10262 5747
rect 10228 5663 10262 5675
rect 10228 5586 10262 5603
rect 10324 6573 10358 6590
rect 10324 6501 10358 6513
rect 10324 6429 10358 6445
rect 10324 6357 10358 6377
rect 10324 6285 10358 6309
rect 10324 6213 10358 6241
rect 10324 6141 10358 6173
rect 10324 6071 10358 6105
rect 10324 6003 10358 6035
rect 10324 5935 10358 5963
rect 10324 5867 10358 5891
rect 10324 5799 10358 5819
rect 10324 5731 10358 5747
rect 10324 5663 10358 5675
rect 10324 5532 10358 5603
rect 10420 6573 10454 6648
rect 10420 6501 10454 6513
rect 10420 6429 10454 6445
rect 10420 6357 10454 6377
rect 10420 6285 10454 6309
rect 10420 6213 10454 6241
rect 10420 6141 10454 6173
rect 10420 6071 10454 6105
rect 10420 6003 10454 6035
rect 10420 5935 10454 5963
rect 10420 5867 10454 5891
rect 10420 5799 10454 5819
rect 10420 5731 10454 5747
rect 10420 5663 10454 5675
rect 10420 5586 10454 5603
rect 11034 6569 11068 6650
rect 11034 6497 11068 6509
rect 11034 6425 11068 6441
rect 11034 6353 11068 6373
rect 11034 6281 11068 6305
rect 11034 6209 11068 6237
rect 11034 6137 11068 6169
rect 11034 6067 11068 6101
rect 11034 5999 11068 6031
rect 11034 5931 11068 5959
rect 11034 5863 11068 5887
rect 11034 5795 11068 5815
rect 11034 5727 11068 5743
rect 11034 5659 11068 5671
rect 11034 5580 11068 5599
rect 11130 6569 11164 6586
rect 11130 6497 11164 6509
rect 11130 6425 11164 6441
rect 11130 6353 11164 6373
rect 11130 6281 11164 6305
rect 11130 6209 11164 6237
rect 11130 6137 11164 6169
rect 11130 6067 11164 6101
rect 11130 5999 11164 6031
rect 11130 5931 11164 5959
rect 11130 5863 11164 5887
rect 11130 5795 11164 5815
rect 11130 5727 11164 5743
rect 11130 5659 11164 5671
rect 9364 5498 10358 5532
rect 11130 5530 11164 5599
rect 11226 6569 11260 6650
rect 11226 6497 11260 6509
rect 11226 6425 11260 6441
rect 11226 6353 11260 6373
rect 11226 6281 11260 6305
rect 11226 6209 11260 6237
rect 11226 6137 11260 6169
rect 11226 6067 11260 6101
rect 11226 5999 11260 6031
rect 11226 5931 11260 5959
rect 11226 5863 11260 5887
rect 11226 5795 11260 5815
rect 11226 5727 11260 5743
rect 11226 5659 11260 5671
rect 11226 5580 11260 5599
rect 11322 6569 11356 6586
rect 11322 6497 11356 6509
rect 11322 6425 11356 6441
rect 11322 6353 11356 6373
rect 11322 6281 11356 6305
rect 11322 6209 11356 6237
rect 11322 6137 11356 6169
rect 11322 6067 11356 6101
rect 11322 5999 11356 6031
rect 11322 5931 11356 5959
rect 11322 5863 11356 5887
rect 11322 5795 11356 5815
rect 11322 5727 11356 5743
rect 11322 5659 11356 5671
rect 11322 5530 11356 5599
rect 11418 6569 11452 6650
rect 11418 6497 11452 6509
rect 11418 6425 11452 6441
rect 11418 6353 11452 6373
rect 11418 6281 11452 6305
rect 11418 6209 11452 6237
rect 11418 6137 11452 6169
rect 11418 6067 11452 6101
rect 11418 5999 11452 6031
rect 11418 5931 11452 5959
rect 11418 5863 11452 5887
rect 11418 5795 11452 5815
rect 11418 5727 11452 5743
rect 11418 5659 11452 5671
rect 11418 5580 11452 5599
rect 11514 6569 11548 6586
rect 11514 6497 11548 6509
rect 11514 6425 11548 6441
rect 11514 6353 11548 6373
rect 11514 6281 11548 6305
rect 11514 6209 11548 6237
rect 11514 6137 11548 6169
rect 11514 6067 11548 6101
rect 11514 5999 11548 6031
rect 11514 5931 11548 5959
rect 11514 5863 11548 5887
rect 11514 5795 11548 5815
rect 11514 5727 11548 5743
rect 11514 5659 11548 5671
rect 11514 5530 11548 5599
rect 11610 6569 11644 6650
rect 11610 6497 11644 6509
rect 11610 6425 11644 6441
rect 11610 6353 11644 6373
rect 11610 6281 11644 6305
rect 11610 6209 11644 6237
rect 11610 6137 11644 6169
rect 11610 6067 11644 6101
rect 11610 5999 11644 6031
rect 11610 5931 11644 5959
rect 11610 5863 11644 5887
rect 11610 5795 11644 5815
rect 11610 5727 11644 5743
rect 11610 5659 11644 5671
rect 11610 5580 11644 5599
rect 11706 6569 11740 6586
rect 11706 6497 11740 6509
rect 11706 6425 11740 6441
rect 11706 6353 11740 6373
rect 11706 6281 11740 6305
rect 11706 6209 11740 6237
rect 11706 6137 11740 6169
rect 11706 6067 11740 6101
rect 11706 5999 11740 6031
rect 11706 5931 11740 5959
rect 11706 5863 11740 5887
rect 11706 5795 11740 5815
rect 11706 5727 11740 5743
rect 11706 5659 11740 5671
rect 11706 5530 11740 5599
rect 11802 6569 11836 6650
rect 11802 6497 11836 6509
rect 11802 6425 11836 6441
rect 11802 6353 11836 6373
rect 11802 6281 11836 6305
rect 11802 6209 11836 6237
rect 11802 6137 11836 6169
rect 11802 6067 11836 6101
rect 11802 5999 11836 6031
rect 11802 5931 11836 5959
rect 11802 5863 11836 5887
rect 11802 5795 11836 5815
rect 11802 5727 11836 5743
rect 11802 5659 11836 5671
rect 11802 5582 11836 5599
rect 12424 6622 13618 6656
rect 14190 6624 14998 6658
rect 12424 6547 12458 6622
rect 12424 6475 12458 6487
rect 12424 6403 12458 6419
rect 12424 6331 12458 6351
rect 12424 6259 12458 6283
rect 12424 6187 12458 6215
rect 12424 6115 12458 6147
rect 12424 6045 12458 6079
rect 12424 5977 12458 6009
rect 12424 5909 12458 5937
rect 12424 5841 12458 5865
rect 12424 5773 12458 5793
rect 12424 5705 12458 5721
rect 12424 5637 12458 5649
rect 12424 5558 12458 5577
rect 12520 6547 12554 6564
rect 12520 6475 12554 6487
rect 12520 6403 12554 6419
rect 12520 6331 12554 6351
rect 12520 6259 12554 6283
rect 12520 6187 12554 6215
rect 12520 6115 12554 6147
rect 12520 6045 12554 6079
rect 12520 5977 12554 6009
rect 12520 5909 12554 5937
rect 12520 5841 12554 5865
rect 12520 5773 12554 5793
rect 12520 5705 12554 5721
rect 12520 5637 12554 5649
rect 6780 5352 6854 5398
rect 6956 5352 6978 5398
rect 6780 5334 6978 5352
rect 8246 5402 8444 5498
rect 8246 5356 8268 5402
rect 8370 5356 8444 5402
rect 8246 5332 8444 5356
rect 9872 5392 10070 5498
rect 11130 5496 11740 5530
rect 12520 5506 12554 5577
rect 12616 6547 12650 6622
rect 12616 6475 12650 6487
rect 12616 6403 12650 6419
rect 12616 6331 12650 6351
rect 12616 6259 12650 6283
rect 12616 6187 12650 6215
rect 12616 6115 12650 6147
rect 12616 6045 12650 6079
rect 12616 5977 12650 6009
rect 12616 5909 12650 5937
rect 12616 5841 12650 5865
rect 12616 5773 12650 5793
rect 12616 5705 12650 5721
rect 12616 5637 12650 5649
rect 12616 5560 12650 5577
rect 12712 6547 12746 6564
rect 12712 6475 12746 6487
rect 12712 6403 12746 6419
rect 12712 6331 12746 6351
rect 12712 6259 12746 6283
rect 12712 6187 12746 6215
rect 12712 6115 12746 6147
rect 12712 6045 12746 6079
rect 12712 5977 12746 6009
rect 12712 5909 12746 5937
rect 12712 5841 12746 5865
rect 12712 5773 12746 5793
rect 12712 5705 12746 5721
rect 12712 5637 12746 5649
rect 12712 5506 12746 5577
rect 12808 6547 12842 6622
rect 12808 6475 12842 6487
rect 12808 6403 12842 6419
rect 12808 6331 12842 6351
rect 12808 6259 12842 6283
rect 12808 6187 12842 6215
rect 12808 6115 12842 6147
rect 12808 6045 12842 6079
rect 12808 5977 12842 6009
rect 12808 5909 12842 5937
rect 12808 5841 12842 5865
rect 12808 5773 12842 5793
rect 12808 5705 12842 5721
rect 12808 5637 12842 5649
rect 12808 5560 12842 5577
rect 12904 6547 12938 6564
rect 12904 6475 12938 6487
rect 12904 6403 12938 6419
rect 12904 6331 12938 6351
rect 12904 6259 12938 6283
rect 12904 6187 12938 6215
rect 12904 6115 12938 6147
rect 12904 6045 12938 6079
rect 12904 5977 12938 6009
rect 12904 5909 12938 5937
rect 12904 5841 12938 5865
rect 12904 5773 12938 5793
rect 12904 5705 12938 5721
rect 12904 5637 12938 5649
rect 12904 5506 12938 5577
rect 13000 6547 13034 6622
rect 13000 6475 13034 6487
rect 13000 6403 13034 6419
rect 13000 6331 13034 6351
rect 13000 6259 13034 6283
rect 13000 6187 13034 6215
rect 13000 6115 13034 6147
rect 13000 6045 13034 6079
rect 13000 5977 13034 6009
rect 13000 5909 13034 5937
rect 13000 5841 13034 5865
rect 13000 5773 13034 5793
rect 13000 5705 13034 5721
rect 13000 5637 13034 5649
rect 13000 5560 13034 5577
rect 13096 6547 13130 6564
rect 13096 6475 13130 6487
rect 13096 6403 13130 6419
rect 13096 6331 13130 6351
rect 13096 6259 13130 6283
rect 13096 6187 13130 6215
rect 13096 6115 13130 6147
rect 13096 6045 13130 6079
rect 13096 5977 13130 6009
rect 13096 5909 13130 5937
rect 13096 5841 13130 5865
rect 13096 5773 13130 5793
rect 13096 5705 13130 5721
rect 13096 5637 13130 5649
rect 13096 5506 13130 5577
rect 13192 6547 13226 6622
rect 13192 6475 13226 6487
rect 13192 6403 13226 6419
rect 13192 6331 13226 6351
rect 13192 6259 13226 6283
rect 13192 6187 13226 6215
rect 13192 6115 13226 6147
rect 13192 6045 13226 6079
rect 13192 5977 13226 6009
rect 13192 5909 13226 5937
rect 13192 5841 13226 5865
rect 13192 5773 13226 5793
rect 13192 5705 13226 5721
rect 13192 5637 13226 5649
rect 13192 5560 13226 5577
rect 13288 6547 13322 6564
rect 13288 6475 13322 6487
rect 13288 6403 13322 6419
rect 13288 6331 13322 6351
rect 13288 6259 13322 6283
rect 13288 6187 13322 6215
rect 13288 6115 13322 6147
rect 13288 6045 13322 6079
rect 13288 5977 13322 6009
rect 13288 5909 13322 5937
rect 13288 5841 13322 5865
rect 13288 5773 13322 5793
rect 13288 5705 13322 5721
rect 13288 5637 13322 5649
rect 13288 5506 13322 5577
rect 13384 6547 13418 6622
rect 13384 6475 13418 6487
rect 13384 6403 13418 6419
rect 13384 6331 13418 6351
rect 13384 6259 13418 6283
rect 13384 6187 13418 6215
rect 13384 6115 13418 6147
rect 13384 6045 13418 6079
rect 13384 5977 13418 6009
rect 13384 5909 13418 5937
rect 13384 5841 13418 5865
rect 13384 5773 13418 5793
rect 13384 5705 13418 5721
rect 13384 5637 13418 5649
rect 13384 5560 13418 5577
rect 13480 6547 13514 6564
rect 13480 6475 13514 6487
rect 13480 6403 13514 6419
rect 13480 6331 13514 6351
rect 13480 6259 13514 6283
rect 13480 6187 13514 6215
rect 13480 6115 13514 6147
rect 13480 6045 13514 6079
rect 13480 5977 13514 6009
rect 13480 5909 13514 5937
rect 13480 5841 13514 5865
rect 13480 5773 13514 5793
rect 13480 5705 13514 5721
rect 13480 5637 13514 5649
rect 13480 5506 13514 5577
rect 13576 6547 13610 6622
rect 13576 6475 13610 6487
rect 13576 6403 13610 6419
rect 13576 6331 13610 6351
rect 13576 6259 13610 6283
rect 13576 6187 13610 6215
rect 13576 6115 13610 6147
rect 13576 6045 13610 6079
rect 13576 5977 13610 6009
rect 13576 5909 13610 5937
rect 13576 5841 13610 5865
rect 13576 5773 13610 5793
rect 13576 5705 13610 5721
rect 13576 5637 13610 5649
rect 13576 5560 13610 5577
rect 14190 6543 14224 6624
rect 14190 6471 14224 6483
rect 14190 6399 14224 6415
rect 14190 6327 14224 6347
rect 14190 6255 14224 6279
rect 14190 6183 14224 6211
rect 14190 6111 14224 6143
rect 14190 6041 14224 6075
rect 14190 5973 14224 6005
rect 14190 5905 14224 5933
rect 14190 5837 14224 5861
rect 14190 5769 14224 5789
rect 14190 5701 14224 5717
rect 14190 5633 14224 5645
rect 14190 5554 14224 5573
rect 14286 6543 14320 6560
rect 14286 6471 14320 6483
rect 14286 6399 14320 6415
rect 14286 6327 14320 6347
rect 14286 6255 14320 6279
rect 14286 6183 14320 6211
rect 14286 6111 14320 6143
rect 14286 6041 14320 6075
rect 14286 5973 14320 6005
rect 14286 5905 14320 5933
rect 14286 5837 14320 5861
rect 14286 5769 14320 5789
rect 14286 5701 14320 5717
rect 14286 5633 14320 5645
rect 9872 5346 9950 5392
rect 10052 5346 10070 5392
rect 9872 5332 10070 5346
rect 11334 5398 11532 5496
rect 12520 5472 13514 5506
rect 14286 5504 14320 5573
rect 14382 6543 14416 6624
rect 14382 6471 14416 6483
rect 14382 6399 14416 6415
rect 14382 6327 14416 6347
rect 14382 6255 14416 6279
rect 14382 6183 14416 6211
rect 14382 6111 14416 6143
rect 14382 6041 14416 6075
rect 14382 5973 14416 6005
rect 14382 5905 14416 5933
rect 14382 5837 14416 5861
rect 14382 5769 14416 5789
rect 14382 5701 14416 5717
rect 14382 5633 14416 5645
rect 14382 5554 14416 5573
rect 14478 6543 14512 6560
rect 14478 6471 14512 6483
rect 14478 6399 14512 6415
rect 14478 6327 14512 6347
rect 14478 6255 14512 6279
rect 14478 6183 14512 6211
rect 14478 6111 14512 6143
rect 14478 6041 14512 6075
rect 14478 5973 14512 6005
rect 14478 5905 14512 5933
rect 14478 5837 14512 5861
rect 14478 5769 14512 5789
rect 14478 5701 14512 5717
rect 14478 5633 14512 5645
rect 14478 5504 14512 5573
rect 14574 6543 14608 6624
rect 14574 6471 14608 6483
rect 14574 6399 14608 6415
rect 14574 6327 14608 6347
rect 14574 6255 14608 6279
rect 14574 6183 14608 6211
rect 14574 6111 14608 6143
rect 14574 6041 14608 6075
rect 14574 5973 14608 6005
rect 14574 5905 14608 5933
rect 14574 5837 14608 5861
rect 14574 5769 14608 5789
rect 14574 5701 14608 5717
rect 14574 5633 14608 5645
rect 14574 5554 14608 5573
rect 14670 6543 14704 6560
rect 14670 6471 14704 6483
rect 14670 6399 14704 6415
rect 14670 6327 14704 6347
rect 14670 6255 14704 6279
rect 14670 6183 14704 6211
rect 14670 6111 14704 6143
rect 14670 6041 14704 6075
rect 14670 5973 14704 6005
rect 14670 5905 14704 5933
rect 14670 5837 14704 5861
rect 14670 5769 14704 5789
rect 14670 5701 14704 5717
rect 14670 5633 14704 5645
rect 14670 5504 14704 5573
rect 14766 6543 14800 6624
rect 14766 6471 14800 6483
rect 14766 6399 14800 6415
rect 14766 6327 14800 6347
rect 14766 6255 14800 6279
rect 14766 6183 14800 6211
rect 14766 6111 14800 6143
rect 14766 6041 14800 6075
rect 14766 5973 14800 6005
rect 14766 5905 14800 5933
rect 14766 5837 14800 5861
rect 14766 5769 14800 5789
rect 14766 5701 14800 5717
rect 14766 5633 14800 5645
rect 14766 5554 14800 5573
rect 14862 6543 14896 6560
rect 14862 6471 14896 6483
rect 14862 6399 14896 6415
rect 14862 6327 14896 6347
rect 14862 6255 14896 6279
rect 14862 6183 14896 6211
rect 14862 6111 14896 6143
rect 14862 6041 14896 6075
rect 14862 5973 14896 6005
rect 14862 5905 14896 5933
rect 14862 5837 14896 5861
rect 14862 5769 14896 5789
rect 14862 5701 14896 5717
rect 14862 5633 14896 5645
rect 14862 5504 14896 5573
rect 14958 6543 14992 6624
rect 14958 6471 14992 6483
rect 14958 6399 14992 6415
rect 14958 6327 14992 6347
rect 14958 6255 14992 6279
rect 14958 6183 14992 6211
rect 14958 6111 14992 6143
rect 14958 6041 14992 6075
rect 15614 6032 15648 6148
rect 14958 5973 14992 6005
rect 14958 5905 14992 5933
rect 14958 5837 14992 5861
rect 14958 5769 14992 5789
rect 14958 5701 14992 5717
rect 14958 5633 14992 5645
rect 14958 5556 14992 5573
rect 15518 5996 15744 6032
rect 15518 5895 15552 5996
rect 15518 5827 15552 5845
rect 15518 5759 15552 5773
rect 15518 5691 15552 5701
rect 15518 5623 15552 5629
rect 11334 5352 11354 5398
rect 11456 5352 11532 5398
rect 11334 5330 11532 5352
rect 13032 5366 13230 5472
rect 14286 5470 14896 5504
rect 15518 5555 15552 5557
rect 15518 5519 15552 5521
rect -868 5283 -834 5311
rect 13032 5320 13094 5366
rect 13196 5320 13230 5366
rect 13032 5306 13230 5320
rect 14488 5372 14686 5470
rect 14488 5326 14510 5372
rect 14612 5326 14686 5372
rect 14488 5310 14686 5326
rect 15518 5447 15552 5453
rect 15518 5375 15552 5385
rect -868 5215 -834 5239
rect -868 5147 -834 5167
rect 15518 5303 15552 5317
rect 15518 5231 15552 5249
rect 15518 5159 15552 5181
rect -868 5079 -834 5095
rect 1580 5028 1614 5090
rect -868 5011 -834 5023
rect 1482 4994 1908 5028
rect 4536 5012 4570 5074
rect 7566 5012 7600 5074
rect 15518 5087 15552 5113
rect -868 4934 -834 4951
rect -1554 4842 -932 4876
rect 1484 4929 1518 4994
rect 1484 4857 1518 4869
rect -1162 4840 -1124 4842
rect -23596 4805 -18094 4826
rect -23596 4635 -23548 4805
rect -18142 4635 -18094 4805
rect -23596 4614 -18094 4635
rect -16766 4817 -11264 4838
rect -16766 4647 -16718 4817
rect -11312 4647 -11264 4817
rect -16766 4626 -11264 4647
rect -10300 4815 -4798 4836
rect -10300 4645 -10252 4815
rect -4846 4645 -4798 4815
rect -1158 4768 -1124 4840
rect 1484 4785 1518 4801
rect -1083 4768 -1067 4769
rect -1158 4735 -1067 4768
rect -1033 4735 -1017 4769
rect -1158 4734 -1068 4735
rect -23584 4534 -18104 4614
rect -16756 4546 -11276 4626
rect -10300 4624 -4798 4645
rect 1484 4713 1518 4733
rect 1484 4641 1518 4665
rect -23586 4522 -18076 4534
rect -23586 4500 -21632 4522
rect -23586 4427 -23552 4500
rect -23586 4355 -23552 4367
rect -23586 4283 -23552 4299
rect -23586 4211 -23552 4231
rect -23586 4139 -23552 4163
rect -23586 4067 -23552 4095
rect -23586 3995 -23552 4027
rect -23586 3925 -23552 3959
rect -23586 3857 -23552 3889
rect -23586 3789 -23552 3817
rect -23586 3721 -23552 3745
rect -23586 3653 -23552 3673
rect -23586 3585 -23552 3601
rect -23586 3517 -23552 3529
rect -23586 3438 -23552 3457
rect -23490 4427 -23456 4446
rect -23490 4355 -23456 4367
rect -23490 4283 -23456 4299
rect -23490 4211 -23456 4231
rect -23490 4139 -23456 4163
rect -23490 4067 -23456 4095
rect -23490 3995 -23456 4027
rect -23490 3925 -23456 3959
rect -23490 3857 -23456 3889
rect -23490 3789 -23456 3817
rect -23490 3721 -23456 3745
rect -23490 3653 -23456 3673
rect -23490 3585 -23456 3601
rect -23490 3517 -23456 3529
rect -23490 3392 -23456 3457
rect -23394 4427 -23360 4500
rect -23394 4355 -23360 4367
rect -23394 4283 -23360 4299
rect -23394 4211 -23360 4231
rect -23394 4139 -23360 4163
rect -23394 4067 -23360 4095
rect -23394 3995 -23360 4027
rect -23394 3925 -23360 3959
rect -23394 3857 -23360 3889
rect -23394 3789 -23360 3817
rect -23394 3721 -23360 3745
rect -23394 3653 -23360 3673
rect -23394 3585 -23360 3601
rect -23394 3517 -23360 3529
rect -23394 3438 -23360 3457
rect -23298 4427 -23264 4446
rect -23298 4355 -23264 4367
rect -23298 4283 -23264 4299
rect -23298 4211 -23264 4231
rect -23298 4139 -23264 4163
rect -23298 4067 -23264 4095
rect -23298 3995 -23264 4027
rect -23298 3925 -23264 3959
rect -23298 3857 -23264 3889
rect -23298 3789 -23264 3817
rect -23298 3721 -23264 3745
rect -23298 3653 -23264 3673
rect -23298 3585 -23264 3601
rect -23298 3517 -23264 3529
rect -23298 3392 -23264 3457
rect -23202 4427 -23168 4500
rect -23202 4355 -23168 4367
rect -23202 4283 -23168 4299
rect -23202 4211 -23168 4231
rect -23202 4139 -23168 4163
rect -23202 4067 -23168 4095
rect -23202 3995 -23168 4027
rect -23202 3925 -23168 3959
rect -23202 3857 -23168 3889
rect -23202 3789 -23168 3817
rect -23202 3721 -23168 3745
rect -23202 3653 -23168 3673
rect -23202 3585 -23168 3601
rect -23202 3517 -23168 3529
rect -23202 3438 -23168 3457
rect -23106 4427 -23072 4446
rect -23106 4355 -23072 4367
rect -23106 4283 -23072 4299
rect -23106 4211 -23072 4231
rect -23106 4139 -23072 4163
rect -23106 4067 -23072 4095
rect -23106 3995 -23072 4027
rect -23106 3925 -23072 3959
rect -23106 3857 -23072 3889
rect -23106 3789 -23072 3817
rect -23106 3721 -23072 3745
rect -23106 3653 -23072 3673
rect -23106 3585 -23072 3601
rect -23106 3517 -23072 3529
rect -23106 3392 -23072 3457
rect -23010 4427 -22976 4500
rect -23010 4355 -22976 4367
rect -23010 4283 -22976 4299
rect -23010 4211 -22976 4231
rect -23010 4139 -22976 4163
rect -23010 4067 -22976 4095
rect -23010 3995 -22976 4027
rect -23010 3925 -22976 3959
rect -23010 3857 -22976 3889
rect -23010 3789 -22976 3817
rect -23010 3721 -22976 3745
rect -23010 3653 -22976 3673
rect -23010 3585 -22976 3601
rect -23010 3517 -22976 3529
rect -23010 3438 -22976 3457
rect -22914 4427 -22880 4446
rect -22914 4355 -22880 4367
rect -22914 4283 -22880 4299
rect -22914 4211 -22880 4231
rect -22914 4139 -22880 4163
rect -22914 4067 -22880 4095
rect -22914 3995 -22880 4027
rect -22914 3925 -22880 3959
rect -22914 3857 -22880 3889
rect -22914 3789 -22880 3817
rect -22914 3721 -22880 3745
rect -22914 3653 -22880 3673
rect -22914 3585 -22880 3601
rect -22914 3517 -22880 3529
rect -22914 3392 -22880 3457
rect -22818 4427 -22784 4500
rect -22818 4355 -22784 4367
rect -22818 4283 -22784 4299
rect -22818 4211 -22784 4231
rect -22818 4139 -22784 4163
rect -22818 4067 -22784 4095
rect -22818 3995 -22784 4027
rect -22818 3925 -22784 3959
rect -22818 3857 -22784 3889
rect -22818 3789 -22784 3817
rect -22818 3721 -22784 3745
rect -22818 3653 -22784 3673
rect -22818 3585 -22784 3601
rect -22818 3517 -22784 3529
rect -22818 3438 -22784 3457
rect -22722 4427 -22688 4446
rect -22722 4355 -22688 4367
rect -22722 4283 -22688 4299
rect -22722 4211 -22688 4231
rect -22722 4139 -22688 4163
rect -22722 4067 -22688 4095
rect -22722 3995 -22688 4027
rect -22722 3925 -22688 3959
rect -22722 3857 -22688 3889
rect -22722 3789 -22688 3817
rect -22722 3721 -22688 3745
rect -22722 3653 -22688 3673
rect -22722 3585 -22688 3601
rect -22722 3517 -22688 3529
rect -22722 3392 -22688 3457
rect -22626 4427 -22592 4500
rect -22626 4355 -22592 4367
rect -22626 4283 -22592 4299
rect -22626 4211 -22592 4231
rect -22626 4139 -22592 4163
rect -22626 4067 -22592 4095
rect -22626 3995 -22592 4027
rect -22626 3925 -22592 3959
rect -22626 3857 -22592 3889
rect -22626 3789 -22592 3817
rect -22626 3721 -22592 3745
rect -22626 3653 -22592 3673
rect -22626 3585 -22592 3601
rect -22626 3517 -22592 3529
rect -22626 3438 -22592 3457
rect -22530 4427 -22496 4446
rect -22530 4355 -22496 4367
rect -22530 4283 -22496 4299
rect -22530 4211 -22496 4231
rect -22530 4139 -22496 4163
rect -22530 4067 -22496 4095
rect -22530 3995 -22496 4027
rect -22530 3925 -22496 3959
rect -22530 3857 -22496 3889
rect -22530 3789 -22496 3817
rect -22530 3721 -22496 3745
rect -22530 3653 -22496 3673
rect -22530 3585 -22496 3601
rect -22530 3517 -22496 3529
rect -22530 3392 -22496 3457
rect -22434 4427 -22400 4500
rect -22434 4355 -22400 4367
rect -22434 4283 -22400 4299
rect -22434 4211 -22400 4231
rect -22434 4139 -22400 4163
rect -22434 4067 -22400 4095
rect -22434 3995 -22400 4027
rect -22434 3925 -22400 3959
rect -22434 3857 -22400 3889
rect -22434 3789 -22400 3817
rect -22434 3721 -22400 3745
rect -22434 3653 -22400 3673
rect -22434 3585 -22400 3601
rect -22434 3517 -22400 3529
rect -22434 3438 -22400 3457
rect -22338 4427 -22304 4446
rect -22338 4355 -22304 4367
rect -22338 4283 -22304 4299
rect -22338 4211 -22304 4231
rect -22338 4139 -22304 4163
rect -22338 4067 -22304 4095
rect -22338 3995 -22304 4027
rect -22338 3925 -22304 3959
rect -22338 3857 -22304 3889
rect -22338 3789 -22304 3817
rect -22338 3721 -22304 3745
rect -22338 3653 -22304 3673
rect -22338 3585 -22304 3601
rect -22338 3517 -22304 3529
rect -22338 3392 -22304 3457
rect -22242 4427 -22208 4500
rect -22242 4355 -22208 4367
rect -22242 4283 -22208 4299
rect -22242 4211 -22208 4231
rect -22242 4139 -22208 4163
rect -22242 4067 -22208 4095
rect -22242 3995 -22208 4027
rect -22242 3925 -22208 3959
rect -22242 3857 -22208 3889
rect -22242 3789 -22208 3817
rect -22242 3721 -22208 3745
rect -22242 3653 -22208 3673
rect -22242 3585 -22208 3601
rect -22242 3517 -22208 3529
rect -22242 3438 -22208 3457
rect -22146 4427 -22112 4446
rect -22146 4355 -22112 4367
rect -22146 4283 -22112 4299
rect -22146 4211 -22112 4231
rect -22146 4139 -22112 4163
rect -22146 4067 -22112 4095
rect -22146 3995 -22112 4027
rect -22146 3925 -22112 3959
rect -22146 3857 -22112 3889
rect -22146 3789 -22112 3817
rect -22146 3721 -22112 3745
rect -22146 3653 -22112 3673
rect -22146 3585 -22112 3601
rect -22146 3517 -22112 3529
rect -22146 3392 -22112 3457
rect -22050 4427 -22016 4500
rect -22050 4355 -22016 4367
rect -22050 4283 -22016 4299
rect -22050 4211 -22016 4231
rect -22050 4139 -22016 4163
rect -22050 4067 -22016 4095
rect -22050 3995 -22016 4027
rect -22050 3925 -22016 3959
rect -22050 3857 -22016 3889
rect -22050 3789 -22016 3817
rect -22050 3721 -22016 3745
rect -22050 3653 -22016 3673
rect -22050 3585 -22016 3601
rect -22050 3517 -22016 3529
rect -22050 3438 -22016 3457
rect -21954 4427 -21920 4446
rect -21954 4355 -21920 4367
rect -21954 4283 -21920 4299
rect -21954 4211 -21920 4231
rect -21954 4139 -21920 4163
rect -21954 4067 -21920 4095
rect -21954 3995 -21920 4027
rect -21954 3925 -21920 3959
rect -21954 3857 -21920 3889
rect -21954 3789 -21920 3817
rect -21954 3721 -21920 3745
rect -21954 3653 -21920 3673
rect -21954 3585 -21920 3601
rect -21954 3517 -21920 3529
rect -21954 3392 -21920 3457
rect -21858 4427 -21824 4500
rect -21858 4355 -21824 4367
rect -21858 4283 -21824 4299
rect -21858 4211 -21824 4231
rect -21858 4139 -21824 4163
rect -21858 4067 -21824 4095
rect -21858 3995 -21824 4027
rect -21858 3925 -21824 3959
rect -21858 3857 -21824 3889
rect -21858 3789 -21824 3817
rect -21858 3721 -21824 3745
rect -21858 3653 -21824 3673
rect -21858 3585 -21824 3601
rect -21858 3517 -21824 3529
rect -21858 3438 -21824 3457
rect -21762 4427 -21728 4446
rect -21762 4355 -21728 4367
rect -21762 4283 -21728 4299
rect -21762 4211 -21728 4231
rect -21762 4139 -21728 4163
rect -21762 4067 -21728 4095
rect -21762 3995 -21728 4027
rect -21762 3925 -21728 3959
rect -21762 3857 -21728 3889
rect -21762 3789 -21728 3817
rect -21762 3721 -21728 3745
rect -21762 3653 -21728 3673
rect -21762 3585 -21728 3601
rect -21762 3517 -21728 3529
rect -21762 3392 -21728 3457
rect -21666 4427 -21632 4500
rect -21346 4494 -19968 4522
rect -21666 4355 -21632 4367
rect -21666 4283 -21632 4299
rect -21666 4211 -21632 4231
rect -21666 4139 -21632 4163
rect -21666 4067 -21632 4095
rect -21666 3995 -21632 4027
rect -21666 3925 -21632 3959
rect -21666 3857 -21632 3889
rect -21666 3789 -21632 3817
rect -21666 3721 -21632 3745
rect -21666 3653 -21632 3673
rect -21666 3585 -21632 3601
rect -21666 3517 -21632 3529
rect -21666 3438 -21632 3457
rect -21442 4433 -21408 4452
rect -21442 4361 -21408 4373
rect -21442 4289 -21408 4305
rect -21442 4217 -21408 4237
rect -21442 4145 -21408 4169
rect -21442 4073 -21408 4101
rect -21442 4001 -21408 4033
rect -21442 3931 -21408 3965
rect -21442 3863 -21408 3895
rect -21442 3795 -21408 3823
rect -21442 3727 -21408 3751
rect -21442 3659 -21408 3679
rect -21442 3591 -21408 3607
rect -21442 3523 -21408 3535
rect -23490 3358 -21728 3392
rect -21442 3386 -21408 3463
rect -21346 4433 -21312 4494
rect -21346 4361 -21312 4373
rect -21346 4289 -21312 4305
rect -21346 4217 -21312 4237
rect -21346 4145 -21312 4169
rect -21346 4073 -21312 4101
rect -21346 4001 -21312 4033
rect -21346 3931 -21312 3965
rect -21346 3863 -21312 3895
rect -21346 3795 -21312 3823
rect -21346 3727 -21312 3751
rect -21346 3659 -21312 3679
rect -21346 3591 -21312 3607
rect -21346 3523 -21312 3535
rect -21346 3444 -21312 3463
rect -21250 4433 -21216 4452
rect -21250 4361 -21216 4373
rect -21250 4289 -21216 4305
rect -21250 4217 -21216 4237
rect -21250 4145 -21216 4169
rect -21250 4073 -21216 4101
rect -21250 4001 -21216 4033
rect -21250 3931 -21216 3965
rect -21250 3863 -21216 3895
rect -21250 3795 -21216 3823
rect -21250 3727 -21216 3751
rect -21250 3659 -21216 3679
rect -21250 3591 -21216 3607
rect -21250 3523 -21216 3535
rect -21250 3386 -21216 3463
rect -21154 4433 -21120 4494
rect -21154 4361 -21120 4373
rect -21154 4289 -21120 4305
rect -21154 4217 -21120 4237
rect -21154 4145 -21120 4169
rect -21154 4073 -21120 4101
rect -21154 4001 -21120 4033
rect -21154 3931 -21120 3965
rect -21154 3863 -21120 3895
rect -21154 3795 -21120 3823
rect -21154 3727 -21120 3751
rect -21154 3659 -21120 3679
rect -21154 3591 -21120 3607
rect -21154 3523 -21120 3535
rect -21154 3444 -21120 3463
rect -21058 4433 -21024 4452
rect -21058 4361 -21024 4373
rect -21058 4289 -21024 4305
rect -21058 4217 -21024 4237
rect -21058 4145 -21024 4169
rect -21058 4073 -21024 4101
rect -21058 4001 -21024 4033
rect -21058 3931 -21024 3965
rect -21058 3863 -21024 3895
rect -21058 3795 -21024 3823
rect -21058 3727 -21024 3751
rect -21058 3659 -21024 3679
rect -21058 3591 -21024 3607
rect -21058 3523 -21024 3535
rect -21058 3386 -21024 3463
rect -20962 4433 -20928 4494
rect -20962 4361 -20928 4373
rect -20962 4289 -20928 4305
rect -20962 4217 -20928 4237
rect -20962 4145 -20928 4169
rect -20962 4073 -20928 4101
rect -20962 4001 -20928 4033
rect -20962 3931 -20928 3965
rect -20962 3863 -20928 3895
rect -20962 3795 -20928 3823
rect -20962 3727 -20928 3751
rect -20962 3659 -20928 3679
rect -20962 3591 -20928 3607
rect -20962 3523 -20928 3535
rect -20962 3444 -20928 3463
rect -20866 4433 -20832 4452
rect -20866 4361 -20832 4373
rect -20866 4289 -20832 4305
rect -20866 4217 -20832 4237
rect -20866 4145 -20832 4169
rect -20866 4073 -20832 4101
rect -20866 4001 -20832 4033
rect -20866 3931 -20832 3965
rect -20866 3863 -20832 3895
rect -20866 3795 -20832 3823
rect -20866 3727 -20832 3751
rect -20866 3659 -20832 3679
rect -20866 3591 -20832 3607
rect -20866 3523 -20832 3535
rect -20866 3386 -20832 3463
rect -20770 4433 -20736 4494
rect -20770 4361 -20736 4373
rect -20770 4289 -20736 4305
rect -20770 4217 -20736 4237
rect -20770 4145 -20736 4169
rect -20770 4073 -20736 4101
rect -20770 4001 -20736 4033
rect -20770 3931 -20736 3965
rect -20770 3863 -20736 3895
rect -20770 3795 -20736 3823
rect -20770 3727 -20736 3751
rect -20770 3659 -20736 3679
rect -20770 3591 -20736 3607
rect -20770 3523 -20736 3535
rect -20770 3444 -20736 3463
rect -20674 4433 -20640 4452
rect -20674 4361 -20640 4373
rect -20674 4289 -20640 4305
rect -20674 4217 -20640 4237
rect -20674 4145 -20640 4169
rect -20674 4073 -20640 4101
rect -20674 4001 -20640 4033
rect -20674 3931 -20640 3965
rect -20674 3863 -20640 3895
rect -20674 3795 -20640 3823
rect -20674 3727 -20640 3751
rect -20674 3659 -20640 3679
rect -20674 3591 -20640 3607
rect -20674 3523 -20640 3535
rect -20674 3386 -20640 3463
rect -20578 4433 -20544 4494
rect -20578 4361 -20544 4373
rect -20578 4289 -20544 4305
rect -20578 4217 -20544 4237
rect -20578 4145 -20544 4169
rect -20578 4073 -20544 4101
rect -20578 4001 -20544 4033
rect -20578 3931 -20544 3965
rect -20578 3863 -20544 3895
rect -20578 3795 -20544 3823
rect -20578 3727 -20544 3751
rect -20578 3659 -20544 3679
rect -20578 3591 -20544 3607
rect -20578 3523 -20544 3535
rect -20578 3444 -20544 3463
rect -20482 4433 -20448 4452
rect -20482 4361 -20448 4373
rect -20482 4289 -20448 4305
rect -20482 4217 -20448 4237
rect -20482 4145 -20448 4169
rect -20482 4073 -20448 4101
rect -20482 4001 -20448 4033
rect -20482 3931 -20448 3965
rect -20482 3863 -20448 3895
rect -20482 3795 -20448 3823
rect -20482 3727 -20448 3751
rect -20482 3659 -20448 3679
rect -20482 3591 -20448 3607
rect -20482 3523 -20448 3535
rect -20482 3386 -20448 3463
rect -20386 4433 -20352 4494
rect -20386 4361 -20352 4373
rect -20386 4289 -20352 4305
rect -20386 4217 -20352 4237
rect -20386 4145 -20352 4169
rect -20386 4073 -20352 4101
rect -20386 4001 -20352 4033
rect -20386 3931 -20352 3965
rect -20386 3863 -20352 3895
rect -20386 3795 -20352 3823
rect -20386 3727 -20352 3751
rect -20386 3659 -20352 3679
rect -20386 3591 -20352 3607
rect -20386 3523 -20352 3535
rect -20386 3444 -20352 3463
rect -20290 4433 -20256 4452
rect -20290 4361 -20256 4373
rect -20290 4289 -20256 4305
rect -20290 4217 -20256 4237
rect -20290 4145 -20256 4169
rect -20290 4073 -20256 4101
rect -20290 4001 -20256 4033
rect -20290 3931 -20256 3965
rect -20290 3863 -20256 3895
rect -20290 3795 -20256 3823
rect -20290 3727 -20256 3751
rect -20290 3659 -20256 3679
rect -20290 3591 -20256 3607
rect -20290 3523 -20256 3535
rect -20290 3386 -20256 3463
rect -20194 4433 -20160 4494
rect -20194 4361 -20160 4373
rect -20194 4289 -20160 4305
rect -20194 4217 -20160 4237
rect -20194 4145 -20160 4169
rect -20194 4073 -20160 4101
rect -20194 4001 -20160 4033
rect -20194 3931 -20160 3965
rect -20194 3863 -20160 3895
rect -20194 3795 -20160 3823
rect -20194 3727 -20160 3751
rect -20194 3659 -20160 3679
rect -20194 3591 -20160 3607
rect -20194 3523 -20160 3535
rect -20194 3444 -20160 3463
rect -20098 4433 -20064 4452
rect -20098 4361 -20064 4373
rect -20098 4289 -20064 4305
rect -20098 4217 -20064 4237
rect -20098 4145 -20064 4169
rect -20098 4073 -20064 4101
rect -20098 4001 -20064 4033
rect -20098 3931 -20064 3965
rect -20098 3863 -20064 3895
rect -20098 3795 -20064 3823
rect -20098 3727 -20064 3751
rect -20098 3659 -20064 3679
rect -20098 3591 -20064 3607
rect -20098 3523 -20064 3535
rect -20098 3386 -20064 3463
rect -20002 4433 -19968 4494
rect -20002 4361 -19968 4373
rect -20002 4289 -19968 4305
rect -20002 4217 -19968 4237
rect -20002 4145 -19968 4169
rect -20002 4073 -19968 4101
rect -20002 4001 -19968 4033
rect -20002 3931 -19968 3965
rect -20002 3863 -19968 3895
rect -20002 3795 -19968 3823
rect -20002 3727 -19968 3751
rect -20002 3659 -19968 3679
rect -20002 3591 -19968 3607
rect -20002 3523 -19968 3535
rect -20002 3444 -19968 3463
rect -19758 4498 -18764 4522
rect -19758 4439 -19724 4498
rect -19758 4367 -19724 4379
rect -19758 4295 -19724 4311
rect -19758 4223 -19724 4243
rect -19758 4151 -19724 4175
rect -19758 4079 -19724 4107
rect -19758 4007 -19724 4039
rect -19758 3937 -19724 3971
rect -19758 3869 -19724 3901
rect -19758 3801 -19724 3829
rect -19758 3733 -19724 3757
rect -19758 3665 -19724 3685
rect -19758 3597 -19724 3613
rect -19758 3529 -19724 3541
rect -19758 3450 -19724 3469
rect -19662 4439 -19628 4458
rect -19662 4367 -19628 4379
rect -19662 4295 -19628 4311
rect -19662 4223 -19628 4243
rect -19662 4151 -19628 4175
rect -19662 4079 -19628 4107
rect -19662 4007 -19628 4039
rect -19662 3937 -19628 3971
rect -19662 3869 -19628 3901
rect -19662 3801 -19628 3829
rect -19662 3733 -19628 3757
rect -19662 3665 -19628 3685
rect -19662 3597 -19628 3613
rect -19662 3529 -19628 3541
rect -22980 3130 -22934 3358
rect -21442 3352 -20064 3386
rect -19662 3392 -19628 3469
rect -19566 4439 -19532 4498
rect -19566 4367 -19532 4379
rect -19566 4295 -19532 4311
rect -19566 4223 -19532 4243
rect -19566 4151 -19532 4175
rect -19566 4079 -19532 4107
rect -19566 4007 -19532 4039
rect -19566 3937 -19532 3971
rect -19566 3869 -19532 3901
rect -19566 3801 -19532 3829
rect -19566 3733 -19532 3757
rect -19566 3665 -19532 3685
rect -19566 3597 -19532 3613
rect -19566 3529 -19532 3541
rect -19566 3450 -19532 3469
rect -19470 4439 -19436 4458
rect -19470 4367 -19436 4379
rect -19470 4295 -19436 4311
rect -19470 4223 -19436 4243
rect -19470 4151 -19436 4175
rect -19470 4079 -19436 4107
rect -19470 4007 -19436 4039
rect -19470 3937 -19436 3971
rect -19470 3869 -19436 3901
rect -19470 3801 -19436 3829
rect -19470 3733 -19436 3757
rect -19470 3665 -19436 3685
rect -19470 3597 -19436 3613
rect -19470 3529 -19436 3541
rect -19470 3392 -19436 3469
rect -19374 4439 -19340 4498
rect -19374 4367 -19340 4379
rect -19374 4295 -19340 4311
rect -19374 4223 -19340 4243
rect -19374 4151 -19340 4175
rect -19374 4079 -19340 4107
rect -19374 4007 -19340 4039
rect -19374 3937 -19340 3971
rect -19374 3869 -19340 3901
rect -19374 3801 -19340 3829
rect -19374 3733 -19340 3757
rect -19374 3665 -19340 3685
rect -19374 3597 -19340 3613
rect -19374 3529 -19340 3541
rect -19374 3450 -19340 3469
rect -19278 4439 -19244 4458
rect -19278 4367 -19244 4379
rect -19278 4295 -19244 4311
rect -19278 4223 -19244 4243
rect -19278 4151 -19244 4175
rect -19278 4079 -19244 4107
rect -19278 4007 -19244 4039
rect -19278 3937 -19244 3971
rect -19278 3869 -19244 3901
rect -19278 3801 -19244 3829
rect -19278 3733 -19244 3757
rect -19278 3665 -19244 3685
rect -19278 3597 -19244 3613
rect -19278 3529 -19244 3541
rect -19278 3392 -19244 3469
rect -19182 4439 -19148 4498
rect -19182 4367 -19148 4379
rect -19182 4295 -19148 4311
rect -19182 4223 -19148 4243
rect -19182 4151 -19148 4175
rect -19182 4079 -19148 4107
rect -19182 4007 -19148 4039
rect -19182 3937 -19148 3971
rect -19182 3869 -19148 3901
rect -19182 3801 -19148 3829
rect -19182 3733 -19148 3757
rect -19182 3665 -19148 3685
rect -19182 3597 -19148 3613
rect -19182 3529 -19148 3541
rect -19182 3450 -19148 3469
rect -19086 4439 -19052 4458
rect -19086 4367 -19052 4379
rect -19086 4295 -19052 4311
rect -19086 4223 -19052 4243
rect -19086 4151 -19052 4175
rect -19086 4079 -19052 4107
rect -19086 4007 -19052 4039
rect -19086 3937 -19052 3971
rect -19086 3869 -19052 3901
rect -19086 3801 -19052 3829
rect -19086 3733 -19052 3757
rect -19086 3665 -19052 3685
rect -19086 3597 -19052 3613
rect -19086 3529 -19052 3541
rect -19086 3392 -19052 3469
rect -18990 4439 -18956 4498
rect -18990 4367 -18956 4379
rect -18990 4295 -18956 4311
rect -18990 4223 -18956 4243
rect -18990 4151 -18956 4175
rect -18990 4079 -18956 4107
rect -18990 4007 -18956 4039
rect -18990 3937 -18956 3971
rect -18990 3869 -18956 3901
rect -18990 3801 -18956 3829
rect -18990 3733 -18956 3757
rect -18990 3665 -18956 3685
rect -18990 3597 -18956 3613
rect -18990 3529 -18956 3541
rect -18990 3450 -18956 3469
rect -18894 4439 -18860 4458
rect -18894 4367 -18860 4379
rect -18894 4295 -18860 4311
rect -18894 4223 -18860 4243
rect -18894 4151 -18860 4175
rect -18894 4079 -18860 4107
rect -18894 4007 -18860 4039
rect -18894 3937 -18860 3971
rect -18894 3869 -18860 3901
rect -18894 3801 -18860 3829
rect -18894 3733 -18860 3757
rect -18894 3665 -18860 3685
rect -18894 3597 -18860 3613
rect -18894 3529 -18860 3541
rect -18894 3392 -18860 3469
rect -18798 4439 -18764 4498
rect -18494 4500 -18076 4522
rect -18798 4367 -18764 4379
rect -18798 4295 -18764 4311
rect -18798 4223 -18764 4243
rect -18798 4151 -18764 4175
rect -18798 4079 -18764 4107
rect -18798 4007 -18764 4039
rect -18798 3937 -18764 3971
rect -18798 3869 -18764 3901
rect -18798 3801 -18764 3829
rect -18798 3733 -18764 3757
rect -18798 3665 -18764 3685
rect -18798 3597 -18764 3613
rect -18798 3529 -18764 3541
rect -18798 3450 -18764 3469
rect -18590 4441 -18556 4460
rect -18590 4369 -18556 4381
rect -18590 4297 -18556 4313
rect -18590 4225 -18556 4245
rect -18590 4153 -18556 4177
rect -18590 4081 -18556 4109
rect -18590 4009 -18556 4041
rect -18590 3939 -18556 3973
rect -18590 3871 -18556 3903
rect -18590 3803 -18556 3831
rect -18590 3735 -18556 3759
rect -18590 3667 -18556 3687
rect -18590 3599 -18556 3615
rect -18590 3531 -18556 3543
rect -19662 3358 -18860 3392
rect -18590 3400 -18556 3471
rect -18494 4441 -18460 4500
rect -18494 4369 -18460 4381
rect -18494 4297 -18460 4313
rect -18494 4225 -18460 4245
rect -18494 4153 -18460 4177
rect -18494 4081 -18460 4109
rect -18494 4009 -18460 4041
rect -18494 3939 -18460 3973
rect -18494 3871 -18460 3903
rect -18494 3803 -18460 3831
rect -18494 3735 -18460 3759
rect -18494 3667 -18460 3687
rect -18494 3599 -18460 3615
rect -18494 3531 -18460 3543
rect -18494 3452 -18460 3471
rect -18398 4441 -18364 4460
rect -18398 4369 -18364 4381
rect -18398 4297 -18364 4313
rect -18398 4225 -18364 4245
rect -18398 4153 -18364 4177
rect -18398 4081 -18364 4109
rect -18398 4009 -18364 4041
rect -18398 3939 -18364 3973
rect -18398 3871 -18364 3903
rect -18398 3803 -18364 3831
rect -18398 3735 -18364 3759
rect -18398 3667 -18364 3687
rect -18398 3599 -18364 3615
rect -18398 3531 -18364 3543
rect -18398 3400 -18364 3471
rect -18302 4441 -18268 4500
rect -18302 4369 -18268 4381
rect -18302 4297 -18268 4313
rect -18302 4225 -18268 4245
rect -18302 4153 -18268 4177
rect -18302 4081 -18268 4109
rect -18302 4009 -18268 4041
rect -18302 3939 -18268 3973
rect -18302 3871 -18268 3903
rect -18302 3803 -18268 3831
rect -18302 3735 -18268 3759
rect -18302 3667 -18268 3687
rect -18302 3599 -18268 3615
rect -18302 3531 -18268 3543
rect -18302 3452 -18268 3471
rect -18206 4441 -18172 4460
rect -18206 4369 -18172 4381
rect -18206 4297 -18172 4313
rect -18206 4225 -18172 4245
rect -18206 4153 -18172 4177
rect -18206 4081 -18172 4109
rect -18206 4009 -18172 4041
rect -18206 3939 -18172 3973
rect -18206 3871 -18172 3903
rect -18206 3803 -18172 3831
rect -18206 3735 -18172 3759
rect -18206 3667 -18172 3687
rect -18206 3599 -18172 3615
rect -18206 3531 -18172 3543
rect -18206 3400 -18172 3471
rect -18110 4441 -18076 4500
rect -18110 4369 -18076 4381
rect -18110 4297 -18076 4313
rect -18110 4225 -18076 4245
rect -18110 4153 -18076 4177
rect -18110 4081 -18076 4109
rect -18110 4009 -18076 4041
rect -18110 3939 -18076 3973
rect -18110 3871 -18076 3903
rect -18110 3803 -18076 3831
rect -18110 3735 -18076 3759
rect -18110 3667 -18076 3687
rect -18110 3599 -18076 3615
rect -18110 3531 -18076 3543
rect -18110 3452 -18076 3471
rect -16756 4524 -11246 4546
rect -10292 4544 -4812 4624
rect 1484 4569 1518 4597
rect -10292 4532 -4780 4544
rect -16756 4512 -14802 4524
rect -16756 4439 -16722 4512
rect -16756 4367 -16722 4379
rect -16756 4295 -16722 4311
rect -16756 4223 -16722 4243
rect -16756 4151 -16722 4175
rect -16756 4079 -16722 4107
rect -16756 4007 -16722 4039
rect -16756 3937 -16722 3971
rect -16756 3869 -16722 3901
rect -16756 3801 -16722 3829
rect -16756 3733 -16722 3757
rect -16756 3665 -16722 3685
rect -16756 3597 -16722 3613
rect -16756 3529 -16722 3541
rect -16756 3450 -16722 3469
rect -16660 4439 -16626 4458
rect -16660 4367 -16626 4379
rect -16660 4295 -16626 4311
rect -16660 4223 -16626 4243
rect -16660 4151 -16626 4175
rect -16660 4079 -16626 4107
rect -16660 4007 -16626 4039
rect -16660 3937 -16626 3971
rect -16660 3869 -16626 3901
rect -16660 3801 -16626 3829
rect -16660 3733 -16626 3757
rect -16660 3665 -16626 3685
rect -16660 3597 -16626 3613
rect -16660 3529 -16626 3541
rect -16660 3404 -16626 3469
rect -16564 4439 -16530 4512
rect -16564 4367 -16530 4379
rect -16564 4295 -16530 4311
rect -16564 4223 -16530 4243
rect -16564 4151 -16530 4175
rect -16564 4079 -16530 4107
rect -16564 4007 -16530 4039
rect -16564 3937 -16530 3971
rect -16564 3869 -16530 3901
rect -16564 3801 -16530 3829
rect -16564 3733 -16530 3757
rect -16564 3665 -16530 3685
rect -16564 3597 -16530 3613
rect -16564 3529 -16530 3541
rect -16564 3450 -16530 3469
rect -16468 4439 -16434 4458
rect -16468 4367 -16434 4379
rect -16468 4295 -16434 4311
rect -16468 4223 -16434 4243
rect -16468 4151 -16434 4175
rect -16468 4079 -16434 4107
rect -16468 4007 -16434 4039
rect -16468 3937 -16434 3971
rect -16468 3869 -16434 3901
rect -16468 3801 -16434 3829
rect -16468 3733 -16434 3757
rect -16468 3665 -16434 3685
rect -16468 3597 -16434 3613
rect -16468 3529 -16434 3541
rect -16468 3404 -16434 3469
rect -16372 4439 -16338 4512
rect -16372 4367 -16338 4379
rect -16372 4295 -16338 4311
rect -16372 4223 -16338 4243
rect -16372 4151 -16338 4175
rect -16372 4079 -16338 4107
rect -16372 4007 -16338 4039
rect -16372 3937 -16338 3971
rect -16372 3869 -16338 3901
rect -16372 3801 -16338 3829
rect -16372 3733 -16338 3757
rect -16372 3665 -16338 3685
rect -16372 3597 -16338 3613
rect -16372 3529 -16338 3541
rect -16372 3450 -16338 3469
rect -16276 4439 -16242 4458
rect -16276 4367 -16242 4379
rect -16276 4295 -16242 4311
rect -16276 4223 -16242 4243
rect -16276 4151 -16242 4175
rect -16276 4079 -16242 4107
rect -16276 4007 -16242 4039
rect -16276 3937 -16242 3971
rect -16276 3869 -16242 3901
rect -16276 3801 -16242 3829
rect -16276 3733 -16242 3757
rect -16276 3665 -16242 3685
rect -16276 3597 -16242 3613
rect -16276 3529 -16242 3541
rect -16276 3404 -16242 3469
rect -16180 4439 -16146 4512
rect -16180 4367 -16146 4379
rect -16180 4295 -16146 4311
rect -16180 4223 -16146 4243
rect -16180 4151 -16146 4175
rect -16180 4079 -16146 4107
rect -16180 4007 -16146 4039
rect -16180 3937 -16146 3971
rect -16180 3869 -16146 3901
rect -16180 3801 -16146 3829
rect -16180 3733 -16146 3757
rect -16180 3665 -16146 3685
rect -16180 3597 -16146 3613
rect -16180 3529 -16146 3541
rect -16180 3450 -16146 3469
rect -16084 4439 -16050 4458
rect -16084 4367 -16050 4379
rect -16084 4295 -16050 4311
rect -16084 4223 -16050 4243
rect -16084 4151 -16050 4175
rect -16084 4079 -16050 4107
rect -16084 4007 -16050 4039
rect -16084 3937 -16050 3971
rect -16084 3869 -16050 3901
rect -16084 3801 -16050 3829
rect -16084 3733 -16050 3757
rect -16084 3665 -16050 3685
rect -16084 3597 -16050 3613
rect -16084 3529 -16050 3541
rect -16084 3404 -16050 3469
rect -15988 4439 -15954 4512
rect -15988 4367 -15954 4379
rect -15988 4295 -15954 4311
rect -15988 4223 -15954 4243
rect -15988 4151 -15954 4175
rect -15988 4079 -15954 4107
rect -15988 4007 -15954 4039
rect -15988 3937 -15954 3971
rect -15988 3869 -15954 3901
rect -15988 3801 -15954 3829
rect -15988 3733 -15954 3757
rect -15988 3665 -15954 3685
rect -15988 3597 -15954 3613
rect -15988 3529 -15954 3541
rect -15988 3450 -15954 3469
rect -15892 4439 -15858 4458
rect -15892 4367 -15858 4379
rect -15892 4295 -15858 4311
rect -15892 4223 -15858 4243
rect -15892 4151 -15858 4175
rect -15892 4079 -15858 4107
rect -15892 4007 -15858 4039
rect -15892 3937 -15858 3971
rect -15892 3869 -15858 3901
rect -15892 3801 -15858 3829
rect -15892 3733 -15858 3757
rect -15892 3665 -15858 3685
rect -15892 3597 -15858 3613
rect -15892 3529 -15858 3541
rect -15892 3404 -15858 3469
rect -15796 4439 -15762 4512
rect -15796 4367 -15762 4379
rect -15796 4295 -15762 4311
rect -15796 4223 -15762 4243
rect -15796 4151 -15762 4175
rect -15796 4079 -15762 4107
rect -15796 4007 -15762 4039
rect -15796 3937 -15762 3971
rect -15796 3869 -15762 3901
rect -15796 3801 -15762 3829
rect -15796 3733 -15762 3757
rect -15796 3665 -15762 3685
rect -15796 3597 -15762 3613
rect -15796 3529 -15762 3541
rect -15796 3450 -15762 3469
rect -15700 4439 -15666 4458
rect -15700 4367 -15666 4379
rect -15700 4295 -15666 4311
rect -15700 4223 -15666 4243
rect -15700 4151 -15666 4175
rect -15700 4079 -15666 4107
rect -15700 4007 -15666 4039
rect -15700 3937 -15666 3971
rect -15700 3869 -15666 3901
rect -15700 3801 -15666 3829
rect -15700 3733 -15666 3757
rect -15700 3665 -15666 3685
rect -15700 3597 -15666 3613
rect -15700 3529 -15666 3541
rect -15700 3404 -15666 3469
rect -15604 4439 -15570 4512
rect -15604 4367 -15570 4379
rect -15604 4295 -15570 4311
rect -15604 4223 -15570 4243
rect -15604 4151 -15570 4175
rect -15604 4079 -15570 4107
rect -15604 4007 -15570 4039
rect -15604 3937 -15570 3971
rect -15604 3869 -15570 3901
rect -15604 3801 -15570 3829
rect -15604 3733 -15570 3757
rect -15604 3665 -15570 3685
rect -15604 3597 -15570 3613
rect -15604 3529 -15570 3541
rect -15604 3450 -15570 3469
rect -15508 4439 -15474 4458
rect -15508 4367 -15474 4379
rect -15508 4295 -15474 4311
rect -15508 4223 -15474 4243
rect -15508 4151 -15474 4175
rect -15508 4079 -15474 4107
rect -15508 4007 -15474 4039
rect -15508 3937 -15474 3971
rect -15508 3869 -15474 3901
rect -15508 3801 -15474 3829
rect -15508 3733 -15474 3757
rect -15508 3665 -15474 3685
rect -15508 3597 -15474 3613
rect -15508 3529 -15474 3541
rect -15508 3404 -15474 3469
rect -15412 4439 -15378 4512
rect -15412 4367 -15378 4379
rect -15412 4295 -15378 4311
rect -15412 4223 -15378 4243
rect -15412 4151 -15378 4175
rect -15412 4079 -15378 4107
rect -15412 4007 -15378 4039
rect -15412 3937 -15378 3971
rect -15412 3869 -15378 3901
rect -15412 3801 -15378 3829
rect -15412 3733 -15378 3757
rect -15412 3665 -15378 3685
rect -15412 3597 -15378 3613
rect -15412 3529 -15378 3541
rect -15412 3450 -15378 3469
rect -15316 4439 -15282 4458
rect -15316 4367 -15282 4379
rect -15316 4295 -15282 4311
rect -15316 4223 -15282 4243
rect -15316 4151 -15282 4175
rect -15316 4079 -15282 4107
rect -15316 4007 -15282 4039
rect -15316 3937 -15282 3971
rect -15316 3869 -15282 3901
rect -15316 3801 -15282 3829
rect -15316 3733 -15282 3757
rect -15316 3665 -15282 3685
rect -15316 3597 -15282 3613
rect -15316 3529 -15282 3541
rect -15316 3404 -15282 3469
rect -15220 4439 -15186 4512
rect -15220 4367 -15186 4379
rect -15220 4295 -15186 4311
rect -15220 4223 -15186 4243
rect -15220 4151 -15186 4175
rect -15220 4079 -15186 4107
rect -15220 4007 -15186 4039
rect -15220 3937 -15186 3971
rect -15220 3869 -15186 3901
rect -15220 3801 -15186 3829
rect -15220 3733 -15186 3757
rect -15220 3665 -15186 3685
rect -15220 3597 -15186 3613
rect -15220 3529 -15186 3541
rect -15220 3450 -15186 3469
rect -15124 4439 -15090 4458
rect -15124 4367 -15090 4379
rect -15124 4295 -15090 4311
rect -15124 4223 -15090 4243
rect -15124 4151 -15090 4175
rect -15124 4079 -15090 4107
rect -15124 4007 -15090 4039
rect -15124 3937 -15090 3971
rect -15124 3869 -15090 3901
rect -15124 3801 -15090 3829
rect -15124 3733 -15090 3757
rect -15124 3665 -15090 3685
rect -15124 3597 -15090 3613
rect -15124 3529 -15090 3541
rect -15124 3404 -15090 3469
rect -15028 4439 -14994 4512
rect -15028 4367 -14994 4379
rect -15028 4295 -14994 4311
rect -15028 4223 -14994 4243
rect -15028 4151 -14994 4175
rect -15028 4079 -14994 4107
rect -15028 4007 -14994 4039
rect -15028 3937 -14994 3971
rect -15028 3869 -14994 3901
rect -15028 3801 -14994 3829
rect -15028 3733 -14994 3757
rect -15028 3665 -14994 3685
rect -15028 3597 -14994 3613
rect -15028 3529 -14994 3541
rect -15028 3450 -14994 3469
rect -14932 4439 -14898 4458
rect -14932 4367 -14898 4379
rect -14932 4295 -14898 4311
rect -14932 4223 -14898 4243
rect -14932 4151 -14898 4175
rect -14932 4079 -14898 4107
rect -14932 4007 -14898 4039
rect -14932 3937 -14898 3971
rect -14932 3869 -14898 3901
rect -14932 3801 -14898 3829
rect -14932 3733 -14898 3757
rect -14932 3665 -14898 3685
rect -14932 3597 -14898 3613
rect -14932 3529 -14898 3541
rect -14932 3404 -14898 3469
rect -14836 4439 -14802 4512
rect -14516 4506 -13138 4524
rect -14836 4367 -14802 4379
rect -14836 4295 -14802 4311
rect -14836 4223 -14802 4243
rect -14836 4151 -14802 4175
rect -14836 4079 -14802 4107
rect -14836 4007 -14802 4039
rect -14836 3937 -14802 3971
rect -14836 3869 -14802 3901
rect -14836 3801 -14802 3829
rect -14836 3733 -14802 3757
rect -14836 3665 -14802 3685
rect -14836 3597 -14802 3613
rect -14836 3529 -14802 3541
rect -14836 3450 -14802 3469
rect -14612 4445 -14578 4464
rect -14612 4373 -14578 4385
rect -14612 4301 -14578 4317
rect -14612 4229 -14578 4249
rect -14612 4157 -14578 4181
rect -14612 4085 -14578 4113
rect -14612 4013 -14578 4045
rect -14612 3943 -14578 3977
rect -14612 3875 -14578 3907
rect -14612 3807 -14578 3835
rect -14612 3739 -14578 3763
rect -14612 3671 -14578 3691
rect -14612 3603 -14578 3619
rect -14612 3535 -14578 3547
rect -18590 3366 -18170 3400
rect -16660 3370 -14898 3404
rect -14612 3398 -14578 3475
rect -14516 4445 -14482 4506
rect -14516 4373 -14482 4385
rect -14516 4301 -14482 4317
rect -14516 4229 -14482 4249
rect -14516 4157 -14482 4181
rect -14516 4085 -14482 4113
rect -14516 4013 -14482 4045
rect -14516 3943 -14482 3977
rect -14516 3875 -14482 3907
rect -14516 3807 -14482 3835
rect -14516 3739 -14482 3763
rect -14516 3671 -14482 3691
rect -14516 3603 -14482 3619
rect -14516 3535 -14482 3547
rect -14516 3456 -14482 3475
rect -14420 4445 -14386 4464
rect -14420 4373 -14386 4385
rect -14420 4301 -14386 4317
rect -14420 4229 -14386 4249
rect -14420 4157 -14386 4181
rect -14420 4085 -14386 4113
rect -14420 4013 -14386 4045
rect -14420 3943 -14386 3977
rect -14420 3875 -14386 3907
rect -14420 3807 -14386 3835
rect -14420 3739 -14386 3763
rect -14420 3671 -14386 3691
rect -14420 3603 -14386 3619
rect -14420 3535 -14386 3547
rect -14420 3398 -14386 3475
rect -14324 4445 -14290 4506
rect -14324 4373 -14290 4385
rect -14324 4301 -14290 4317
rect -14324 4229 -14290 4249
rect -14324 4157 -14290 4181
rect -14324 4085 -14290 4113
rect -14324 4013 -14290 4045
rect -14324 3943 -14290 3977
rect -14324 3875 -14290 3907
rect -14324 3807 -14290 3835
rect -14324 3739 -14290 3763
rect -14324 3671 -14290 3691
rect -14324 3603 -14290 3619
rect -14324 3535 -14290 3547
rect -14324 3456 -14290 3475
rect -14228 4445 -14194 4464
rect -14228 4373 -14194 4385
rect -14228 4301 -14194 4317
rect -14228 4229 -14194 4249
rect -14228 4157 -14194 4181
rect -14228 4085 -14194 4113
rect -14228 4013 -14194 4045
rect -14228 3943 -14194 3977
rect -14228 3875 -14194 3907
rect -14228 3807 -14194 3835
rect -14228 3739 -14194 3763
rect -14228 3671 -14194 3691
rect -14228 3603 -14194 3619
rect -14228 3535 -14194 3547
rect -14228 3398 -14194 3475
rect -14132 4445 -14098 4506
rect -14132 4373 -14098 4385
rect -14132 4301 -14098 4317
rect -14132 4229 -14098 4249
rect -14132 4157 -14098 4181
rect -14132 4085 -14098 4113
rect -14132 4013 -14098 4045
rect -14132 3943 -14098 3977
rect -14132 3875 -14098 3907
rect -14132 3807 -14098 3835
rect -14132 3739 -14098 3763
rect -14132 3671 -14098 3691
rect -14132 3603 -14098 3619
rect -14132 3535 -14098 3547
rect -14132 3456 -14098 3475
rect -14036 4445 -14002 4464
rect -14036 4373 -14002 4385
rect -14036 4301 -14002 4317
rect -14036 4229 -14002 4249
rect -14036 4157 -14002 4181
rect -14036 4085 -14002 4113
rect -14036 4013 -14002 4045
rect -14036 3943 -14002 3977
rect -14036 3875 -14002 3907
rect -14036 3807 -14002 3835
rect -14036 3739 -14002 3763
rect -14036 3671 -14002 3691
rect -14036 3603 -14002 3619
rect -14036 3535 -14002 3547
rect -14036 3398 -14002 3475
rect -13940 4445 -13906 4506
rect -13940 4373 -13906 4385
rect -13940 4301 -13906 4317
rect -13940 4229 -13906 4249
rect -13940 4157 -13906 4181
rect -13940 4085 -13906 4113
rect -13940 4013 -13906 4045
rect -13940 3943 -13906 3977
rect -13940 3875 -13906 3907
rect -13940 3807 -13906 3835
rect -13940 3739 -13906 3763
rect -13940 3671 -13906 3691
rect -13940 3603 -13906 3619
rect -13940 3535 -13906 3547
rect -13940 3456 -13906 3475
rect -13844 4445 -13810 4464
rect -13844 4373 -13810 4385
rect -13844 4301 -13810 4317
rect -13844 4229 -13810 4249
rect -13844 4157 -13810 4181
rect -13844 4085 -13810 4113
rect -13844 4013 -13810 4045
rect -13844 3943 -13810 3977
rect -13844 3875 -13810 3907
rect -13844 3807 -13810 3835
rect -13844 3739 -13810 3763
rect -13844 3671 -13810 3691
rect -13844 3603 -13810 3619
rect -13844 3535 -13810 3547
rect -13844 3398 -13810 3475
rect -13748 4445 -13714 4506
rect -13748 4373 -13714 4385
rect -13748 4301 -13714 4317
rect -13748 4229 -13714 4249
rect -13748 4157 -13714 4181
rect -13748 4085 -13714 4113
rect -13748 4013 -13714 4045
rect -13748 3943 -13714 3977
rect -13748 3875 -13714 3907
rect -13748 3807 -13714 3835
rect -13748 3739 -13714 3763
rect -13748 3671 -13714 3691
rect -13748 3603 -13714 3619
rect -13748 3535 -13714 3547
rect -13748 3456 -13714 3475
rect -13652 4445 -13618 4464
rect -13652 4373 -13618 4385
rect -13652 4301 -13618 4317
rect -13652 4229 -13618 4249
rect -13652 4157 -13618 4181
rect -13652 4085 -13618 4113
rect -13652 4013 -13618 4045
rect -13652 3943 -13618 3977
rect -13652 3875 -13618 3907
rect -13652 3807 -13618 3835
rect -13652 3739 -13618 3763
rect -13652 3671 -13618 3691
rect -13652 3603 -13618 3619
rect -13652 3535 -13618 3547
rect -13652 3398 -13618 3475
rect -13556 4445 -13522 4506
rect -13556 4373 -13522 4385
rect -13556 4301 -13522 4317
rect -13556 4229 -13522 4249
rect -13556 4157 -13522 4181
rect -13556 4085 -13522 4113
rect -13556 4013 -13522 4045
rect -13556 3943 -13522 3977
rect -13556 3875 -13522 3907
rect -13556 3807 -13522 3835
rect -13556 3739 -13522 3763
rect -13556 3671 -13522 3691
rect -13556 3603 -13522 3619
rect -13556 3535 -13522 3547
rect -13556 3456 -13522 3475
rect -13460 4445 -13426 4464
rect -13460 4373 -13426 4385
rect -13460 4301 -13426 4317
rect -13460 4229 -13426 4249
rect -13460 4157 -13426 4181
rect -13460 4085 -13426 4113
rect -13460 4013 -13426 4045
rect -13460 3943 -13426 3977
rect -13460 3875 -13426 3907
rect -13460 3807 -13426 3835
rect -13460 3739 -13426 3763
rect -13460 3671 -13426 3691
rect -13460 3603 -13426 3619
rect -13460 3535 -13426 3547
rect -13460 3398 -13426 3475
rect -13364 4445 -13330 4506
rect -13364 4373 -13330 4385
rect -13364 4301 -13330 4317
rect -13364 4229 -13330 4249
rect -13364 4157 -13330 4181
rect -13364 4085 -13330 4113
rect -13364 4013 -13330 4045
rect -13364 3943 -13330 3977
rect -13364 3875 -13330 3907
rect -13364 3807 -13330 3835
rect -13364 3739 -13330 3763
rect -13364 3671 -13330 3691
rect -13364 3603 -13330 3619
rect -13364 3535 -13330 3547
rect -13364 3456 -13330 3475
rect -13268 4445 -13234 4464
rect -13268 4373 -13234 4385
rect -13268 4301 -13234 4317
rect -13268 4229 -13234 4249
rect -13268 4157 -13234 4181
rect -13268 4085 -13234 4113
rect -13268 4013 -13234 4045
rect -13268 3943 -13234 3977
rect -13268 3875 -13234 3907
rect -13268 3807 -13234 3835
rect -13268 3739 -13234 3763
rect -13268 3671 -13234 3691
rect -13268 3603 -13234 3619
rect -13268 3535 -13234 3547
rect -13268 3398 -13234 3475
rect -13172 4445 -13138 4506
rect -13172 4373 -13138 4385
rect -13172 4301 -13138 4317
rect -13172 4229 -13138 4249
rect -13172 4157 -13138 4181
rect -13172 4085 -13138 4113
rect -13172 4013 -13138 4045
rect -13172 3943 -13138 3977
rect -13172 3875 -13138 3907
rect -13172 3807 -13138 3835
rect -13172 3739 -13138 3763
rect -13172 3671 -13138 3691
rect -13172 3603 -13138 3619
rect -13172 3535 -13138 3547
rect -13172 3456 -13138 3475
rect -12928 4510 -11934 4524
rect -12928 4451 -12894 4510
rect -12928 4379 -12894 4391
rect -12928 4307 -12894 4323
rect -12928 4235 -12894 4255
rect -12928 4163 -12894 4187
rect -12928 4091 -12894 4119
rect -12928 4019 -12894 4051
rect -12928 3949 -12894 3983
rect -12928 3881 -12894 3913
rect -12928 3813 -12894 3841
rect -12928 3745 -12894 3769
rect -12928 3677 -12894 3697
rect -12928 3609 -12894 3625
rect -12928 3541 -12894 3553
rect -12928 3462 -12894 3481
rect -12832 4451 -12798 4470
rect -12832 4379 -12798 4391
rect -12832 4307 -12798 4323
rect -12832 4235 -12798 4255
rect -12832 4163 -12798 4187
rect -12832 4091 -12798 4119
rect -12832 4019 -12798 4051
rect -12832 3949 -12798 3983
rect -12832 3881 -12798 3913
rect -12832 3813 -12798 3841
rect -12832 3745 -12798 3769
rect -12832 3677 -12798 3697
rect -12832 3609 -12798 3625
rect -12832 3541 -12798 3553
rect -21730 3241 -21714 3275
rect -21680 3241 -21664 3275
rect -22980 3096 -22974 3130
rect -22940 3096 -22934 3130
rect -22980 2930 -22934 3096
rect -20774 3132 -20734 3352
rect -20066 3247 -20050 3281
rect -20016 3247 -20000 3281
rect -20774 3098 -20771 3132
rect -20737 3098 -20734 3132
rect -21732 2982 -21716 3016
rect -21682 2982 -21666 3016
rect -20774 2934 -20734 3098
rect -19120 3145 -19082 3358
rect -18862 3253 -18846 3287
rect -18812 3253 -18796 3287
rect -19120 3111 -19118 3145
rect -19084 3111 -19082 3145
rect -20064 2984 -20048 3018
rect -20014 2984 -19998 3018
rect -19120 2942 -19082 3111
rect -18302 3147 -18268 3366
rect -18174 3235 -18158 3269
rect -18124 3235 -18108 3269
rect -18866 3028 -18850 3062
rect -18816 3028 -18800 3062
rect -23398 2896 -21634 2930
rect -23492 2839 -23458 2858
rect -23492 2767 -23458 2779
rect -23492 2695 -23458 2711
rect -23492 2623 -23458 2643
rect -23492 2551 -23458 2575
rect -23492 2479 -23458 2507
rect -23492 2407 -23458 2439
rect -23492 2337 -23458 2371
rect -23492 2269 -23458 2301
rect -23492 2201 -23458 2229
rect -23492 2133 -23458 2157
rect -23492 2065 -23458 2085
rect -23492 1997 -23458 2013
rect -23492 1929 -23458 1941
rect -23492 1808 -23458 1869
rect -23396 2839 -23362 2896
rect -23396 2767 -23362 2779
rect -23396 2695 -23362 2711
rect -23396 2623 -23362 2643
rect -23396 2551 -23362 2575
rect -23396 2479 -23362 2507
rect -23396 2407 -23362 2439
rect -23396 2337 -23362 2371
rect -23396 2269 -23362 2301
rect -23396 2201 -23362 2229
rect -23396 2133 -23362 2157
rect -23396 2065 -23362 2085
rect -23396 1997 -23362 2013
rect -23396 1929 -23362 1941
rect -23396 1850 -23362 1869
rect -23300 2839 -23266 2858
rect -23300 2767 -23266 2779
rect -23300 2695 -23266 2711
rect -23300 2623 -23266 2643
rect -23300 2551 -23266 2575
rect -23300 2479 -23266 2507
rect -23300 2407 -23266 2439
rect -23300 2337 -23266 2371
rect -23300 2269 -23266 2301
rect -23300 2201 -23266 2229
rect -23300 2133 -23266 2157
rect -23300 2065 -23266 2085
rect -23300 1997 -23266 2013
rect -23300 1929 -23266 1941
rect -23300 1808 -23266 1869
rect -23204 2839 -23170 2896
rect -23204 2767 -23170 2779
rect -23204 2695 -23170 2711
rect -23204 2623 -23170 2643
rect -23204 2551 -23170 2575
rect -23204 2479 -23170 2507
rect -23204 2407 -23170 2439
rect -23204 2337 -23170 2371
rect -23204 2269 -23170 2301
rect -23204 2201 -23170 2229
rect -23204 2133 -23170 2157
rect -23204 2065 -23170 2085
rect -23204 1997 -23170 2013
rect -23204 1929 -23170 1941
rect -23204 1850 -23170 1869
rect -23108 2839 -23074 2858
rect -23108 2767 -23074 2779
rect -23108 2695 -23074 2711
rect -23108 2623 -23074 2643
rect -23108 2551 -23074 2575
rect -23108 2479 -23074 2507
rect -23108 2407 -23074 2439
rect -23108 2337 -23074 2371
rect -23108 2269 -23074 2301
rect -23108 2201 -23074 2229
rect -23108 2133 -23074 2157
rect -23108 2065 -23074 2085
rect -23108 1997 -23074 2013
rect -23108 1929 -23074 1941
rect -23108 1808 -23074 1869
rect -23012 2839 -22978 2896
rect -23012 2767 -22978 2779
rect -23012 2695 -22978 2711
rect -23012 2623 -22978 2643
rect -23012 2551 -22978 2575
rect -23012 2479 -22978 2507
rect -23012 2407 -22978 2439
rect -23012 2337 -22978 2371
rect -23012 2269 -22978 2301
rect -23012 2201 -22978 2229
rect -23012 2133 -22978 2157
rect -23012 2065 -22978 2085
rect -23012 1997 -22978 2013
rect -23012 1929 -22978 1941
rect -23012 1850 -22978 1869
rect -22916 2839 -22882 2858
rect -22916 2767 -22882 2779
rect -22916 2695 -22882 2711
rect -22916 2623 -22882 2643
rect -22916 2551 -22882 2575
rect -22916 2479 -22882 2507
rect -22916 2407 -22882 2439
rect -22916 2337 -22882 2371
rect -22916 2269 -22882 2301
rect -22916 2201 -22882 2229
rect -22916 2133 -22882 2157
rect -22916 2065 -22882 2085
rect -22916 1997 -22882 2013
rect -22916 1929 -22882 1941
rect -22916 1808 -22882 1869
rect -22820 2839 -22786 2896
rect -22820 2767 -22786 2779
rect -22820 2695 -22786 2711
rect -22820 2623 -22786 2643
rect -22820 2551 -22786 2575
rect -22820 2479 -22786 2507
rect -22820 2407 -22786 2439
rect -22820 2337 -22786 2371
rect -22820 2269 -22786 2301
rect -22820 2201 -22786 2229
rect -22820 2133 -22786 2157
rect -22820 2065 -22786 2085
rect -22820 1997 -22786 2013
rect -22820 1929 -22786 1941
rect -22820 1850 -22786 1869
rect -22724 2839 -22690 2858
rect -22724 2767 -22690 2779
rect -22724 2695 -22690 2711
rect -22724 2623 -22690 2643
rect -22724 2551 -22690 2575
rect -22724 2479 -22690 2507
rect -22724 2407 -22690 2439
rect -22724 2337 -22690 2371
rect -22724 2269 -22690 2301
rect -22724 2201 -22690 2229
rect -22724 2133 -22690 2157
rect -22724 2065 -22690 2085
rect -22724 1997 -22690 2013
rect -22724 1929 -22690 1941
rect -22724 1808 -22690 1869
rect -22628 2839 -22594 2896
rect -22628 2767 -22594 2779
rect -22628 2695 -22594 2711
rect -22628 2623 -22594 2643
rect -22628 2551 -22594 2575
rect -22628 2479 -22594 2507
rect -22628 2407 -22594 2439
rect -22628 2337 -22594 2371
rect -22628 2269 -22594 2301
rect -22628 2201 -22594 2229
rect -22628 2133 -22594 2157
rect -22628 2065 -22594 2085
rect -22628 1997 -22594 2013
rect -22628 1929 -22594 1941
rect -22628 1850 -22594 1869
rect -22532 2839 -22498 2858
rect -22532 2767 -22498 2779
rect -22532 2695 -22498 2711
rect -22532 2623 -22498 2643
rect -22532 2551 -22498 2575
rect -22532 2479 -22498 2507
rect -22532 2407 -22498 2439
rect -22532 2337 -22498 2371
rect -22532 2269 -22498 2301
rect -22532 2201 -22498 2229
rect -22532 2133 -22498 2157
rect -22532 2065 -22498 2085
rect -22532 1997 -22498 2013
rect -22532 1929 -22498 1941
rect -22532 1808 -22498 1869
rect -22436 2839 -22402 2896
rect -22436 2767 -22402 2779
rect -22436 2695 -22402 2711
rect -22436 2623 -22402 2643
rect -22436 2551 -22402 2575
rect -22436 2479 -22402 2507
rect -22436 2407 -22402 2439
rect -22436 2337 -22402 2371
rect -22436 2269 -22402 2301
rect -22436 2201 -22402 2229
rect -22436 2133 -22402 2157
rect -22436 2065 -22402 2085
rect -22436 1997 -22402 2013
rect -22436 1929 -22402 1941
rect -22436 1850 -22402 1869
rect -22340 2839 -22306 2858
rect -22340 2767 -22306 2779
rect -22340 2695 -22306 2711
rect -22340 2623 -22306 2643
rect -22340 2551 -22306 2575
rect -22340 2479 -22306 2507
rect -22340 2407 -22306 2439
rect -22340 2337 -22306 2371
rect -22340 2269 -22306 2301
rect -22340 2201 -22306 2229
rect -22340 2133 -22306 2157
rect -22340 2065 -22306 2085
rect -22340 1997 -22306 2013
rect -22340 1929 -22306 1941
rect -22340 1808 -22306 1869
rect -22244 2839 -22210 2896
rect -22244 2767 -22210 2779
rect -22244 2695 -22210 2711
rect -22244 2623 -22210 2643
rect -22244 2551 -22210 2575
rect -22244 2479 -22210 2507
rect -22244 2407 -22210 2439
rect -22244 2337 -22210 2371
rect -22244 2269 -22210 2301
rect -22244 2201 -22210 2229
rect -22244 2133 -22210 2157
rect -22244 2065 -22210 2085
rect -22244 1997 -22210 2013
rect -22244 1929 -22210 1941
rect -22244 1850 -22210 1869
rect -22148 2839 -22114 2858
rect -22148 2767 -22114 2779
rect -22148 2695 -22114 2711
rect -22148 2623 -22114 2643
rect -22148 2551 -22114 2575
rect -22148 2479 -22114 2507
rect -22148 2407 -22114 2439
rect -22148 2337 -22114 2371
rect -22148 2269 -22114 2301
rect -22148 2201 -22114 2229
rect -22148 2133 -22114 2157
rect -22148 2065 -22114 2085
rect -22148 1997 -22114 2013
rect -22148 1929 -22114 1941
rect -22148 1808 -22114 1869
rect -22052 2839 -22018 2896
rect -22052 2767 -22018 2779
rect -22052 2695 -22018 2711
rect -22052 2623 -22018 2643
rect -22052 2551 -22018 2575
rect -22052 2479 -22018 2507
rect -22052 2407 -22018 2439
rect -22052 2337 -22018 2371
rect -22052 2269 -22018 2301
rect -22052 2201 -22018 2229
rect -22052 2133 -22018 2157
rect -22052 2065 -22018 2085
rect -22052 1997 -22018 2013
rect -22052 1929 -22018 1941
rect -22052 1850 -22018 1869
rect -21956 2839 -21922 2858
rect -21956 2767 -21922 2779
rect -21956 2695 -21922 2711
rect -21956 2623 -21922 2643
rect -21956 2551 -21922 2575
rect -21956 2479 -21922 2507
rect -21956 2407 -21922 2439
rect -21956 2337 -21922 2371
rect -21956 2269 -21922 2301
rect -21956 2201 -21922 2229
rect -21956 2133 -21922 2157
rect -21956 2065 -21922 2085
rect -21956 1997 -21922 2013
rect -21956 1929 -21922 1941
rect -21956 1808 -21922 1869
rect -21860 2839 -21826 2896
rect -21860 2767 -21826 2779
rect -21860 2695 -21826 2711
rect -21860 2623 -21826 2643
rect -21860 2551 -21826 2575
rect -21860 2479 -21826 2507
rect -21860 2407 -21826 2439
rect -21860 2337 -21826 2371
rect -21860 2269 -21826 2301
rect -21860 2201 -21826 2229
rect -21860 2133 -21826 2157
rect -21860 2065 -21826 2085
rect -21860 1997 -21826 2013
rect -21860 1929 -21826 1941
rect -21860 1850 -21826 1869
rect -21764 2839 -21730 2858
rect -21764 2767 -21730 2779
rect -21764 2695 -21730 2711
rect -21764 2623 -21730 2643
rect -21764 2551 -21730 2575
rect -21764 2479 -21730 2507
rect -21764 2407 -21730 2439
rect -21764 2337 -21730 2371
rect -21764 2269 -21730 2301
rect -21764 2201 -21730 2229
rect -21764 2133 -21730 2157
rect -21764 2065 -21730 2085
rect -21764 1997 -21730 2013
rect -21764 1929 -21730 1941
rect -21764 1808 -21730 1869
rect -21668 2839 -21634 2896
rect -21344 2900 -19966 2934
rect -21668 2767 -21634 2779
rect -21668 2695 -21634 2711
rect -21668 2623 -21634 2643
rect -21668 2551 -21634 2575
rect -21668 2479 -21634 2507
rect -21668 2407 -21634 2439
rect -21668 2337 -21634 2371
rect -21668 2269 -21634 2301
rect -21668 2201 -21634 2229
rect -21668 2133 -21634 2157
rect -21668 2065 -21634 2085
rect -21668 1997 -21634 2013
rect -21668 1929 -21634 1941
rect -21668 1850 -21634 1869
rect -21572 2839 -21538 2858
rect -21572 2767 -21538 2779
rect -21572 2695 -21538 2711
rect -21572 2623 -21538 2643
rect -21572 2551 -21538 2575
rect -21572 2479 -21538 2507
rect -21572 2407 -21538 2439
rect -21572 2337 -21538 2371
rect -21572 2269 -21538 2301
rect -21572 2201 -21538 2229
rect -21572 2133 -21538 2157
rect -21572 2065 -21538 2085
rect -21572 1997 -21538 2013
rect -21572 1929 -21538 1941
rect -21572 1808 -21538 1869
rect -21344 2831 -21310 2900
rect -21344 2759 -21310 2771
rect -21344 2687 -21310 2703
rect -21344 2615 -21310 2635
rect -21344 2543 -21310 2567
rect -21344 2471 -21310 2499
rect -21344 2399 -21310 2431
rect -21344 2329 -21310 2363
rect -21344 2261 -21310 2293
rect -21344 2193 -21310 2221
rect -21344 2125 -21310 2149
rect -21344 2057 -21310 2077
rect -21344 1989 -21310 2005
rect -21344 1921 -21310 1933
rect -21344 1842 -21310 1861
rect -21248 2831 -21214 2850
rect -21248 2759 -21214 2771
rect -21248 2687 -21214 2703
rect -21248 2615 -21214 2635
rect -21248 2543 -21214 2567
rect -21248 2471 -21214 2499
rect -21248 2399 -21214 2431
rect -21248 2329 -21214 2363
rect -21248 2261 -21214 2293
rect -21248 2193 -21214 2221
rect -21248 2125 -21214 2149
rect -21248 2057 -21214 2077
rect -21248 1989 -21214 2005
rect -21248 1921 -21214 1933
rect -23492 1790 -21538 1808
rect -21248 1800 -21214 1861
rect -21152 2831 -21118 2900
rect -21152 2759 -21118 2771
rect -21152 2687 -21118 2703
rect -21152 2615 -21118 2635
rect -21152 2543 -21118 2567
rect -21152 2471 -21118 2499
rect -21152 2399 -21118 2431
rect -21152 2329 -21118 2363
rect -21152 2261 -21118 2293
rect -21152 2193 -21118 2221
rect -21152 2125 -21118 2149
rect -21152 2057 -21118 2077
rect -21152 1989 -21118 2005
rect -21152 1921 -21118 1933
rect -21152 1842 -21118 1861
rect -21056 2831 -21022 2850
rect -21056 2759 -21022 2771
rect -21056 2687 -21022 2703
rect -21056 2615 -21022 2635
rect -21056 2543 -21022 2567
rect -21056 2471 -21022 2499
rect -21056 2399 -21022 2431
rect -21056 2329 -21022 2363
rect -21056 2261 -21022 2293
rect -21056 2193 -21022 2221
rect -21056 2125 -21022 2149
rect -21056 2057 -21022 2077
rect -21056 1989 -21022 2005
rect -21056 1921 -21022 1933
rect -21056 1800 -21022 1861
rect -20960 2831 -20926 2900
rect -20960 2759 -20926 2771
rect -20960 2687 -20926 2703
rect -20960 2615 -20926 2635
rect -20960 2543 -20926 2567
rect -20960 2471 -20926 2499
rect -20960 2399 -20926 2431
rect -20960 2329 -20926 2363
rect -20960 2261 -20926 2293
rect -20960 2193 -20926 2221
rect -20960 2125 -20926 2149
rect -20960 2057 -20926 2077
rect -20960 1989 -20926 2005
rect -20960 1921 -20926 1933
rect -20960 1842 -20926 1861
rect -20864 2831 -20830 2850
rect -20864 2759 -20830 2771
rect -20864 2687 -20830 2703
rect -20864 2615 -20830 2635
rect -20864 2543 -20830 2567
rect -20864 2471 -20830 2499
rect -20864 2399 -20830 2431
rect -20864 2329 -20830 2363
rect -20864 2261 -20830 2293
rect -20864 2193 -20830 2221
rect -20864 2125 -20830 2149
rect -20864 2057 -20830 2077
rect -20864 1989 -20830 2005
rect -20864 1921 -20830 1933
rect -20864 1800 -20830 1861
rect -20768 2831 -20734 2900
rect -20768 2759 -20734 2771
rect -20768 2687 -20734 2703
rect -20768 2615 -20734 2635
rect -20768 2543 -20734 2567
rect -20768 2471 -20734 2499
rect -20768 2399 -20734 2431
rect -20768 2329 -20734 2363
rect -20768 2261 -20734 2293
rect -20768 2193 -20734 2221
rect -20768 2125 -20734 2149
rect -20768 2057 -20734 2077
rect -20768 1989 -20734 2005
rect -20768 1921 -20734 1933
rect -20768 1842 -20734 1861
rect -20672 2831 -20638 2850
rect -20672 2759 -20638 2771
rect -20672 2687 -20638 2703
rect -20672 2615 -20638 2635
rect -20672 2543 -20638 2567
rect -20672 2471 -20638 2499
rect -20672 2399 -20638 2431
rect -20672 2329 -20638 2363
rect -20672 2261 -20638 2293
rect -20672 2193 -20638 2221
rect -20672 2125 -20638 2149
rect -20672 2057 -20638 2077
rect -20672 1989 -20638 2005
rect -20672 1921 -20638 1933
rect -20672 1800 -20638 1861
rect -20576 2831 -20542 2900
rect -20576 2759 -20542 2771
rect -20576 2687 -20542 2703
rect -20576 2615 -20542 2635
rect -20576 2543 -20542 2567
rect -20576 2471 -20542 2499
rect -20576 2399 -20542 2431
rect -20576 2329 -20542 2363
rect -20576 2261 -20542 2293
rect -20576 2193 -20542 2221
rect -20576 2125 -20542 2149
rect -20576 2057 -20542 2077
rect -20576 1989 -20542 2005
rect -20576 1921 -20542 1933
rect -20576 1842 -20542 1861
rect -20480 2831 -20446 2850
rect -20480 2759 -20446 2771
rect -20480 2687 -20446 2703
rect -20480 2615 -20446 2635
rect -20480 2543 -20446 2567
rect -20480 2471 -20446 2499
rect -20480 2399 -20446 2431
rect -20480 2329 -20446 2363
rect -20480 2261 -20446 2293
rect -20480 2193 -20446 2221
rect -20480 2125 -20446 2149
rect -20480 2057 -20446 2077
rect -20480 1989 -20446 2005
rect -20480 1921 -20446 1933
rect -20480 1800 -20446 1861
rect -20384 2831 -20350 2900
rect -20384 2759 -20350 2771
rect -20384 2687 -20350 2703
rect -20384 2615 -20350 2635
rect -20384 2543 -20350 2567
rect -20384 2471 -20350 2499
rect -20384 2399 -20350 2431
rect -20384 2329 -20350 2363
rect -20384 2261 -20350 2293
rect -20384 2193 -20350 2221
rect -20384 2125 -20350 2149
rect -20384 2057 -20350 2077
rect -20384 1989 -20350 2005
rect -20384 1921 -20350 1933
rect -20384 1842 -20350 1861
rect -20288 2831 -20254 2850
rect -20288 2759 -20254 2771
rect -20288 2687 -20254 2703
rect -20288 2615 -20254 2635
rect -20288 2543 -20254 2567
rect -20288 2471 -20254 2499
rect -20288 2399 -20254 2431
rect -20288 2329 -20254 2363
rect -20288 2261 -20254 2293
rect -20288 2193 -20254 2221
rect -20288 2125 -20254 2149
rect -20288 2057 -20254 2077
rect -20288 1989 -20254 2005
rect -20288 1921 -20254 1933
rect -20288 1800 -20254 1861
rect -20192 2831 -20158 2900
rect -20192 2759 -20158 2771
rect -20192 2687 -20158 2703
rect -20192 2615 -20158 2635
rect -20192 2543 -20158 2567
rect -20192 2471 -20158 2499
rect -20192 2399 -20158 2431
rect -20192 2329 -20158 2363
rect -20192 2261 -20158 2293
rect -20192 2193 -20158 2221
rect -20192 2125 -20158 2149
rect -20192 2057 -20158 2077
rect -20192 1989 -20158 2005
rect -20192 1921 -20158 1933
rect -20192 1842 -20158 1861
rect -20096 2831 -20062 2850
rect -20096 2759 -20062 2771
rect -20096 2687 -20062 2703
rect -20096 2615 -20062 2635
rect -20096 2543 -20062 2567
rect -20096 2471 -20062 2499
rect -20096 2399 -20062 2431
rect -20096 2329 -20062 2363
rect -20096 2261 -20062 2293
rect -20096 2193 -20062 2221
rect -20096 2125 -20062 2149
rect -20096 2057 -20062 2077
rect -20096 1989 -20062 2005
rect -20096 1921 -20062 1933
rect -20096 1800 -20062 1861
rect -20000 2831 -19966 2900
rect -19570 2908 -18768 2942
rect -18302 2932 -18268 3113
rect -16150 3142 -16104 3370
rect -14612 3364 -13234 3398
rect -12832 3404 -12798 3481
rect -12736 4451 -12702 4510
rect -12736 4379 -12702 4391
rect -12736 4307 -12702 4323
rect -12736 4235 -12702 4255
rect -12736 4163 -12702 4187
rect -12736 4091 -12702 4119
rect -12736 4019 -12702 4051
rect -12736 3949 -12702 3983
rect -12736 3881 -12702 3913
rect -12736 3813 -12702 3841
rect -12736 3745 -12702 3769
rect -12736 3677 -12702 3697
rect -12736 3609 -12702 3625
rect -12736 3541 -12702 3553
rect -12736 3462 -12702 3481
rect -12640 4451 -12606 4470
rect -12640 4379 -12606 4391
rect -12640 4307 -12606 4323
rect -12640 4235 -12606 4255
rect -12640 4163 -12606 4187
rect -12640 4091 -12606 4119
rect -12640 4019 -12606 4051
rect -12640 3949 -12606 3983
rect -12640 3881 -12606 3913
rect -12640 3813 -12606 3841
rect -12640 3745 -12606 3769
rect -12640 3677 -12606 3697
rect -12640 3609 -12606 3625
rect -12640 3541 -12606 3553
rect -12640 3404 -12606 3481
rect -12544 4451 -12510 4510
rect -12544 4379 -12510 4391
rect -12544 4307 -12510 4323
rect -12544 4235 -12510 4255
rect -12544 4163 -12510 4187
rect -12544 4091 -12510 4119
rect -12544 4019 -12510 4051
rect -12544 3949 -12510 3983
rect -12544 3881 -12510 3913
rect -12544 3813 -12510 3841
rect -12544 3745 -12510 3769
rect -12544 3677 -12510 3697
rect -12544 3609 -12510 3625
rect -12544 3541 -12510 3553
rect -12544 3462 -12510 3481
rect -12448 4451 -12414 4470
rect -12448 4379 -12414 4391
rect -12448 4307 -12414 4323
rect -12448 4235 -12414 4255
rect -12448 4163 -12414 4187
rect -12448 4091 -12414 4119
rect -12448 4019 -12414 4051
rect -12448 3949 -12414 3983
rect -12448 3881 -12414 3913
rect -12448 3813 -12414 3841
rect -12448 3745 -12414 3769
rect -12448 3677 -12414 3697
rect -12448 3609 -12414 3625
rect -12448 3541 -12414 3553
rect -12448 3404 -12414 3481
rect -12352 4451 -12318 4510
rect -12352 4379 -12318 4391
rect -12352 4307 -12318 4323
rect -12352 4235 -12318 4255
rect -12352 4163 -12318 4187
rect -12352 4091 -12318 4119
rect -12352 4019 -12318 4051
rect -12352 3949 -12318 3983
rect -12352 3881 -12318 3913
rect -12352 3813 -12318 3841
rect -12352 3745 -12318 3769
rect -12352 3677 -12318 3697
rect -12352 3609 -12318 3625
rect -12352 3541 -12318 3553
rect -12352 3462 -12318 3481
rect -12256 4451 -12222 4470
rect -12256 4379 -12222 4391
rect -12256 4307 -12222 4323
rect -12256 4235 -12222 4255
rect -12256 4163 -12222 4187
rect -12256 4091 -12222 4119
rect -12256 4019 -12222 4051
rect -12256 3949 -12222 3983
rect -12256 3881 -12222 3913
rect -12256 3813 -12222 3841
rect -12256 3745 -12222 3769
rect -12256 3677 -12222 3697
rect -12256 3609 -12222 3625
rect -12256 3541 -12222 3553
rect -12256 3404 -12222 3481
rect -12160 4451 -12126 4510
rect -12160 4379 -12126 4391
rect -12160 4307 -12126 4323
rect -12160 4235 -12126 4255
rect -12160 4163 -12126 4187
rect -12160 4091 -12126 4119
rect -12160 4019 -12126 4051
rect -12160 3949 -12126 3983
rect -12160 3881 -12126 3913
rect -12160 3813 -12126 3841
rect -12160 3745 -12126 3769
rect -12160 3677 -12126 3697
rect -12160 3609 -12126 3625
rect -12160 3541 -12126 3553
rect -12160 3462 -12126 3481
rect -12064 4451 -12030 4470
rect -12064 4379 -12030 4391
rect -12064 4307 -12030 4323
rect -12064 4235 -12030 4255
rect -12064 4163 -12030 4187
rect -12064 4091 -12030 4119
rect -12064 4019 -12030 4051
rect -12064 3949 -12030 3983
rect -12064 3881 -12030 3913
rect -12064 3813 -12030 3841
rect -12064 3745 -12030 3769
rect -12064 3677 -12030 3697
rect -12064 3609 -12030 3625
rect -12064 3541 -12030 3553
rect -12064 3404 -12030 3481
rect -11968 4451 -11934 4510
rect -11664 4512 -11246 4524
rect -11968 4379 -11934 4391
rect -11968 4307 -11934 4323
rect -11968 4235 -11934 4255
rect -11968 4163 -11934 4187
rect -11968 4091 -11934 4119
rect -11968 4019 -11934 4051
rect -11968 3949 -11934 3983
rect -11968 3881 -11934 3913
rect -11968 3813 -11934 3841
rect -11968 3745 -11934 3769
rect -11968 3677 -11934 3697
rect -11968 3609 -11934 3625
rect -11968 3541 -11934 3553
rect -11968 3462 -11934 3481
rect -11760 4453 -11726 4472
rect -11760 4381 -11726 4393
rect -11760 4309 -11726 4325
rect -11760 4237 -11726 4257
rect -11760 4165 -11726 4189
rect -11760 4093 -11726 4121
rect -11760 4021 -11726 4053
rect -11760 3951 -11726 3985
rect -11760 3883 -11726 3915
rect -11760 3815 -11726 3843
rect -11760 3747 -11726 3771
rect -11760 3679 -11726 3699
rect -11760 3611 -11726 3627
rect -11760 3543 -11726 3555
rect -12832 3370 -12030 3404
rect -11760 3412 -11726 3483
rect -11664 4453 -11630 4512
rect -11664 4381 -11630 4393
rect -11664 4309 -11630 4325
rect -11664 4237 -11630 4257
rect -11664 4165 -11630 4189
rect -11664 4093 -11630 4121
rect -11664 4021 -11630 4053
rect -11664 3951 -11630 3985
rect -11664 3883 -11630 3915
rect -11664 3815 -11630 3843
rect -11664 3747 -11630 3771
rect -11664 3679 -11630 3699
rect -11664 3611 -11630 3627
rect -11664 3543 -11630 3555
rect -11664 3464 -11630 3483
rect -11568 4453 -11534 4472
rect -11568 4381 -11534 4393
rect -11568 4309 -11534 4325
rect -11568 4237 -11534 4257
rect -11568 4165 -11534 4189
rect -11568 4093 -11534 4121
rect -11568 4021 -11534 4053
rect -11568 3951 -11534 3985
rect -11568 3883 -11534 3915
rect -11568 3815 -11534 3843
rect -11568 3747 -11534 3771
rect -11568 3679 -11534 3699
rect -11568 3611 -11534 3627
rect -11568 3543 -11534 3555
rect -11568 3412 -11534 3483
rect -11472 4453 -11438 4512
rect -11472 4381 -11438 4393
rect -11472 4309 -11438 4325
rect -11472 4237 -11438 4257
rect -11472 4165 -11438 4189
rect -11472 4093 -11438 4121
rect -11472 4021 -11438 4053
rect -11472 3951 -11438 3985
rect -11472 3883 -11438 3915
rect -11472 3815 -11438 3843
rect -11472 3747 -11438 3771
rect -11472 3679 -11438 3699
rect -11472 3611 -11438 3627
rect -11472 3543 -11438 3555
rect -11472 3464 -11438 3483
rect -11376 4453 -11342 4472
rect -11376 4381 -11342 4393
rect -11376 4309 -11342 4325
rect -11376 4237 -11342 4257
rect -11376 4165 -11342 4189
rect -11376 4093 -11342 4121
rect -11376 4021 -11342 4053
rect -11376 3951 -11342 3985
rect -11376 3883 -11342 3915
rect -11376 3815 -11342 3843
rect -11376 3747 -11342 3771
rect -11376 3679 -11342 3699
rect -11376 3611 -11342 3627
rect -11376 3543 -11342 3555
rect -11376 3412 -11342 3483
rect -11280 4453 -11246 4512
rect -11280 4381 -11246 4393
rect -11280 4309 -11246 4325
rect -11280 4237 -11246 4257
rect -11280 4165 -11246 4189
rect -11280 4093 -11246 4121
rect -11280 4021 -11246 4053
rect -11280 3951 -11246 3985
rect -11280 3883 -11246 3915
rect -11280 3815 -11246 3843
rect -11280 3747 -11246 3771
rect -11280 3679 -11246 3699
rect -11280 3611 -11246 3627
rect -11280 3543 -11246 3555
rect -11280 3464 -11246 3483
rect -10290 4510 -8336 4532
rect -10290 4437 -10256 4510
rect -10290 4365 -10256 4377
rect -10290 4293 -10256 4309
rect -10290 4221 -10256 4241
rect -10290 4149 -10256 4173
rect -10290 4077 -10256 4105
rect -10290 4005 -10256 4037
rect -10290 3935 -10256 3969
rect -10290 3867 -10256 3899
rect -10290 3799 -10256 3827
rect -10290 3731 -10256 3755
rect -10290 3663 -10256 3683
rect -10290 3595 -10256 3611
rect -10290 3527 -10256 3539
rect -10290 3448 -10256 3467
rect -10194 4437 -10160 4456
rect -10194 4365 -10160 4377
rect -10194 4293 -10160 4309
rect -10194 4221 -10160 4241
rect -10194 4149 -10160 4173
rect -10194 4077 -10160 4105
rect -10194 4005 -10160 4037
rect -10194 3935 -10160 3969
rect -10194 3867 -10160 3899
rect -10194 3799 -10160 3827
rect -10194 3731 -10160 3755
rect -10194 3663 -10160 3683
rect -10194 3595 -10160 3611
rect -10194 3527 -10160 3539
rect -11760 3378 -11340 3412
rect -10194 3402 -10160 3467
rect -10098 4437 -10064 4510
rect -10098 4365 -10064 4377
rect -10098 4293 -10064 4309
rect -10098 4221 -10064 4241
rect -10098 4149 -10064 4173
rect -10098 4077 -10064 4105
rect -10098 4005 -10064 4037
rect -10098 3935 -10064 3969
rect -10098 3867 -10064 3899
rect -10098 3799 -10064 3827
rect -10098 3731 -10064 3755
rect -10098 3663 -10064 3683
rect -10098 3595 -10064 3611
rect -10098 3527 -10064 3539
rect -10098 3448 -10064 3467
rect -10002 4437 -9968 4456
rect -10002 4365 -9968 4377
rect -10002 4293 -9968 4309
rect -10002 4221 -9968 4241
rect -10002 4149 -9968 4173
rect -10002 4077 -9968 4105
rect -10002 4005 -9968 4037
rect -10002 3935 -9968 3969
rect -10002 3867 -9968 3899
rect -10002 3799 -9968 3827
rect -10002 3731 -9968 3755
rect -10002 3663 -9968 3683
rect -10002 3595 -9968 3611
rect -10002 3527 -9968 3539
rect -10002 3402 -9968 3467
rect -9906 4437 -9872 4510
rect -9906 4365 -9872 4377
rect -9906 4293 -9872 4309
rect -9906 4221 -9872 4241
rect -9906 4149 -9872 4173
rect -9906 4077 -9872 4105
rect -9906 4005 -9872 4037
rect -9906 3935 -9872 3969
rect -9906 3867 -9872 3899
rect -9906 3799 -9872 3827
rect -9906 3731 -9872 3755
rect -9906 3663 -9872 3683
rect -9906 3595 -9872 3611
rect -9906 3527 -9872 3539
rect -9906 3448 -9872 3467
rect -9810 4437 -9776 4456
rect -9810 4365 -9776 4377
rect -9810 4293 -9776 4309
rect -9810 4221 -9776 4241
rect -9810 4149 -9776 4173
rect -9810 4077 -9776 4105
rect -9810 4005 -9776 4037
rect -9810 3935 -9776 3969
rect -9810 3867 -9776 3899
rect -9810 3799 -9776 3827
rect -9810 3731 -9776 3755
rect -9810 3663 -9776 3683
rect -9810 3595 -9776 3611
rect -9810 3527 -9776 3539
rect -9810 3402 -9776 3467
rect -9714 4437 -9680 4510
rect -9714 4365 -9680 4377
rect -9714 4293 -9680 4309
rect -9714 4221 -9680 4241
rect -9714 4149 -9680 4173
rect -9714 4077 -9680 4105
rect -9714 4005 -9680 4037
rect -9714 3935 -9680 3969
rect -9714 3867 -9680 3899
rect -9714 3799 -9680 3827
rect -9714 3731 -9680 3755
rect -9714 3663 -9680 3683
rect -9714 3595 -9680 3611
rect -9714 3527 -9680 3539
rect -9714 3448 -9680 3467
rect -9618 4437 -9584 4456
rect -9618 4365 -9584 4377
rect -9618 4293 -9584 4309
rect -9618 4221 -9584 4241
rect -9618 4149 -9584 4173
rect -9618 4077 -9584 4105
rect -9618 4005 -9584 4037
rect -9618 3935 -9584 3969
rect -9618 3867 -9584 3899
rect -9618 3799 -9584 3827
rect -9618 3731 -9584 3755
rect -9618 3663 -9584 3683
rect -9618 3595 -9584 3611
rect -9618 3527 -9584 3539
rect -9618 3402 -9584 3467
rect -9522 4437 -9488 4510
rect -9522 4365 -9488 4377
rect -9522 4293 -9488 4309
rect -9522 4221 -9488 4241
rect -9522 4149 -9488 4173
rect -9522 4077 -9488 4105
rect -9522 4005 -9488 4037
rect -9522 3935 -9488 3969
rect -9522 3867 -9488 3899
rect -9522 3799 -9488 3827
rect -9522 3731 -9488 3755
rect -9522 3663 -9488 3683
rect -9522 3595 -9488 3611
rect -9522 3527 -9488 3539
rect -9522 3448 -9488 3467
rect -9426 4437 -9392 4456
rect -9426 4365 -9392 4377
rect -9426 4293 -9392 4309
rect -9426 4221 -9392 4241
rect -9426 4149 -9392 4173
rect -9426 4077 -9392 4105
rect -9426 4005 -9392 4037
rect -9426 3935 -9392 3969
rect -9426 3867 -9392 3899
rect -9426 3799 -9392 3827
rect -9426 3731 -9392 3755
rect -9426 3663 -9392 3683
rect -9426 3595 -9392 3611
rect -9426 3527 -9392 3539
rect -9426 3402 -9392 3467
rect -9330 4437 -9296 4510
rect -9330 4365 -9296 4377
rect -9330 4293 -9296 4309
rect -9330 4221 -9296 4241
rect -9330 4149 -9296 4173
rect -9330 4077 -9296 4105
rect -9330 4005 -9296 4037
rect -9330 3935 -9296 3969
rect -9330 3867 -9296 3899
rect -9330 3799 -9296 3827
rect -9330 3731 -9296 3755
rect -9330 3663 -9296 3683
rect -9330 3595 -9296 3611
rect -9330 3527 -9296 3539
rect -9330 3448 -9296 3467
rect -9234 4437 -9200 4456
rect -9234 4365 -9200 4377
rect -9234 4293 -9200 4309
rect -9234 4221 -9200 4241
rect -9234 4149 -9200 4173
rect -9234 4077 -9200 4105
rect -9234 4005 -9200 4037
rect -9234 3935 -9200 3969
rect -9234 3867 -9200 3899
rect -9234 3799 -9200 3827
rect -9234 3731 -9200 3755
rect -9234 3663 -9200 3683
rect -9234 3595 -9200 3611
rect -9234 3527 -9200 3539
rect -9234 3402 -9200 3467
rect -9138 4437 -9104 4510
rect -9138 4365 -9104 4377
rect -9138 4293 -9104 4309
rect -9138 4221 -9104 4241
rect -9138 4149 -9104 4173
rect -9138 4077 -9104 4105
rect -9138 4005 -9104 4037
rect -9138 3935 -9104 3969
rect -9138 3867 -9104 3899
rect -9138 3799 -9104 3827
rect -9138 3731 -9104 3755
rect -9138 3663 -9104 3683
rect -9138 3595 -9104 3611
rect -9138 3527 -9104 3539
rect -9138 3448 -9104 3467
rect -9042 4437 -9008 4456
rect -9042 4365 -9008 4377
rect -9042 4293 -9008 4309
rect -9042 4221 -9008 4241
rect -9042 4149 -9008 4173
rect -9042 4077 -9008 4105
rect -9042 4005 -9008 4037
rect -9042 3935 -9008 3969
rect -9042 3867 -9008 3899
rect -9042 3799 -9008 3827
rect -9042 3731 -9008 3755
rect -9042 3663 -9008 3683
rect -9042 3595 -9008 3611
rect -9042 3527 -9008 3539
rect -9042 3402 -9008 3467
rect -8946 4437 -8912 4510
rect -8946 4365 -8912 4377
rect -8946 4293 -8912 4309
rect -8946 4221 -8912 4241
rect -8946 4149 -8912 4173
rect -8946 4077 -8912 4105
rect -8946 4005 -8912 4037
rect -8946 3935 -8912 3969
rect -8946 3867 -8912 3899
rect -8946 3799 -8912 3827
rect -8946 3731 -8912 3755
rect -8946 3663 -8912 3683
rect -8946 3595 -8912 3611
rect -8946 3527 -8912 3539
rect -8946 3448 -8912 3467
rect -8850 4437 -8816 4456
rect -8850 4365 -8816 4377
rect -8850 4293 -8816 4309
rect -8850 4221 -8816 4241
rect -8850 4149 -8816 4173
rect -8850 4077 -8816 4105
rect -8850 4005 -8816 4037
rect -8850 3935 -8816 3969
rect -8850 3867 -8816 3899
rect -8850 3799 -8816 3827
rect -8850 3731 -8816 3755
rect -8850 3663 -8816 3683
rect -8850 3595 -8816 3611
rect -8850 3527 -8816 3539
rect -8850 3402 -8816 3467
rect -8754 4437 -8720 4510
rect -8754 4365 -8720 4377
rect -8754 4293 -8720 4309
rect -8754 4221 -8720 4241
rect -8754 4149 -8720 4173
rect -8754 4077 -8720 4105
rect -8754 4005 -8720 4037
rect -8754 3935 -8720 3969
rect -8754 3867 -8720 3899
rect -8754 3799 -8720 3827
rect -8754 3731 -8720 3755
rect -8754 3663 -8720 3683
rect -8754 3595 -8720 3611
rect -8754 3527 -8720 3539
rect -8754 3448 -8720 3467
rect -8658 4437 -8624 4456
rect -8658 4365 -8624 4377
rect -8658 4293 -8624 4309
rect -8658 4221 -8624 4241
rect -8658 4149 -8624 4173
rect -8658 4077 -8624 4105
rect -8658 4005 -8624 4037
rect -8658 3935 -8624 3969
rect -8658 3867 -8624 3899
rect -8658 3799 -8624 3827
rect -8658 3731 -8624 3755
rect -8658 3663 -8624 3683
rect -8658 3595 -8624 3611
rect -8658 3527 -8624 3539
rect -8658 3402 -8624 3467
rect -8562 4437 -8528 4510
rect -8562 4365 -8528 4377
rect -8562 4293 -8528 4309
rect -8562 4221 -8528 4241
rect -8562 4149 -8528 4173
rect -8562 4077 -8528 4105
rect -8562 4005 -8528 4037
rect -8562 3935 -8528 3969
rect -8562 3867 -8528 3899
rect -8562 3799 -8528 3827
rect -8562 3731 -8528 3755
rect -8562 3663 -8528 3683
rect -8562 3595 -8528 3611
rect -8562 3527 -8528 3539
rect -8562 3448 -8528 3467
rect -8466 4437 -8432 4456
rect -8466 4365 -8432 4377
rect -8466 4293 -8432 4309
rect -8466 4221 -8432 4241
rect -8466 4149 -8432 4173
rect -8466 4077 -8432 4105
rect -8466 4005 -8432 4037
rect -8466 3935 -8432 3969
rect -8466 3867 -8432 3899
rect -8466 3799 -8432 3827
rect -8466 3731 -8432 3755
rect -8466 3663 -8432 3683
rect -8466 3595 -8432 3611
rect -8466 3527 -8432 3539
rect -8466 3402 -8432 3467
rect -8370 4437 -8336 4510
rect -8050 4504 -6672 4532
rect -8370 4365 -8336 4377
rect -8370 4293 -8336 4309
rect -8370 4221 -8336 4241
rect -8370 4149 -8336 4173
rect -8370 4077 -8336 4105
rect -8370 4005 -8336 4037
rect -8370 3935 -8336 3969
rect -8370 3867 -8336 3899
rect -8370 3799 -8336 3827
rect -8370 3731 -8336 3755
rect -8370 3663 -8336 3683
rect -8370 3595 -8336 3611
rect -8370 3527 -8336 3539
rect -8370 3448 -8336 3467
rect -8146 4443 -8112 4462
rect -8146 4371 -8112 4383
rect -8146 4299 -8112 4315
rect -8146 4227 -8112 4247
rect -8146 4155 -8112 4179
rect -8146 4083 -8112 4111
rect -8146 4011 -8112 4043
rect -8146 3941 -8112 3975
rect -8146 3873 -8112 3905
rect -8146 3805 -8112 3833
rect -8146 3737 -8112 3761
rect -8146 3669 -8112 3689
rect -8146 3601 -8112 3617
rect -8146 3533 -8112 3545
rect -14900 3253 -14884 3287
rect -14850 3253 -14834 3287
rect -16150 3108 -16144 3142
rect -16110 3108 -16104 3142
rect -18174 2998 -18158 3032
rect -18124 2998 -18108 3032
rect -16150 2942 -16104 3108
rect -13944 3144 -13904 3364
rect -13236 3259 -13220 3293
rect -13186 3259 -13170 3293
rect -13944 3110 -13941 3144
rect -13907 3110 -13904 3144
rect -14902 2994 -14886 3028
rect -14852 2994 -14836 3028
rect -13944 2946 -13904 3110
rect -12290 3157 -12252 3370
rect -12032 3265 -12016 3299
rect -11982 3265 -11966 3299
rect -12290 3123 -12288 3157
rect -12254 3123 -12252 3157
rect -13234 2996 -13218 3030
rect -13184 2996 -13168 3030
rect -12290 2954 -12252 3123
rect -11472 3159 -11438 3378
rect -10194 3368 -8432 3402
rect -8146 3396 -8112 3473
rect -8050 4443 -8016 4504
rect -8050 4371 -8016 4383
rect -8050 4299 -8016 4315
rect -8050 4227 -8016 4247
rect -8050 4155 -8016 4179
rect -8050 4083 -8016 4111
rect -8050 4011 -8016 4043
rect -8050 3941 -8016 3975
rect -8050 3873 -8016 3905
rect -8050 3805 -8016 3833
rect -8050 3737 -8016 3761
rect -8050 3669 -8016 3689
rect -8050 3601 -8016 3617
rect -8050 3533 -8016 3545
rect -8050 3454 -8016 3473
rect -7954 4443 -7920 4462
rect -7954 4371 -7920 4383
rect -7954 4299 -7920 4315
rect -7954 4227 -7920 4247
rect -7954 4155 -7920 4179
rect -7954 4083 -7920 4111
rect -7954 4011 -7920 4043
rect -7954 3941 -7920 3975
rect -7954 3873 -7920 3905
rect -7954 3805 -7920 3833
rect -7954 3737 -7920 3761
rect -7954 3669 -7920 3689
rect -7954 3601 -7920 3617
rect -7954 3533 -7920 3545
rect -7954 3396 -7920 3473
rect -7858 4443 -7824 4504
rect -7858 4371 -7824 4383
rect -7858 4299 -7824 4315
rect -7858 4227 -7824 4247
rect -7858 4155 -7824 4179
rect -7858 4083 -7824 4111
rect -7858 4011 -7824 4043
rect -7858 3941 -7824 3975
rect -7858 3873 -7824 3905
rect -7858 3805 -7824 3833
rect -7858 3737 -7824 3761
rect -7858 3669 -7824 3689
rect -7858 3601 -7824 3617
rect -7858 3533 -7824 3545
rect -7858 3454 -7824 3473
rect -7762 4443 -7728 4462
rect -7762 4371 -7728 4383
rect -7762 4299 -7728 4315
rect -7762 4227 -7728 4247
rect -7762 4155 -7728 4179
rect -7762 4083 -7728 4111
rect -7762 4011 -7728 4043
rect -7762 3941 -7728 3975
rect -7762 3873 -7728 3905
rect -7762 3805 -7728 3833
rect -7762 3737 -7728 3761
rect -7762 3669 -7728 3689
rect -7762 3601 -7728 3617
rect -7762 3533 -7728 3545
rect -7762 3396 -7728 3473
rect -7666 4443 -7632 4504
rect -7666 4371 -7632 4383
rect -7666 4299 -7632 4315
rect -7666 4227 -7632 4247
rect -7666 4155 -7632 4179
rect -7666 4083 -7632 4111
rect -7666 4011 -7632 4043
rect -7666 3941 -7632 3975
rect -7666 3873 -7632 3905
rect -7666 3805 -7632 3833
rect -7666 3737 -7632 3761
rect -7666 3669 -7632 3689
rect -7666 3601 -7632 3617
rect -7666 3533 -7632 3545
rect -7666 3454 -7632 3473
rect -7570 4443 -7536 4462
rect -7570 4371 -7536 4383
rect -7570 4299 -7536 4315
rect -7570 4227 -7536 4247
rect -7570 4155 -7536 4179
rect -7570 4083 -7536 4111
rect -7570 4011 -7536 4043
rect -7570 3941 -7536 3975
rect -7570 3873 -7536 3905
rect -7570 3805 -7536 3833
rect -7570 3737 -7536 3761
rect -7570 3669 -7536 3689
rect -7570 3601 -7536 3617
rect -7570 3533 -7536 3545
rect -7570 3396 -7536 3473
rect -7474 4443 -7440 4504
rect -7474 4371 -7440 4383
rect -7474 4299 -7440 4315
rect -7474 4227 -7440 4247
rect -7474 4155 -7440 4179
rect -7474 4083 -7440 4111
rect -7474 4011 -7440 4043
rect -7474 3941 -7440 3975
rect -7474 3873 -7440 3905
rect -7474 3805 -7440 3833
rect -7474 3737 -7440 3761
rect -7474 3669 -7440 3689
rect -7474 3601 -7440 3617
rect -7474 3533 -7440 3545
rect -7474 3454 -7440 3473
rect -7378 4443 -7344 4462
rect -7378 4371 -7344 4383
rect -7378 4299 -7344 4315
rect -7378 4227 -7344 4247
rect -7378 4155 -7344 4179
rect -7378 4083 -7344 4111
rect -7378 4011 -7344 4043
rect -7378 3941 -7344 3975
rect -7378 3873 -7344 3905
rect -7378 3805 -7344 3833
rect -7378 3737 -7344 3761
rect -7378 3669 -7344 3689
rect -7378 3601 -7344 3617
rect -7378 3533 -7344 3545
rect -7378 3396 -7344 3473
rect -7282 4443 -7248 4504
rect -7282 4371 -7248 4383
rect -7282 4299 -7248 4315
rect -7282 4227 -7248 4247
rect -7282 4155 -7248 4179
rect -7282 4083 -7248 4111
rect -7282 4011 -7248 4043
rect -7282 3941 -7248 3975
rect -7282 3873 -7248 3905
rect -7282 3805 -7248 3833
rect -7282 3737 -7248 3761
rect -7282 3669 -7248 3689
rect -7282 3601 -7248 3617
rect -7282 3533 -7248 3545
rect -7282 3454 -7248 3473
rect -7186 4443 -7152 4462
rect -7186 4371 -7152 4383
rect -7186 4299 -7152 4315
rect -7186 4227 -7152 4247
rect -7186 4155 -7152 4179
rect -7186 4083 -7152 4111
rect -7186 4011 -7152 4043
rect -7186 3941 -7152 3975
rect -7186 3873 -7152 3905
rect -7186 3805 -7152 3833
rect -7186 3737 -7152 3761
rect -7186 3669 -7152 3689
rect -7186 3601 -7152 3617
rect -7186 3533 -7152 3545
rect -7186 3396 -7152 3473
rect -7090 4443 -7056 4504
rect -7090 4371 -7056 4383
rect -7090 4299 -7056 4315
rect -7090 4227 -7056 4247
rect -7090 4155 -7056 4179
rect -7090 4083 -7056 4111
rect -7090 4011 -7056 4043
rect -7090 3941 -7056 3975
rect -7090 3873 -7056 3905
rect -7090 3805 -7056 3833
rect -7090 3737 -7056 3761
rect -7090 3669 -7056 3689
rect -7090 3601 -7056 3617
rect -7090 3533 -7056 3545
rect -7090 3454 -7056 3473
rect -6994 4443 -6960 4462
rect -6994 4371 -6960 4383
rect -6994 4299 -6960 4315
rect -6994 4227 -6960 4247
rect -6994 4155 -6960 4179
rect -6994 4083 -6960 4111
rect -6994 4011 -6960 4043
rect -6994 3941 -6960 3975
rect -6994 3873 -6960 3905
rect -6994 3805 -6960 3833
rect -6994 3737 -6960 3761
rect -6994 3669 -6960 3689
rect -6994 3601 -6960 3617
rect -6994 3533 -6960 3545
rect -6994 3396 -6960 3473
rect -6898 4443 -6864 4504
rect -6898 4371 -6864 4383
rect -6898 4299 -6864 4315
rect -6898 4227 -6864 4247
rect -6898 4155 -6864 4179
rect -6898 4083 -6864 4111
rect -6898 4011 -6864 4043
rect -6898 3941 -6864 3975
rect -6898 3873 -6864 3905
rect -6898 3805 -6864 3833
rect -6898 3737 -6864 3761
rect -6898 3669 -6864 3689
rect -6898 3601 -6864 3617
rect -6898 3533 -6864 3545
rect -6898 3454 -6864 3473
rect -6802 4443 -6768 4462
rect -6802 4371 -6768 4383
rect -6802 4299 -6768 4315
rect -6802 4227 -6768 4247
rect -6802 4155 -6768 4179
rect -6802 4083 -6768 4111
rect -6802 4011 -6768 4043
rect -6802 3941 -6768 3975
rect -6802 3873 -6768 3905
rect -6802 3805 -6768 3833
rect -6802 3737 -6768 3761
rect -6802 3669 -6768 3689
rect -6802 3601 -6768 3617
rect -6802 3533 -6768 3545
rect -6802 3396 -6768 3473
rect -6706 4443 -6672 4504
rect -6706 4371 -6672 4383
rect -6706 4299 -6672 4315
rect -6706 4227 -6672 4247
rect -6706 4155 -6672 4179
rect -6706 4083 -6672 4111
rect -6706 4011 -6672 4043
rect -6706 3941 -6672 3975
rect -6706 3873 -6672 3905
rect -6706 3805 -6672 3833
rect -6706 3737 -6672 3761
rect -6706 3669 -6672 3689
rect -6706 3601 -6672 3617
rect -6706 3533 -6672 3545
rect -6706 3454 -6672 3473
rect -6462 4508 -5468 4532
rect -6462 4449 -6428 4508
rect -6462 4377 -6428 4389
rect -6462 4305 -6428 4321
rect -6462 4233 -6428 4253
rect -6462 4161 -6428 4185
rect -6462 4089 -6428 4117
rect -6462 4017 -6428 4049
rect -6462 3947 -6428 3981
rect -6462 3879 -6428 3911
rect -6462 3811 -6428 3839
rect -6462 3743 -6428 3767
rect -6462 3675 -6428 3695
rect -6462 3607 -6428 3623
rect -6462 3539 -6428 3551
rect -6462 3460 -6428 3479
rect -6366 4449 -6332 4468
rect -6366 4377 -6332 4389
rect -6366 4305 -6332 4321
rect -6366 4233 -6332 4253
rect -6366 4161 -6332 4185
rect -6366 4089 -6332 4117
rect -6366 4017 -6332 4049
rect -6366 3947 -6332 3981
rect -6366 3879 -6332 3911
rect -6366 3811 -6332 3839
rect -6366 3743 -6332 3767
rect -6366 3675 -6332 3695
rect -6366 3607 -6332 3623
rect -6366 3539 -6332 3551
rect -11344 3247 -11328 3281
rect -11294 3247 -11278 3281
rect -12036 3040 -12020 3074
rect -11986 3040 -11970 3074
rect -20000 2759 -19966 2771
rect -20000 2687 -19966 2703
rect -20000 2615 -19966 2635
rect -20000 2543 -19966 2567
rect -20000 2471 -19966 2499
rect -20000 2399 -19966 2431
rect -20000 2329 -19966 2363
rect -20000 2261 -19966 2293
rect -20000 2193 -19966 2221
rect -20000 2125 -19966 2149
rect -20000 2057 -19966 2077
rect -20000 1989 -19966 2005
rect -20000 1921 -19966 1933
rect -20000 1842 -19966 1861
rect -19904 2831 -19870 2850
rect -19904 2759 -19870 2771
rect -19904 2687 -19870 2703
rect -19904 2615 -19870 2635
rect -19904 2543 -19870 2567
rect -19904 2471 -19870 2499
rect -19904 2399 -19870 2431
rect -19904 2329 -19870 2363
rect -19904 2261 -19870 2293
rect -19904 2193 -19870 2221
rect -19904 2125 -19870 2149
rect -19904 2057 -19870 2077
rect -19904 1989 -19870 2005
rect -19904 1921 -19870 1933
rect -19904 1800 -19870 1861
rect -21260 1790 -19870 1800
rect -19666 2835 -19632 2854
rect -19666 2763 -19632 2775
rect -19666 2691 -19632 2707
rect -19666 2619 -19632 2639
rect -19666 2547 -19632 2571
rect -19666 2475 -19632 2503
rect -19666 2403 -19632 2435
rect -19666 2333 -19632 2367
rect -19666 2265 -19632 2297
rect -19666 2197 -19632 2225
rect -19666 2129 -19632 2153
rect -19666 2061 -19632 2081
rect -19666 1993 -19632 2009
rect -19666 1925 -19632 1937
rect -19666 1812 -19632 1865
rect -19570 2835 -19536 2908
rect -19570 2763 -19536 2775
rect -19570 2691 -19536 2707
rect -19570 2619 -19536 2639
rect -19570 2547 -19536 2571
rect -19570 2475 -19536 2503
rect -19570 2403 -19536 2435
rect -19570 2333 -19536 2367
rect -19570 2265 -19536 2297
rect -19570 2197 -19536 2225
rect -19570 2129 -19536 2153
rect -19570 2061 -19536 2081
rect -19570 1993 -19536 2009
rect -19570 1925 -19536 1937
rect -19570 1846 -19536 1865
rect -19474 2835 -19440 2854
rect -19474 2763 -19440 2775
rect -19474 2691 -19440 2707
rect -19474 2619 -19440 2639
rect -19474 2547 -19440 2571
rect -19474 2475 -19440 2503
rect -19474 2403 -19440 2435
rect -19474 2333 -19440 2367
rect -19474 2265 -19440 2297
rect -19474 2197 -19440 2225
rect -19474 2129 -19440 2153
rect -19474 2061 -19440 2081
rect -19474 1993 -19440 2009
rect -19474 1925 -19440 1937
rect -19474 1812 -19440 1865
rect -19378 2835 -19344 2908
rect -19378 2763 -19344 2775
rect -19378 2691 -19344 2707
rect -19378 2619 -19344 2639
rect -19378 2547 -19344 2571
rect -19378 2475 -19344 2503
rect -19378 2403 -19344 2435
rect -19378 2333 -19344 2367
rect -19378 2265 -19344 2297
rect -19378 2197 -19344 2225
rect -19378 2129 -19344 2153
rect -19378 2061 -19344 2081
rect -19378 1993 -19344 2009
rect -19378 1925 -19344 1937
rect -19378 1846 -19344 1865
rect -19282 2835 -19248 2854
rect -19282 2763 -19248 2775
rect -19282 2691 -19248 2707
rect -19282 2619 -19248 2639
rect -19282 2547 -19248 2571
rect -19282 2475 -19248 2503
rect -19282 2403 -19248 2435
rect -19282 2333 -19248 2367
rect -19282 2265 -19248 2297
rect -19282 2197 -19248 2225
rect -19282 2129 -19248 2153
rect -19282 2061 -19248 2081
rect -19282 1993 -19248 2009
rect -19282 1925 -19248 1937
rect -19282 1812 -19248 1865
rect -19186 2835 -19152 2908
rect -19186 2763 -19152 2775
rect -19186 2691 -19152 2707
rect -19186 2619 -19152 2639
rect -19186 2547 -19152 2571
rect -19186 2475 -19152 2503
rect -19186 2403 -19152 2435
rect -19186 2333 -19152 2367
rect -19186 2265 -19152 2297
rect -19186 2197 -19152 2225
rect -19186 2129 -19152 2153
rect -19186 2061 -19152 2081
rect -19186 1993 -19152 2009
rect -19186 1925 -19152 1937
rect -19186 1846 -19152 1865
rect -19090 2835 -19056 2854
rect -19090 2763 -19056 2775
rect -19090 2691 -19056 2707
rect -19090 2619 -19056 2639
rect -19090 2547 -19056 2571
rect -19090 2475 -19056 2503
rect -19090 2403 -19056 2435
rect -19090 2333 -19056 2367
rect -19090 2265 -19056 2297
rect -19090 2197 -19056 2225
rect -19090 2129 -19056 2153
rect -19090 2061 -19056 2081
rect -19090 1993 -19056 2009
rect -19090 1925 -19056 1937
rect -19090 1812 -19056 1865
rect -18994 2835 -18960 2908
rect -18994 2763 -18960 2775
rect -18994 2691 -18960 2707
rect -18994 2619 -18960 2639
rect -18994 2547 -18960 2571
rect -18994 2475 -18960 2503
rect -18994 2403 -18960 2435
rect -18994 2333 -18960 2367
rect -18994 2265 -18960 2297
rect -18994 2197 -18960 2225
rect -18994 2129 -18960 2153
rect -18994 2061 -18960 2081
rect -18994 1993 -18960 2009
rect -18994 1925 -18960 1937
rect -18994 1846 -18960 1865
rect -18898 2835 -18864 2854
rect -18898 2763 -18864 2775
rect -18898 2691 -18864 2707
rect -18898 2619 -18864 2639
rect -18898 2547 -18864 2571
rect -18898 2475 -18864 2503
rect -18898 2403 -18864 2435
rect -18898 2333 -18864 2367
rect -18898 2265 -18864 2297
rect -18898 2197 -18864 2225
rect -18898 2129 -18864 2153
rect -18898 2061 -18864 2081
rect -18898 1993 -18864 2009
rect -18898 1925 -18864 1937
rect -18898 1812 -18864 1865
rect -18802 2835 -18768 2908
rect -18494 2898 -18076 2932
rect -16568 2908 -14804 2942
rect -18802 2763 -18768 2775
rect -18802 2691 -18768 2707
rect -18802 2619 -18768 2639
rect -18802 2547 -18768 2571
rect -18802 2475 -18768 2503
rect -18802 2403 -18768 2435
rect -18802 2333 -18768 2367
rect -18802 2265 -18768 2297
rect -18802 2197 -18768 2225
rect -18802 2129 -18768 2153
rect -18802 2061 -18768 2081
rect -18802 1993 -18768 2009
rect -18802 1925 -18768 1937
rect -18802 1846 -18768 1865
rect -18706 2835 -18672 2854
rect -18706 2763 -18672 2775
rect -18706 2691 -18672 2707
rect -18706 2619 -18672 2639
rect -18706 2547 -18672 2571
rect -18706 2475 -18672 2503
rect -18706 2403 -18672 2435
rect -18706 2333 -18672 2367
rect -18706 2265 -18672 2297
rect -18706 2197 -18672 2225
rect -18706 2129 -18672 2153
rect -18706 2061 -18672 2081
rect -18706 1993 -18672 2009
rect -18706 1925 -18672 1937
rect -18706 1812 -18672 1865
rect -18494 2845 -18460 2898
rect -18494 2773 -18460 2785
rect -18494 2701 -18460 2717
rect -18494 2629 -18460 2649
rect -18494 2557 -18460 2581
rect -18494 2485 -18460 2513
rect -18494 2413 -18460 2445
rect -18494 2343 -18460 2377
rect -18494 2275 -18460 2307
rect -18494 2207 -18460 2235
rect -18494 2139 -18460 2163
rect -18494 2071 -18460 2091
rect -18494 2003 -18460 2019
rect -18494 1935 -18460 1947
rect -18494 1856 -18460 1875
rect -18398 2845 -18364 2864
rect -18398 2773 -18364 2785
rect -18398 2701 -18364 2717
rect -18398 2629 -18364 2649
rect -18398 2557 -18364 2581
rect -18398 2485 -18364 2513
rect -18398 2413 -18364 2445
rect -18398 2343 -18364 2377
rect -18398 2275 -18364 2307
rect -18398 2207 -18364 2235
rect -18398 2139 -18364 2163
rect -18398 2071 -18364 2091
rect -18398 2003 -18364 2019
rect -18398 1935 -18364 1947
rect -19666 1790 -18672 1812
rect -18398 1808 -18364 1875
rect -18302 2845 -18268 2898
rect -18302 2773 -18268 2785
rect -18302 2701 -18268 2717
rect -18302 2629 -18268 2649
rect -18302 2557 -18268 2581
rect -18302 2485 -18268 2513
rect -18302 2413 -18268 2445
rect -18302 2343 -18268 2377
rect -18302 2275 -18268 2307
rect -18302 2207 -18268 2235
rect -18302 2139 -18268 2163
rect -18302 2071 -18268 2091
rect -18302 2003 -18268 2019
rect -18302 1935 -18268 1947
rect -18302 1856 -18268 1875
rect -18206 2845 -18172 2864
rect -18206 2773 -18172 2785
rect -18206 2701 -18172 2717
rect -18206 2629 -18172 2649
rect -18206 2557 -18172 2581
rect -18206 2485 -18172 2513
rect -18206 2413 -18172 2445
rect -18206 2343 -18172 2377
rect -18206 2275 -18172 2307
rect -18206 2207 -18172 2235
rect -18206 2139 -18172 2163
rect -18206 2071 -18172 2091
rect -18206 2003 -18172 2019
rect -18206 1935 -18172 1947
rect -18206 1808 -18172 1875
rect -18110 2845 -18076 2898
rect -18110 2773 -18076 2785
rect -18110 2701 -18076 2717
rect -18110 2629 -18076 2649
rect -18110 2557 -18076 2581
rect -18110 2485 -18076 2513
rect -18110 2413 -18076 2445
rect -18110 2343 -18076 2377
rect -18110 2275 -18076 2307
rect -18110 2207 -18076 2235
rect -18110 2139 -18076 2163
rect -18110 2071 -18076 2091
rect -18110 2003 -18076 2019
rect -18110 1935 -18076 1947
rect -18110 1856 -18076 1875
rect -18014 2845 -17980 2864
rect -18014 2773 -17980 2785
rect -18014 2701 -17980 2717
rect -18014 2629 -17980 2649
rect -18014 2557 -17980 2581
rect -18014 2485 -17980 2513
rect -18014 2413 -17980 2445
rect -18014 2343 -17980 2377
rect -18014 2275 -17980 2307
rect -18014 2207 -17980 2235
rect -18014 2139 -17980 2163
rect -18014 2071 -17980 2091
rect -18014 2003 -17980 2019
rect -18014 1935 -17980 1947
rect -18014 1808 -17980 1875
rect -18398 1790 -17980 1808
rect -23492 1774 -17980 1790
rect -16662 2851 -16628 2870
rect -16662 2779 -16628 2791
rect -16662 2707 -16628 2723
rect -16662 2635 -16628 2655
rect -16662 2563 -16628 2587
rect -16662 2491 -16628 2519
rect -16662 2419 -16628 2451
rect -16662 2349 -16628 2383
rect -16662 2281 -16628 2313
rect -16662 2213 -16628 2241
rect -16662 2145 -16628 2169
rect -16662 2077 -16628 2097
rect -16662 2009 -16628 2025
rect -16662 1941 -16628 1953
rect -16662 1820 -16628 1881
rect -16566 2851 -16532 2908
rect -16566 2779 -16532 2791
rect -16566 2707 -16532 2723
rect -16566 2635 -16532 2655
rect -16566 2563 -16532 2587
rect -16566 2491 -16532 2519
rect -16566 2419 -16532 2451
rect -16566 2349 -16532 2383
rect -16566 2281 -16532 2313
rect -16566 2213 -16532 2241
rect -16566 2145 -16532 2169
rect -16566 2077 -16532 2097
rect -16566 2009 -16532 2025
rect -16566 1941 -16532 1953
rect -16566 1862 -16532 1881
rect -16470 2851 -16436 2870
rect -16470 2779 -16436 2791
rect -16470 2707 -16436 2723
rect -16470 2635 -16436 2655
rect -16470 2563 -16436 2587
rect -16470 2491 -16436 2519
rect -16470 2419 -16436 2451
rect -16470 2349 -16436 2383
rect -16470 2281 -16436 2313
rect -16470 2213 -16436 2241
rect -16470 2145 -16436 2169
rect -16470 2077 -16436 2097
rect -16470 2009 -16436 2025
rect -16470 1941 -16436 1953
rect -16470 1820 -16436 1881
rect -16374 2851 -16340 2908
rect -16374 2779 -16340 2791
rect -16374 2707 -16340 2723
rect -16374 2635 -16340 2655
rect -16374 2563 -16340 2587
rect -16374 2491 -16340 2519
rect -16374 2419 -16340 2451
rect -16374 2349 -16340 2383
rect -16374 2281 -16340 2313
rect -16374 2213 -16340 2241
rect -16374 2145 -16340 2169
rect -16374 2077 -16340 2097
rect -16374 2009 -16340 2025
rect -16374 1941 -16340 1953
rect -16374 1862 -16340 1881
rect -16278 2851 -16244 2870
rect -16278 2779 -16244 2791
rect -16278 2707 -16244 2723
rect -16278 2635 -16244 2655
rect -16278 2563 -16244 2587
rect -16278 2491 -16244 2519
rect -16278 2419 -16244 2451
rect -16278 2349 -16244 2383
rect -16278 2281 -16244 2313
rect -16278 2213 -16244 2241
rect -16278 2145 -16244 2169
rect -16278 2077 -16244 2097
rect -16278 2009 -16244 2025
rect -16278 1941 -16244 1953
rect -16278 1820 -16244 1881
rect -16182 2851 -16148 2908
rect -16182 2779 -16148 2791
rect -16182 2707 -16148 2723
rect -16182 2635 -16148 2655
rect -16182 2563 -16148 2587
rect -16182 2491 -16148 2519
rect -16182 2419 -16148 2451
rect -16182 2349 -16148 2383
rect -16182 2281 -16148 2313
rect -16182 2213 -16148 2241
rect -16182 2145 -16148 2169
rect -16182 2077 -16148 2097
rect -16182 2009 -16148 2025
rect -16182 1941 -16148 1953
rect -16182 1862 -16148 1881
rect -16086 2851 -16052 2870
rect -16086 2779 -16052 2791
rect -16086 2707 -16052 2723
rect -16086 2635 -16052 2655
rect -16086 2563 -16052 2587
rect -16086 2491 -16052 2519
rect -16086 2419 -16052 2451
rect -16086 2349 -16052 2383
rect -16086 2281 -16052 2313
rect -16086 2213 -16052 2241
rect -16086 2145 -16052 2169
rect -16086 2077 -16052 2097
rect -16086 2009 -16052 2025
rect -16086 1941 -16052 1953
rect -16086 1820 -16052 1881
rect -15990 2851 -15956 2908
rect -15990 2779 -15956 2791
rect -15990 2707 -15956 2723
rect -15990 2635 -15956 2655
rect -15990 2563 -15956 2587
rect -15990 2491 -15956 2519
rect -15990 2419 -15956 2451
rect -15990 2349 -15956 2383
rect -15990 2281 -15956 2313
rect -15990 2213 -15956 2241
rect -15990 2145 -15956 2169
rect -15990 2077 -15956 2097
rect -15990 2009 -15956 2025
rect -15990 1941 -15956 1953
rect -15990 1862 -15956 1881
rect -15894 2851 -15860 2870
rect -15894 2779 -15860 2791
rect -15894 2707 -15860 2723
rect -15894 2635 -15860 2655
rect -15894 2563 -15860 2587
rect -15894 2491 -15860 2519
rect -15894 2419 -15860 2451
rect -15894 2349 -15860 2383
rect -15894 2281 -15860 2313
rect -15894 2213 -15860 2241
rect -15894 2145 -15860 2169
rect -15894 2077 -15860 2097
rect -15894 2009 -15860 2025
rect -15894 1941 -15860 1953
rect -15894 1820 -15860 1881
rect -15798 2851 -15764 2908
rect -15798 2779 -15764 2791
rect -15798 2707 -15764 2723
rect -15798 2635 -15764 2655
rect -15798 2563 -15764 2587
rect -15798 2491 -15764 2519
rect -15798 2419 -15764 2451
rect -15798 2349 -15764 2383
rect -15798 2281 -15764 2313
rect -15798 2213 -15764 2241
rect -15798 2145 -15764 2169
rect -15798 2077 -15764 2097
rect -15798 2009 -15764 2025
rect -15798 1941 -15764 1953
rect -15798 1862 -15764 1881
rect -15702 2851 -15668 2870
rect -15702 2779 -15668 2791
rect -15702 2707 -15668 2723
rect -15702 2635 -15668 2655
rect -15702 2563 -15668 2587
rect -15702 2491 -15668 2519
rect -15702 2419 -15668 2451
rect -15702 2349 -15668 2383
rect -15702 2281 -15668 2313
rect -15702 2213 -15668 2241
rect -15702 2145 -15668 2169
rect -15702 2077 -15668 2097
rect -15702 2009 -15668 2025
rect -15702 1941 -15668 1953
rect -15702 1820 -15668 1881
rect -15606 2851 -15572 2908
rect -15606 2779 -15572 2791
rect -15606 2707 -15572 2723
rect -15606 2635 -15572 2655
rect -15606 2563 -15572 2587
rect -15606 2491 -15572 2519
rect -15606 2419 -15572 2451
rect -15606 2349 -15572 2383
rect -15606 2281 -15572 2313
rect -15606 2213 -15572 2241
rect -15606 2145 -15572 2169
rect -15606 2077 -15572 2097
rect -15606 2009 -15572 2025
rect -15606 1941 -15572 1953
rect -15606 1862 -15572 1881
rect -15510 2851 -15476 2870
rect -15510 2779 -15476 2791
rect -15510 2707 -15476 2723
rect -15510 2635 -15476 2655
rect -15510 2563 -15476 2587
rect -15510 2491 -15476 2519
rect -15510 2419 -15476 2451
rect -15510 2349 -15476 2383
rect -15510 2281 -15476 2313
rect -15510 2213 -15476 2241
rect -15510 2145 -15476 2169
rect -15510 2077 -15476 2097
rect -15510 2009 -15476 2025
rect -15510 1941 -15476 1953
rect -15510 1820 -15476 1881
rect -15414 2851 -15380 2908
rect -15414 2779 -15380 2791
rect -15414 2707 -15380 2723
rect -15414 2635 -15380 2655
rect -15414 2563 -15380 2587
rect -15414 2491 -15380 2519
rect -15414 2419 -15380 2451
rect -15414 2349 -15380 2383
rect -15414 2281 -15380 2313
rect -15414 2213 -15380 2241
rect -15414 2145 -15380 2169
rect -15414 2077 -15380 2097
rect -15414 2009 -15380 2025
rect -15414 1941 -15380 1953
rect -15414 1862 -15380 1881
rect -15318 2851 -15284 2870
rect -15318 2779 -15284 2791
rect -15318 2707 -15284 2723
rect -15318 2635 -15284 2655
rect -15318 2563 -15284 2587
rect -15318 2491 -15284 2519
rect -15318 2419 -15284 2451
rect -15318 2349 -15284 2383
rect -15318 2281 -15284 2313
rect -15318 2213 -15284 2241
rect -15318 2145 -15284 2169
rect -15318 2077 -15284 2097
rect -15318 2009 -15284 2025
rect -15318 1941 -15284 1953
rect -15318 1820 -15284 1881
rect -15222 2851 -15188 2908
rect -15222 2779 -15188 2791
rect -15222 2707 -15188 2723
rect -15222 2635 -15188 2655
rect -15222 2563 -15188 2587
rect -15222 2491 -15188 2519
rect -15222 2419 -15188 2451
rect -15222 2349 -15188 2383
rect -15222 2281 -15188 2313
rect -15222 2213 -15188 2241
rect -15222 2145 -15188 2169
rect -15222 2077 -15188 2097
rect -15222 2009 -15188 2025
rect -15222 1941 -15188 1953
rect -15222 1862 -15188 1881
rect -15126 2851 -15092 2870
rect -15126 2779 -15092 2791
rect -15126 2707 -15092 2723
rect -15126 2635 -15092 2655
rect -15126 2563 -15092 2587
rect -15126 2491 -15092 2519
rect -15126 2419 -15092 2451
rect -15126 2349 -15092 2383
rect -15126 2281 -15092 2313
rect -15126 2213 -15092 2241
rect -15126 2145 -15092 2169
rect -15126 2077 -15092 2097
rect -15126 2009 -15092 2025
rect -15126 1941 -15092 1953
rect -15126 1820 -15092 1881
rect -15030 2851 -14996 2908
rect -15030 2779 -14996 2791
rect -15030 2707 -14996 2723
rect -15030 2635 -14996 2655
rect -15030 2563 -14996 2587
rect -15030 2491 -14996 2519
rect -15030 2419 -14996 2451
rect -15030 2349 -14996 2383
rect -15030 2281 -14996 2313
rect -15030 2213 -14996 2241
rect -15030 2145 -14996 2169
rect -15030 2077 -14996 2097
rect -15030 2009 -14996 2025
rect -15030 1941 -14996 1953
rect -15030 1862 -14996 1881
rect -14934 2851 -14900 2870
rect -14934 2779 -14900 2791
rect -14934 2707 -14900 2723
rect -14934 2635 -14900 2655
rect -14934 2563 -14900 2587
rect -14934 2491 -14900 2519
rect -14934 2419 -14900 2451
rect -14934 2349 -14900 2383
rect -14934 2281 -14900 2313
rect -14934 2213 -14900 2241
rect -14934 2145 -14900 2169
rect -14934 2077 -14900 2097
rect -14934 2009 -14900 2025
rect -14934 1941 -14900 1953
rect -14934 1820 -14900 1881
rect -14838 2851 -14804 2908
rect -14514 2912 -13136 2946
rect -14838 2779 -14804 2791
rect -14838 2707 -14804 2723
rect -14838 2635 -14804 2655
rect -14838 2563 -14804 2587
rect -14838 2491 -14804 2519
rect -14838 2419 -14804 2451
rect -14838 2349 -14804 2383
rect -14838 2281 -14804 2313
rect -14838 2213 -14804 2241
rect -14838 2145 -14804 2169
rect -14838 2077 -14804 2097
rect -14838 2009 -14804 2025
rect -14838 1941 -14804 1953
rect -14838 1862 -14804 1881
rect -14742 2851 -14708 2870
rect -14742 2779 -14708 2791
rect -14742 2707 -14708 2723
rect -14742 2635 -14708 2655
rect -14742 2563 -14708 2587
rect -14742 2491 -14708 2519
rect -14742 2419 -14708 2451
rect -14742 2349 -14708 2383
rect -14742 2281 -14708 2313
rect -14742 2213 -14708 2241
rect -14742 2145 -14708 2169
rect -14742 2077 -14708 2097
rect -14742 2009 -14708 2025
rect -14742 1941 -14708 1953
rect -14742 1820 -14708 1881
rect -14514 2843 -14480 2912
rect -14514 2771 -14480 2783
rect -14514 2699 -14480 2715
rect -14514 2627 -14480 2647
rect -14514 2555 -14480 2579
rect -14514 2483 -14480 2511
rect -14514 2411 -14480 2443
rect -14514 2341 -14480 2375
rect -14514 2273 -14480 2305
rect -14514 2205 -14480 2233
rect -14514 2137 -14480 2161
rect -14514 2069 -14480 2089
rect -14514 2001 -14480 2017
rect -14514 1933 -14480 1945
rect -14514 1854 -14480 1873
rect -14418 2843 -14384 2862
rect -14418 2771 -14384 2783
rect -14418 2699 -14384 2715
rect -14418 2627 -14384 2647
rect -14418 2555 -14384 2579
rect -14418 2483 -14384 2511
rect -14418 2411 -14384 2443
rect -14418 2341 -14384 2375
rect -14418 2273 -14384 2305
rect -14418 2205 -14384 2233
rect -14418 2137 -14384 2161
rect -14418 2069 -14384 2089
rect -14418 2001 -14384 2017
rect -14418 1933 -14384 1945
rect -16662 1798 -14708 1820
rect -14418 1812 -14384 1873
rect -14322 2843 -14288 2912
rect -14322 2771 -14288 2783
rect -14322 2699 -14288 2715
rect -14322 2627 -14288 2647
rect -14322 2555 -14288 2579
rect -14322 2483 -14288 2511
rect -14322 2411 -14288 2443
rect -14322 2341 -14288 2375
rect -14322 2273 -14288 2305
rect -14322 2205 -14288 2233
rect -14322 2137 -14288 2161
rect -14322 2069 -14288 2089
rect -14322 2001 -14288 2017
rect -14322 1933 -14288 1945
rect -14322 1854 -14288 1873
rect -14226 2843 -14192 2862
rect -14226 2771 -14192 2783
rect -14226 2699 -14192 2715
rect -14226 2627 -14192 2647
rect -14226 2555 -14192 2579
rect -14226 2483 -14192 2511
rect -14226 2411 -14192 2443
rect -14226 2341 -14192 2375
rect -14226 2273 -14192 2305
rect -14226 2205 -14192 2233
rect -14226 2137 -14192 2161
rect -14226 2069 -14192 2089
rect -14226 2001 -14192 2017
rect -14226 1933 -14192 1945
rect -14226 1812 -14192 1873
rect -14130 2843 -14096 2912
rect -14130 2771 -14096 2783
rect -14130 2699 -14096 2715
rect -14130 2627 -14096 2647
rect -14130 2555 -14096 2579
rect -14130 2483 -14096 2511
rect -14130 2411 -14096 2443
rect -14130 2341 -14096 2375
rect -14130 2273 -14096 2305
rect -14130 2205 -14096 2233
rect -14130 2137 -14096 2161
rect -14130 2069 -14096 2089
rect -14130 2001 -14096 2017
rect -14130 1933 -14096 1945
rect -14130 1854 -14096 1873
rect -14034 2843 -14000 2862
rect -14034 2771 -14000 2783
rect -14034 2699 -14000 2715
rect -14034 2627 -14000 2647
rect -14034 2555 -14000 2579
rect -14034 2483 -14000 2511
rect -14034 2411 -14000 2443
rect -14034 2341 -14000 2375
rect -14034 2273 -14000 2305
rect -14034 2205 -14000 2233
rect -14034 2137 -14000 2161
rect -14034 2069 -14000 2089
rect -14034 2001 -14000 2017
rect -14034 1933 -14000 1945
rect -14034 1812 -14000 1873
rect -13938 2843 -13904 2912
rect -13938 2771 -13904 2783
rect -13938 2699 -13904 2715
rect -13938 2627 -13904 2647
rect -13938 2555 -13904 2579
rect -13938 2483 -13904 2511
rect -13938 2411 -13904 2443
rect -13938 2341 -13904 2375
rect -13938 2273 -13904 2305
rect -13938 2205 -13904 2233
rect -13938 2137 -13904 2161
rect -13938 2069 -13904 2089
rect -13938 2001 -13904 2017
rect -13938 1933 -13904 1945
rect -13938 1854 -13904 1873
rect -13842 2843 -13808 2862
rect -13842 2771 -13808 2783
rect -13842 2699 -13808 2715
rect -13842 2627 -13808 2647
rect -13842 2555 -13808 2579
rect -13842 2483 -13808 2511
rect -13842 2411 -13808 2443
rect -13842 2341 -13808 2375
rect -13842 2273 -13808 2305
rect -13842 2205 -13808 2233
rect -13842 2137 -13808 2161
rect -13842 2069 -13808 2089
rect -13842 2001 -13808 2017
rect -13842 1933 -13808 1945
rect -13842 1812 -13808 1873
rect -13746 2843 -13712 2912
rect -13746 2771 -13712 2783
rect -13746 2699 -13712 2715
rect -13746 2627 -13712 2647
rect -13746 2555 -13712 2579
rect -13746 2483 -13712 2511
rect -13746 2411 -13712 2443
rect -13746 2341 -13712 2375
rect -13746 2273 -13712 2305
rect -13746 2205 -13712 2233
rect -13746 2137 -13712 2161
rect -13746 2069 -13712 2089
rect -13746 2001 -13712 2017
rect -13746 1933 -13712 1945
rect -13746 1854 -13712 1873
rect -13650 2843 -13616 2862
rect -13650 2771 -13616 2783
rect -13650 2699 -13616 2715
rect -13650 2627 -13616 2647
rect -13650 2555 -13616 2579
rect -13650 2483 -13616 2511
rect -13650 2411 -13616 2443
rect -13650 2341 -13616 2375
rect -13650 2273 -13616 2305
rect -13650 2205 -13616 2233
rect -13650 2137 -13616 2161
rect -13650 2069 -13616 2089
rect -13650 2001 -13616 2017
rect -13650 1933 -13616 1945
rect -13650 1812 -13616 1873
rect -13554 2843 -13520 2912
rect -13554 2771 -13520 2783
rect -13554 2699 -13520 2715
rect -13554 2627 -13520 2647
rect -13554 2555 -13520 2579
rect -13554 2483 -13520 2511
rect -13554 2411 -13520 2443
rect -13554 2341 -13520 2375
rect -13554 2273 -13520 2305
rect -13554 2205 -13520 2233
rect -13554 2137 -13520 2161
rect -13554 2069 -13520 2089
rect -13554 2001 -13520 2017
rect -13554 1933 -13520 1945
rect -13554 1854 -13520 1873
rect -13458 2843 -13424 2862
rect -13458 2771 -13424 2783
rect -13458 2699 -13424 2715
rect -13458 2627 -13424 2647
rect -13458 2555 -13424 2579
rect -13458 2483 -13424 2511
rect -13458 2411 -13424 2443
rect -13458 2341 -13424 2375
rect -13458 2273 -13424 2305
rect -13458 2205 -13424 2233
rect -13458 2137 -13424 2161
rect -13458 2069 -13424 2089
rect -13458 2001 -13424 2017
rect -13458 1933 -13424 1945
rect -13458 1812 -13424 1873
rect -13362 2843 -13328 2912
rect -13362 2771 -13328 2783
rect -13362 2699 -13328 2715
rect -13362 2627 -13328 2647
rect -13362 2555 -13328 2579
rect -13362 2483 -13328 2511
rect -13362 2411 -13328 2443
rect -13362 2341 -13328 2375
rect -13362 2273 -13328 2305
rect -13362 2205 -13328 2233
rect -13362 2137 -13328 2161
rect -13362 2069 -13328 2089
rect -13362 2001 -13328 2017
rect -13362 1933 -13328 1945
rect -13362 1854 -13328 1873
rect -13266 2843 -13232 2862
rect -13266 2771 -13232 2783
rect -13266 2699 -13232 2715
rect -13266 2627 -13232 2647
rect -13266 2555 -13232 2579
rect -13266 2483 -13232 2511
rect -13266 2411 -13232 2443
rect -13266 2341 -13232 2375
rect -13266 2273 -13232 2305
rect -13266 2205 -13232 2233
rect -13266 2137 -13232 2161
rect -13266 2069 -13232 2089
rect -13266 2001 -13232 2017
rect -13266 1933 -13232 1945
rect -13266 1812 -13232 1873
rect -13170 2843 -13136 2912
rect -12740 2920 -11938 2954
rect -11472 2944 -11438 3125
rect -9684 3140 -9638 3368
rect -8146 3362 -6768 3396
rect -6366 3402 -6332 3479
rect -6270 4449 -6236 4508
rect -6270 4377 -6236 4389
rect -6270 4305 -6236 4321
rect -6270 4233 -6236 4253
rect -6270 4161 -6236 4185
rect -6270 4089 -6236 4117
rect -6270 4017 -6236 4049
rect -6270 3947 -6236 3981
rect -6270 3879 -6236 3911
rect -6270 3811 -6236 3839
rect -6270 3743 -6236 3767
rect -6270 3675 -6236 3695
rect -6270 3607 -6236 3623
rect -6270 3539 -6236 3551
rect -6270 3460 -6236 3479
rect -6174 4449 -6140 4468
rect -6174 4377 -6140 4389
rect -6174 4305 -6140 4321
rect -6174 4233 -6140 4253
rect -6174 4161 -6140 4185
rect -6174 4089 -6140 4117
rect -6174 4017 -6140 4049
rect -6174 3947 -6140 3981
rect -6174 3879 -6140 3911
rect -6174 3811 -6140 3839
rect -6174 3743 -6140 3767
rect -6174 3675 -6140 3695
rect -6174 3607 -6140 3623
rect -6174 3539 -6140 3551
rect -6174 3402 -6140 3479
rect -6078 4449 -6044 4508
rect -6078 4377 -6044 4389
rect -6078 4305 -6044 4321
rect -6078 4233 -6044 4253
rect -6078 4161 -6044 4185
rect -6078 4089 -6044 4117
rect -6078 4017 -6044 4049
rect -6078 3947 -6044 3981
rect -6078 3879 -6044 3911
rect -6078 3811 -6044 3839
rect -6078 3743 -6044 3767
rect -6078 3675 -6044 3695
rect -6078 3607 -6044 3623
rect -6078 3539 -6044 3551
rect -6078 3460 -6044 3479
rect -5982 4449 -5948 4468
rect -5982 4377 -5948 4389
rect -5982 4305 -5948 4321
rect -5982 4233 -5948 4253
rect -5982 4161 -5948 4185
rect -5982 4089 -5948 4117
rect -5982 4017 -5948 4049
rect -5982 3947 -5948 3981
rect -5982 3879 -5948 3911
rect -5982 3811 -5948 3839
rect -5982 3743 -5948 3767
rect -5982 3675 -5948 3695
rect -5982 3607 -5948 3623
rect -5982 3539 -5948 3551
rect -5982 3402 -5948 3479
rect -5886 4449 -5852 4508
rect -5886 4377 -5852 4389
rect -5886 4305 -5852 4321
rect -5886 4233 -5852 4253
rect -5886 4161 -5852 4185
rect -5886 4089 -5852 4117
rect -5886 4017 -5852 4049
rect -5886 3947 -5852 3981
rect -5886 3879 -5852 3911
rect -5886 3811 -5852 3839
rect -5886 3743 -5852 3767
rect -5886 3675 -5852 3695
rect -5886 3607 -5852 3623
rect -5886 3539 -5852 3551
rect -5886 3460 -5852 3479
rect -5790 4449 -5756 4468
rect -5790 4377 -5756 4389
rect -5790 4305 -5756 4321
rect -5790 4233 -5756 4253
rect -5790 4161 -5756 4185
rect -5790 4089 -5756 4117
rect -5790 4017 -5756 4049
rect -5790 3947 -5756 3981
rect -5790 3879 -5756 3911
rect -5790 3811 -5756 3839
rect -5790 3743 -5756 3767
rect -5790 3675 -5756 3695
rect -5790 3607 -5756 3623
rect -5790 3539 -5756 3551
rect -5790 3402 -5756 3479
rect -5694 4449 -5660 4508
rect -5694 4377 -5660 4389
rect -5694 4305 -5660 4321
rect -5694 4233 -5660 4253
rect -5694 4161 -5660 4185
rect -5694 4089 -5660 4117
rect -5694 4017 -5660 4049
rect -5694 3947 -5660 3981
rect -5694 3879 -5660 3911
rect -5694 3811 -5660 3839
rect -5694 3743 -5660 3767
rect -5694 3675 -5660 3695
rect -5694 3607 -5660 3623
rect -5694 3539 -5660 3551
rect -5694 3460 -5660 3479
rect -5598 4449 -5564 4468
rect -5598 4377 -5564 4389
rect -5598 4305 -5564 4321
rect -5598 4233 -5564 4253
rect -5598 4161 -5564 4185
rect -5598 4089 -5564 4117
rect -5598 4017 -5564 4049
rect -5598 3947 -5564 3981
rect -5598 3879 -5564 3911
rect -5598 3811 -5564 3839
rect -5598 3743 -5564 3767
rect -5598 3675 -5564 3695
rect -5598 3607 -5564 3623
rect -5598 3539 -5564 3551
rect -5598 3402 -5564 3479
rect -5502 4449 -5468 4508
rect -5198 4510 -4780 4532
rect -5502 4377 -5468 4389
rect -5502 4305 -5468 4321
rect -5502 4233 -5468 4253
rect -5502 4161 -5468 4185
rect -5502 4089 -5468 4117
rect -5502 4017 -5468 4049
rect -5502 3947 -5468 3981
rect -5502 3879 -5468 3911
rect -5502 3811 -5468 3839
rect -5502 3743 -5468 3767
rect -5502 3675 -5468 3695
rect -5502 3607 -5468 3623
rect -5502 3539 -5468 3551
rect -5502 3460 -5468 3479
rect -5294 4451 -5260 4470
rect -5294 4379 -5260 4391
rect -5294 4307 -5260 4323
rect -5294 4235 -5260 4255
rect -5294 4163 -5260 4187
rect -5294 4091 -5260 4119
rect -5294 4019 -5260 4051
rect -5294 3949 -5260 3983
rect -5294 3881 -5260 3913
rect -5294 3813 -5260 3841
rect -5294 3745 -5260 3769
rect -5294 3677 -5260 3697
rect -5294 3609 -5260 3625
rect -5294 3541 -5260 3553
rect -6366 3368 -5564 3402
rect -5294 3410 -5260 3481
rect -5198 4451 -5164 4510
rect -5198 4379 -5164 4391
rect -5198 4307 -5164 4323
rect -5198 4235 -5164 4255
rect -5198 4163 -5164 4187
rect -5198 4091 -5164 4119
rect -5198 4019 -5164 4051
rect -5198 3949 -5164 3983
rect -5198 3881 -5164 3913
rect -5198 3813 -5164 3841
rect -5198 3745 -5164 3769
rect -5198 3677 -5164 3697
rect -5198 3609 -5164 3625
rect -5198 3541 -5164 3553
rect -5198 3462 -5164 3481
rect -5102 4451 -5068 4470
rect -5102 4379 -5068 4391
rect -5102 4307 -5068 4323
rect -5102 4235 -5068 4255
rect -5102 4163 -5068 4187
rect -5102 4091 -5068 4119
rect -5102 4019 -5068 4051
rect -5102 3949 -5068 3983
rect -5102 3881 -5068 3913
rect -5102 3813 -5068 3841
rect -5102 3745 -5068 3769
rect -5102 3677 -5068 3697
rect -5102 3609 -5068 3625
rect -5102 3541 -5068 3553
rect -5102 3410 -5068 3481
rect -5006 4451 -4972 4510
rect -5006 4379 -4972 4391
rect -5006 4307 -4972 4323
rect -5006 4235 -4972 4255
rect -5006 4163 -4972 4187
rect -5006 4091 -4972 4119
rect -5006 4019 -4972 4051
rect -5006 3949 -4972 3983
rect -5006 3881 -4972 3913
rect -5006 3813 -4972 3841
rect -5006 3745 -4972 3769
rect -5006 3677 -4972 3697
rect -5006 3609 -4972 3625
rect -5006 3541 -4972 3553
rect -5006 3462 -4972 3481
rect -4910 4451 -4876 4470
rect -4910 4379 -4876 4391
rect -4910 4307 -4876 4323
rect -4910 4235 -4876 4255
rect -4910 4163 -4876 4187
rect -4910 4091 -4876 4119
rect -4910 4019 -4876 4051
rect -4910 3949 -4876 3983
rect -4910 3881 -4876 3913
rect -4910 3813 -4876 3841
rect -4910 3745 -4876 3769
rect -4910 3677 -4876 3697
rect -4910 3609 -4876 3625
rect -4910 3541 -4876 3553
rect -4910 3410 -4876 3481
rect -4814 4451 -4780 4510
rect -4814 4379 -4780 4391
rect -4814 4307 -4780 4323
rect -4814 4235 -4780 4255
rect -4814 4163 -4780 4187
rect -4814 4091 -4780 4119
rect -4814 4019 -4780 4051
rect -4814 3949 -4780 3983
rect 1484 4497 1518 4529
rect 1484 4427 1518 4461
rect 1484 4359 1518 4391
rect 1484 4291 1518 4319
rect 1484 4223 1518 4247
rect 1484 4155 1518 4175
rect 1484 4087 1518 4103
rect 1484 4019 1518 4031
rect 1484 3940 1518 3959
rect 1580 4929 1614 4946
rect 1580 4857 1614 4869
rect 1580 4785 1614 4801
rect 1580 4713 1614 4733
rect 1580 4641 1614 4665
rect 1580 4569 1614 4597
rect 1580 4497 1614 4529
rect 1580 4427 1614 4461
rect 1580 4359 1614 4391
rect 1580 4291 1614 4319
rect 1580 4223 1614 4247
rect 1580 4155 1614 4175
rect 1580 4087 1614 4103
rect 1580 4019 1614 4031
rect -4814 3881 -4780 3913
rect 1580 3884 1614 3959
rect 1676 4929 1710 4994
rect 1676 4857 1710 4869
rect 1676 4785 1710 4801
rect 1676 4713 1710 4733
rect 1676 4641 1710 4665
rect 1676 4569 1710 4597
rect 1676 4497 1710 4529
rect 1676 4427 1710 4461
rect 1676 4359 1710 4391
rect 1676 4291 1710 4319
rect 1676 4223 1710 4247
rect 1676 4155 1710 4175
rect 1676 4087 1710 4103
rect 1676 4019 1710 4031
rect 1676 3940 1710 3959
rect 1772 4929 1806 4946
rect 1772 4857 1806 4869
rect 1772 4785 1806 4801
rect 1772 4713 1806 4733
rect 1772 4641 1806 4665
rect 1772 4569 1806 4597
rect 1772 4497 1806 4529
rect 1772 4427 1806 4461
rect 1772 4359 1806 4391
rect 1772 4291 1806 4319
rect 1772 4223 1806 4247
rect 1772 4155 1806 4175
rect 1772 4087 1806 4103
rect 1772 4019 1806 4031
rect 1676 3884 1710 3886
rect 1772 3884 1806 3959
rect 1868 4929 1902 4994
rect 4438 4978 4864 5012
rect 7468 4978 7894 5012
rect 10654 5010 10688 5072
rect 1868 4857 1902 4869
rect 1868 4785 1902 4801
rect 1868 4713 1902 4733
rect 1868 4641 1902 4665
rect 1868 4569 1902 4597
rect 1868 4497 1902 4529
rect 1868 4427 1902 4461
rect 1868 4359 1902 4391
rect 1868 4291 1902 4319
rect 1868 4223 1902 4247
rect 1868 4155 1902 4175
rect 1868 4087 1902 4103
rect 1868 4019 1902 4031
rect 1868 3940 1902 3959
rect 4440 4913 4474 4978
rect 4440 4841 4474 4853
rect 4440 4769 4474 4785
rect 4440 4697 4474 4717
rect 4440 4625 4474 4649
rect 4440 4553 4474 4581
rect 4440 4481 4474 4513
rect 4440 4411 4474 4445
rect 4440 4343 4474 4375
rect 4440 4275 4474 4303
rect 4440 4207 4474 4231
rect 4440 4139 4474 4159
rect 4440 4071 4474 4087
rect 4440 4003 4474 4015
rect 4440 3924 4474 3943
rect 4536 4913 4570 4930
rect 4536 4841 4570 4853
rect 4536 4769 4570 4785
rect 4536 4697 4570 4717
rect 4536 4625 4570 4649
rect 4536 4553 4570 4581
rect 4536 4481 4570 4513
rect 4536 4411 4570 4445
rect 4536 4343 4570 4375
rect 4536 4275 4570 4303
rect 4536 4207 4570 4231
rect 4536 4139 4570 4159
rect 4536 4071 4570 4087
rect 4536 4003 4570 4015
rect 1580 3850 1806 3884
rect 4536 3868 4570 3943
rect 4632 4913 4666 4978
rect 4632 4841 4666 4853
rect 4632 4769 4666 4785
rect 4632 4697 4666 4717
rect 4632 4625 4666 4649
rect 4632 4553 4666 4581
rect 4632 4481 4666 4513
rect 4632 4411 4666 4445
rect 4632 4343 4666 4375
rect 4632 4275 4666 4303
rect 4632 4207 4666 4231
rect 4632 4139 4666 4159
rect 4632 4071 4666 4087
rect 4632 4003 4666 4015
rect 4632 3924 4666 3943
rect 4728 4913 4762 4930
rect 4728 4841 4762 4853
rect 4728 4769 4762 4785
rect 4728 4697 4762 4717
rect 4728 4625 4762 4649
rect 4728 4553 4762 4581
rect 4728 4481 4762 4513
rect 4728 4411 4762 4445
rect 4728 4343 4762 4375
rect 4728 4275 4762 4303
rect 4728 4207 4762 4231
rect 4728 4139 4762 4159
rect 4728 4071 4762 4087
rect 4728 4003 4762 4015
rect 4632 3868 4666 3870
rect 4728 3868 4762 3943
rect 4824 4913 4858 4978
rect 4824 4841 4858 4853
rect 4824 4769 4858 4785
rect 4824 4697 4858 4717
rect 4824 4625 4858 4649
rect 4824 4553 4858 4581
rect 4824 4481 4858 4513
rect 4824 4411 4858 4445
rect 4824 4343 4858 4375
rect 4824 4275 4858 4303
rect 4824 4207 4858 4231
rect 4824 4139 4858 4159
rect 4824 4071 4858 4087
rect 4824 4003 4858 4015
rect 4824 3924 4858 3943
rect 7470 4913 7504 4978
rect 7470 4841 7504 4853
rect 7470 4769 7504 4785
rect 7470 4697 7504 4717
rect 7470 4625 7504 4649
rect 7470 4553 7504 4581
rect 7470 4481 7504 4513
rect 7470 4411 7504 4445
rect 7470 4343 7504 4375
rect 7470 4275 7504 4303
rect 7470 4207 7504 4231
rect 7470 4139 7504 4159
rect 7470 4071 7504 4087
rect 7470 4003 7504 4015
rect 7470 3924 7504 3943
rect 7566 4913 7600 4930
rect 7566 4841 7600 4853
rect 7566 4769 7600 4785
rect 7566 4697 7600 4717
rect 7566 4625 7600 4649
rect 7566 4553 7600 4581
rect 7566 4481 7600 4513
rect 7566 4411 7600 4445
rect 7566 4343 7600 4375
rect 7566 4275 7600 4303
rect 7566 4207 7600 4231
rect 7566 4139 7600 4159
rect 7566 4071 7600 4087
rect 7566 4003 7600 4015
rect -4814 3813 -4780 3841
rect -4814 3745 -4780 3769
rect 1564 3743 1580 3777
rect 1614 3743 1630 3777
rect 1676 3754 1710 3850
rect 4536 3834 4762 3868
rect 7566 3868 7600 3943
rect 7662 4913 7696 4978
rect 7662 4841 7696 4853
rect 7662 4769 7696 4785
rect 7662 4697 7696 4717
rect 7662 4625 7696 4649
rect 7662 4553 7696 4581
rect 7662 4481 7696 4513
rect 7662 4411 7696 4445
rect 7662 4343 7696 4375
rect 7662 4275 7696 4303
rect 7662 4207 7696 4231
rect 7662 4139 7696 4159
rect 7662 4071 7696 4087
rect 7662 4003 7696 4015
rect 7662 3924 7696 3943
rect 7758 4913 7792 4930
rect 7758 4841 7792 4853
rect 7758 4769 7792 4785
rect 7758 4697 7792 4717
rect 7758 4625 7792 4649
rect 7758 4553 7792 4581
rect 7758 4481 7792 4513
rect 7758 4411 7792 4445
rect 7758 4343 7792 4375
rect 7758 4275 7792 4303
rect 7758 4207 7792 4231
rect 7758 4139 7792 4159
rect 7758 4071 7792 4087
rect 7758 4003 7792 4015
rect 7662 3868 7696 3870
rect 7758 3868 7792 3943
rect 7854 4913 7888 4978
rect 10556 4976 10982 5010
rect 13810 4984 13844 5046
rect 15518 5015 15552 5045
rect 7854 4841 7888 4853
rect 7854 4769 7888 4785
rect 7854 4697 7888 4717
rect 7854 4625 7888 4649
rect 7854 4553 7888 4581
rect 7854 4481 7888 4513
rect 7854 4411 7888 4445
rect 7854 4343 7888 4375
rect 7854 4275 7888 4303
rect 7854 4207 7888 4231
rect 7854 4139 7888 4159
rect 7854 4071 7888 4087
rect 7854 4003 7888 4015
rect 7854 3924 7888 3943
rect 10558 4911 10592 4976
rect 10558 4839 10592 4851
rect 10558 4767 10592 4783
rect 10558 4695 10592 4715
rect 10558 4623 10592 4647
rect 10558 4551 10592 4579
rect 10558 4479 10592 4511
rect 10558 4409 10592 4443
rect 10558 4341 10592 4373
rect 10558 4273 10592 4301
rect 10558 4205 10592 4229
rect 10558 4137 10592 4157
rect 10558 4069 10592 4085
rect 10558 4001 10592 4013
rect 10558 3922 10592 3941
rect 10654 4911 10688 4928
rect 10654 4839 10688 4851
rect 10654 4767 10688 4783
rect 10654 4695 10688 4715
rect 10654 4623 10688 4647
rect 10654 4551 10688 4579
rect 10654 4479 10688 4511
rect 10654 4409 10688 4443
rect 10654 4341 10688 4373
rect 10654 4273 10688 4301
rect 10654 4205 10688 4229
rect 10654 4137 10688 4157
rect 10654 4069 10688 4085
rect 10654 4001 10688 4013
rect 7566 3834 7792 3868
rect 10654 3866 10688 3941
rect 10750 4911 10784 4976
rect 10750 4839 10784 4851
rect 10750 4767 10784 4783
rect 10750 4695 10784 4715
rect 10750 4623 10784 4647
rect 10750 4551 10784 4579
rect 10750 4479 10784 4511
rect 10750 4409 10784 4443
rect 10750 4341 10784 4373
rect 10750 4273 10784 4301
rect 10750 4205 10784 4229
rect 10750 4137 10784 4157
rect 10750 4069 10784 4085
rect 10750 4001 10784 4013
rect 10750 3922 10784 3941
rect 10846 4911 10880 4928
rect 10846 4839 10880 4851
rect 10846 4767 10880 4783
rect 10846 4695 10880 4715
rect 10846 4623 10880 4647
rect 10846 4551 10880 4579
rect 10846 4479 10880 4511
rect 10846 4409 10880 4443
rect 10846 4341 10880 4373
rect 10846 4273 10880 4301
rect 10846 4205 10880 4229
rect 10846 4137 10880 4157
rect 10846 4069 10880 4085
rect 10846 4001 10880 4013
rect 10750 3866 10784 3868
rect 10846 3866 10880 3941
rect 10942 4911 10976 4976
rect 13712 4950 14138 4984
rect 10942 4839 10976 4851
rect 10942 4767 10976 4783
rect 10942 4695 10976 4715
rect 10942 4623 10976 4647
rect 10942 4551 10976 4579
rect 10942 4479 10976 4511
rect 10942 4409 10976 4443
rect 10942 4341 10976 4373
rect 10942 4273 10976 4301
rect 10942 4205 10976 4229
rect 10942 4137 10976 4157
rect 10942 4069 10976 4085
rect 10942 4001 10976 4013
rect 10942 3922 10976 3941
rect 13714 4885 13748 4950
rect 13714 4813 13748 4825
rect 13714 4741 13748 4757
rect 13714 4669 13748 4689
rect 13714 4597 13748 4621
rect 13714 4525 13748 4553
rect 13714 4453 13748 4485
rect 13714 4383 13748 4417
rect 13714 4315 13748 4347
rect 13714 4247 13748 4275
rect 13714 4179 13748 4203
rect 13714 4111 13748 4131
rect 13714 4043 13748 4059
rect 13714 3975 13748 3987
rect 13714 3896 13748 3915
rect 13810 4885 13844 4902
rect 13810 4813 13844 4825
rect 13810 4741 13844 4757
rect 13810 4669 13844 4689
rect 13810 4597 13844 4621
rect 13810 4525 13844 4553
rect 13810 4453 13844 4485
rect 13810 4383 13844 4417
rect 13810 4315 13844 4347
rect 13810 4247 13844 4275
rect 13810 4179 13844 4203
rect 13810 4111 13844 4131
rect 13810 4043 13844 4059
rect 13810 3975 13844 3987
rect 1756 3743 1772 3777
rect 1806 3743 1822 3777
rect 4520 3727 4536 3761
rect 4570 3727 4586 3761
rect 4632 3738 4666 3834
rect 4712 3727 4728 3761
rect 4762 3727 4778 3761
rect 7550 3727 7566 3761
rect 7600 3727 7616 3761
rect 7662 3738 7696 3834
rect 10654 3832 10880 3866
rect 13810 3840 13844 3915
rect 13906 4885 13940 4950
rect 13906 4813 13940 4825
rect 13906 4741 13940 4757
rect 13906 4669 13940 4689
rect 13906 4597 13940 4621
rect 13906 4525 13940 4553
rect 13906 4453 13940 4485
rect 13906 4383 13940 4417
rect 13906 4315 13940 4347
rect 13906 4247 13940 4275
rect 13906 4179 13940 4203
rect 13906 4111 13940 4131
rect 13906 4043 13940 4059
rect 13906 3975 13940 3987
rect 13906 3896 13940 3915
rect 14002 4885 14036 4902
rect 14002 4813 14036 4825
rect 14002 4741 14036 4757
rect 14002 4669 14036 4689
rect 14002 4597 14036 4621
rect 14002 4525 14036 4553
rect 14002 4453 14036 4485
rect 14002 4383 14036 4417
rect 14002 4315 14036 4347
rect 14002 4247 14036 4275
rect 14002 4179 14036 4203
rect 14002 4111 14036 4131
rect 14002 4043 14036 4059
rect 14002 3975 14036 3987
rect 13906 3840 13940 3842
rect 14002 3840 14036 3915
rect 14098 4885 14132 4950
rect 14098 4813 14132 4825
rect 14098 4741 14132 4757
rect 14098 4669 14132 4689
rect 14098 4597 14132 4621
rect 14098 4525 14132 4553
rect 14098 4453 14132 4485
rect 14098 4383 14132 4417
rect 14098 4315 14132 4347
rect 14098 4247 14132 4275
rect 14098 4179 14132 4203
rect 14098 4111 14132 4131
rect 14098 4043 14132 4059
rect 14098 3975 14132 3987
rect 15518 4943 15552 4977
rect 15518 4875 15552 4909
rect 15518 4807 15552 4837
rect 15518 4739 15552 4765
rect 15518 4671 15552 4693
rect 15518 4603 15552 4621
rect 15518 4535 15552 4549
rect 15518 4467 15552 4477
rect 15518 4399 15552 4405
rect 15518 4331 15552 4333
rect 15518 4295 15552 4297
rect 15518 4223 15552 4229
rect 15518 4151 15552 4161
rect 15518 4079 15552 4093
rect 15518 4007 15552 4025
rect 15518 3918 15552 3957
rect 15614 5895 15648 5930
rect 15614 5827 15648 5845
rect 15614 5759 15648 5773
rect 15614 5691 15648 5701
rect 15614 5623 15648 5629
rect 15614 5555 15648 5557
rect 15614 5519 15648 5521
rect 15614 5447 15648 5453
rect 15614 5375 15648 5385
rect 15614 5303 15648 5317
rect 15614 5231 15648 5249
rect 15614 5159 15648 5181
rect 15614 5087 15648 5113
rect 15614 5015 15648 5045
rect 15614 4943 15648 4977
rect 15614 4875 15648 4909
rect 15614 4807 15648 4837
rect 15614 4739 15648 4765
rect 15614 4671 15648 4693
rect 15614 4603 15648 4621
rect 15614 4535 15648 4549
rect 15614 4467 15648 4477
rect 15614 4399 15648 4405
rect 15614 4331 15648 4333
rect 15614 4295 15648 4297
rect 15614 4223 15648 4229
rect 15614 4151 15648 4161
rect 15614 4079 15648 4093
rect 15614 4007 15648 4025
rect 14098 3896 14132 3915
rect 15614 3884 15648 3957
rect 15710 5895 15744 5996
rect 15710 5827 15744 5845
rect 15710 5759 15744 5773
rect 15710 5691 15744 5701
rect 15710 5623 15744 5629
rect 15710 5555 15744 5557
rect 15710 5519 15744 5521
rect 15710 5447 15744 5453
rect 15710 5375 15744 5385
rect 15710 5303 15744 5317
rect 16800 5479 22302 5500
rect 16800 5309 16848 5479
rect 22254 5309 22302 5479
rect 16800 5288 22302 5309
rect 23288 5477 28790 5498
rect 23288 5307 23336 5477
rect 28742 5307 28790 5477
rect 15710 5231 15744 5249
rect 16806 5208 22286 5288
rect 23288 5286 28790 5307
rect 15710 5159 15744 5181
rect 15710 5087 15744 5113
rect 15710 5015 15744 5045
rect 15710 4943 15744 4977
rect 15710 4875 15744 4909
rect 15710 4807 15744 4837
rect 15710 4739 15744 4765
rect 15710 4671 15744 4693
rect 15710 4603 15744 4621
rect 15710 4535 15744 4549
rect 15710 4467 15744 4477
rect 15710 4399 15744 4405
rect 15710 4331 15744 4333
rect 15710 4295 15744 4297
rect 15710 4223 15744 4229
rect 15710 4151 15744 4161
rect 16782 5196 22292 5208
rect 23302 5206 28782 5286
rect 16782 5174 17200 5196
rect 16782 5115 16816 5174
rect 16782 5043 16816 5055
rect 16782 4971 16816 4987
rect 16782 4899 16816 4919
rect 16782 4827 16816 4851
rect 16782 4755 16816 4783
rect 16782 4683 16816 4715
rect 16782 4613 16816 4647
rect 16782 4545 16816 4577
rect 16782 4477 16816 4505
rect 16782 4409 16816 4433
rect 16782 4341 16816 4361
rect 16782 4273 16816 4289
rect 16782 4205 16816 4217
rect 16782 4126 16816 4145
rect 16878 5115 16912 5134
rect 16878 5043 16912 5055
rect 16878 4971 16912 4987
rect 16878 4899 16912 4919
rect 16878 4827 16912 4851
rect 16878 4755 16912 4783
rect 16878 4683 16912 4715
rect 16878 4613 16912 4647
rect 16878 4545 16912 4577
rect 16878 4477 16912 4505
rect 16878 4409 16912 4433
rect 16878 4341 16912 4361
rect 16878 4273 16912 4289
rect 16878 4205 16912 4217
rect 15710 4079 15744 4093
rect 16878 4074 16912 4145
rect 16974 5115 17008 5174
rect 16974 5043 17008 5055
rect 16974 4971 17008 4987
rect 16974 4899 17008 4919
rect 16974 4827 17008 4851
rect 16974 4755 17008 4783
rect 16974 4683 17008 4715
rect 16974 4613 17008 4647
rect 16974 4545 17008 4577
rect 16974 4477 17008 4505
rect 16974 4409 17008 4433
rect 16974 4341 17008 4361
rect 16974 4273 17008 4289
rect 16974 4205 17008 4217
rect 16974 4126 17008 4145
rect 17070 5115 17104 5134
rect 17070 5043 17104 5055
rect 17070 4971 17104 4987
rect 17070 4899 17104 4919
rect 17070 4827 17104 4851
rect 17070 4755 17104 4783
rect 17070 4683 17104 4715
rect 17070 4613 17104 4647
rect 17070 4545 17104 4577
rect 17070 4477 17104 4505
rect 17070 4409 17104 4433
rect 17070 4341 17104 4361
rect 17070 4273 17104 4289
rect 17070 4205 17104 4217
rect 17070 4074 17104 4145
rect 17166 5115 17200 5174
rect 17470 5172 18464 5196
rect 17166 5043 17200 5055
rect 17166 4971 17200 4987
rect 17166 4899 17200 4919
rect 17166 4827 17200 4851
rect 17166 4755 17200 4783
rect 17166 4683 17200 4715
rect 17166 4613 17200 4647
rect 17166 4545 17200 4577
rect 17166 4477 17200 4505
rect 17166 4409 17200 4433
rect 17166 4341 17200 4361
rect 17166 4273 17200 4289
rect 17166 4205 17200 4217
rect 17166 4126 17200 4145
rect 17262 5115 17296 5134
rect 17262 5043 17296 5055
rect 17262 4971 17296 4987
rect 17262 4899 17296 4919
rect 17262 4827 17296 4851
rect 17262 4755 17296 4783
rect 17262 4683 17296 4715
rect 17262 4613 17296 4647
rect 17262 4545 17296 4577
rect 17262 4477 17296 4505
rect 17262 4409 17296 4433
rect 17262 4341 17296 4361
rect 17262 4273 17296 4289
rect 17262 4205 17296 4217
rect 17262 4074 17296 4145
rect 17470 5113 17504 5172
rect 17470 5041 17504 5053
rect 17470 4969 17504 4985
rect 17470 4897 17504 4917
rect 17470 4825 17504 4849
rect 17470 4753 17504 4781
rect 17470 4681 17504 4713
rect 17470 4611 17504 4645
rect 17470 4543 17504 4575
rect 17470 4475 17504 4503
rect 17470 4407 17504 4431
rect 17470 4339 17504 4359
rect 17470 4271 17504 4287
rect 17470 4203 17504 4215
rect 17470 4124 17504 4143
rect 17566 5113 17600 5132
rect 17566 5041 17600 5053
rect 17566 4969 17600 4985
rect 17566 4897 17600 4917
rect 17566 4825 17600 4849
rect 17566 4753 17600 4781
rect 17566 4681 17600 4713
rect 17566 4611 17600 4645
rect 17566 4543 17600 4575
rect 17566 4475 17600 4503
rect 17566 4407 17600 4431
rect 17566 4339 17600 4359
rect 17566 4271 17600 4287
rect 17566 4203 17600 4215
rect 16876 4040 17296 4074
rect 17566 4066 17600 4143
rect 17662 5113 17696 5172
rect 17662 5041 17696 5053
rect 17662 4969 17696 4985
rect 17662 4897 17696 4917
rect 17662 4825 17696 4849
rect 17662 4753 17696 4781
rect 17662 4681 17696 4713
rect 17662 4611 17696 4645
rect 17662 4543 17696 4575
rect 17662 4475 17696 4503
rect 17662 4407 17696 4431
rect 17662 4339 17696 4359
rect 17662 4271 17696 4287
rect 17662 4203 17696 4215
rect 17662 4124 17696 4143
rect 17758 5113 17792 5132
rect 17758 5041 17792 5053
rect 17758 4969 17792 4985
rect 17758 4897 17792 4917
rect 17758 4825 17792 4849
rect 17758 4753 17792 4781
rect 17758 4681 17792 4713
rect 17758 4611 17792 4645
rect 17758 4543 17792 4575
rect 17758 4475 17792 4503
rect 17758 4407 17792 4431
rect 17758 4339 17792 4359
rect 17758 4271 17792 4287
rect 17758 4203 17792 4215
rect 17758 4066 17792 4143
rect 17854 5113 17888 5172
rect 17854 5041 17888 5053
rect 17854 4969 17888 4985
rect 17854 4897 17888 4917
rect 17854 4825 17888 4849
rect 17854 4753 17888 4781
rect 17854 4681 17888 4713
rect 17854 4611 17888 4645
rect 17854 4543 17888 4575
rect 17854 4475 17888 4503
rect 17854 4407 17888 4431
rect 17854 4339 17888 4359
rect 17854 4271 17888 4287
rect 17854 4203 17888 4215
rect 17854 4124 17888 4143
rect 17950 5113 17984 5132
rect 17950 5041 17984 5053
rect 17950 4969 17984 4985
rect 17950 4897 17984 4917
rect 17950 4825 17984 4849
rect 17950 4753 17984 4781
rect 17950 4681 17984 4713
rect 17950 4611 17984 4645
rect 17950 4543 17984 4575
rect 17950 4475 17984 4503
rect 17950 4407 17984 4431
rect 17950 4339 17984 4359
rect 17950 4271 17984 4287
rect 17950 4203 17984 4215
rect 17950 4066 17984 4143
rect 18046 5113 18080 5172
rect 18046 5041 18080 5053
rect 18046 4969 18080 4985
rect 18046 4897 18080 4917
rect 18046 4825 18080 4849
rect 18046 4753 18080 4781
rect 18046 4681 18080 4713
rect 18046 4611 18080 4645
rect 18046 4543 18080 4575
rect 18046 4475 18080 4503
rect 18046 4407 18080 4431
rect 18046 4339 18080 4359
rect 18046 4271 18080 4287
rect 18046 4203 18080 4215
rect 18046 4124 18080 4143
rect 18142 5113 18176 5132
rect 18142 5041 18176 5053
rect 18142 4969 18176 4985
rect 18142 4897 18176 4917
rect 18142 4825 18176 4849
rect 18142 4753 18176 4781
rect 18142 4681 18176 4713
rect 18142 4611 18176 4645
rect 18142 4543 18176 4575
rect 18142 4475 18176 4503
rect 18142 4407 18176 4431
rect 18142 4339 18176 4359
rect 18142 4271 18176 4287
rect 18142 4203 18176 4215
rect 18142 4066 18176 4143
rect 18238 5113 18272 5172
rect 18238 5041 18272 5053
rect 18238 4969 18272 4985
rect 18238 4897 18272 4917
rect 18238 4825 18272 4849
rect 18238 4753 18272 4781
rect 18238 4681 18272 4713
rect 18238 4611 18272 4645
rect 18238 4543 18272 4575
rect 18238 4475 18272 4503
rect 18238 4407 18272 4431
rect 18238 4339 18272 4359
rect 18238 4271 18272 4287
rect 18238 4203 18272 4215
rect 18238 4124 18272 4143
rect 18334 5113 18368 5132
rect 18334 5041 18368 5053
rect 18334 4969 18368 4985
rect 18334 4897 18368 4917
rect 18334 4825 18368 4849
rect 18334 4753 18368 4781
rect 18334 4681 18368 4713
rect 18334 4611 18368 4645
rect 18334 4543 18368 4575
rect 18334 4475 18368 4503
rect 18334 4407 18368 4431
rect 18334 4339 18368 4359
rect 18334 4271 18368 4287
rect 18334 4203 18368 4215
rect 18334 4066 18368 4143
rect 18430 5113 18464 5172
rect 18430 5041 18464 5053
rect 18430 4969 18464 4985
rect 18430 4897 18464 4917
rect 18430 4825 18464 4849
rect 18430 4753 18464 4781
rect 18430 4681 18464 4713
rect 18430 4611 18464 4645
rect 18430 4543 18464 4575
rect 18430 4475 18464 4503
rect 18430 4407 18464 4431
rect 18430 4339 18464 4359
rect 18430 4271 18464 4287
rect 18430 4203 18464 4215
rect 18430 4124 18464 4143
rect 18674 5168 20052 5196
rect 18674 5107 18708 5168
rect 18674 5035 18708 5047
rect 18674 4963 18708 4979
rect 18674 4891 18708 4911
rect 18674 4819 18708 4843
rect 18674 4747 18708 4775
rect 18674 4675 18708 4707
rect 18674 4605 18708 4639
rect 18674 4537 18708 4569
rect 18674 4469 18708 4497
rect 18674 4401 18708 4425
rect 18674 4333 18708 4353
rect 18674 4265 18708 4281
rect 18674 4197 18708 4209
rect 18674 4118 18708 4137
rect 18770 5107 18804 5126
rect 18770 5035 18804 5047
rect 18770 4963 18804 4979
rect 18770 4891 18804 4911
rect 18770 4819 18804 4843
rect 18770 4747 18804 4775
rect 18770 4675 18804 4707
rect 18770 4605 18804 4639
rect 18770 4537 18804 4569
rect 18770 4469 18804 4497
rect 18770 4401 18804 4425
rect 18770 4333 18804 4353
rect 18770 4265 18804 4281
rect 18770 4197 18804 4209
rect 15710 4007 15744 4025
rect 15710 3922 15744 3957
rect 16814 3909 16830 3943
rect 16864 3909 16880 3943
rect 15614 3850 15744 3884
rect 7742 3727 7758 3761
rect 7792 3727 7808 3761
rect 10638 3725 10654 3759
rect 10688 3725 10704 3759
rect 10750 3736 10784 3832
rect 13810 3806 14036 3840
rect 10830 3725 10846 3759
rect 10880 3725 10896 3759
rect 13794 3699 13810 3733
rect 13844 3699 13860 3733
rect 13906 3710 13940 3806
rect 15550 3779 15616 3780
rect 15550 3745 15566 3779
rect 15600 3745 15616 3779
rect 15550 3744 15616 3745
rect 15710 3760 15744 3850
rect -4814 3677 -4780 3697
rect 13986 3699 14002 3733
rect 14036 3699 14052 3733
rect 16974 3821 17008 4040
rect 17566 4032 18368 4066
rect 18770 4060 18804 4137
rect 18866 5107 18900 5168
rect 18866 5035 18900 5047
rect 18866 4963 18900 4979
rect 18866 4891 18900 4911
rect 18866 4819 18900 4843
rect 18866 4747 18900 4775
rect 18866 4675 18900 4707
rect 18866 4605 18900 4639
rect 18866 4537 18900 4569
rect 18866 4469 18900 4497
rect 18866 4401 18900 4425
rect 18866 4333 18900 4353
rect 18866 4265 18900 4281
rect 18866 4197 18900 4209
rect 18866 4118 18900 4137
rect 18962 5107 18996 5126
rect 18962 5035 18996 5047
rect 18962 4963 18996 4979
rect 18962 4891 18996 4911
rect 18962 4819 18996 4843
rect 18962 4747 18996 4775
rect 18962 4675 18996 4707
rect 18962 4605 18996 4639
rect 18962 4537 18996 4569
rect 18962 4469 18996 4497
rect 18962 4401 18996 4425
rect 18962 4333 18996 4353
rect 18962 4265 18996 4281
rect 18962 4197 18996 4209
rect 18962 4060 18996 4137
rect 19058 5107 19092 5168
rect 19058 5035 19092 5047
rect 19058 4963 19092 4979
rect 19058 4891 19092 4911
rect 19058 4819 19092 4843
rect 19058 4747 19092 4775
rect 19058 4675 19092 4707
rect 19058 4605 19092 4639
rect 19058 4537 19092 4569
rect 19058 4469 19092 4497
rect 19058 4401 19092 4425
rect 19058 4333 19092 4353
rect 19058 4265 19092 4281
rect 19058 4197 19092 4209
rect 19058 4118 19092 4137
rect 19154 5107 19188 5126
rect 19154 5035 19188 5047
rect 19154 4963 19188 4979
rect 19154 4891 19188 4911
rect 19154 4819 19188 4843
rect 19154 4747 19188 4775
rect 19154 4675 19188 4707
rect 19154 4605 19188 4639
rect 19154 4537 19188 4569
rect 19154 4469 19188 4497
rect 19154 4401 19188 4425
rect 19154 4333 19188 4353
rect 19154 4265 19188 4281
rect 19154 4197 19188 4209
rect 19154 4060 19188 4137
rect 19250 5107 19284 5168
rect 19250 5035 19284 5047
rect 19250 4963 19284 4979
rect 19250 4891 19284 4911
rect 19250 4819 19284 4843
rect 19250 4747 19284 4775
rect 19250 4675 19284 4707
rect 19250 4605 19284 4639
rect 19250 4537 19284 4569
rect 19250 4469 19284 4497
rect 19250 4401 19284 4425
rect 19250 4333 19284 4353
rect 19250 4265 19284 4281
rect 19250 4197 19284 4209
rect 19250 4118 19284 4137
rect 19346 5107 19380 5126
rect 19346 5035 19380 5047
rect 19346 4963 19380 4979
rect 19346 4891 19380 4911
rect 19346 4819 19380 4843
rect 19346 4747 19380 4775
rect 19346 4675 19380 4707
rect 19346 4605 19380 4639
rect 19346 4537 19380 4569
rect 19346 4469 19380 4497
rect 19346 4401 19380 4425
rect 19346 4333 19380 4353
rect 19346 4265 19380 4281
rect 19346 4197 19380 4209
rect 19346 4060 19380 4137
rect 19442 5107 19476 5168
rect 19442 5035 19476 5047
rect 19442 4963 19476 4979
rect 19442 4891 19476 4911
rect 19442 4819 19476 4843
rect 19442 4747 19476 4775
rect 19442 4675 19476 4707
rect 19442 4605 19476 4639
rect 19442 4537 19476 4569
rect 19442 4469 19476 4497
rect 19442 4401 19476 4425
rect 19442 4333 19476 4353
rect 19442 4265 19476 4281
rect 19442 4197 19476 4209
rect 19442 4118 19476 4137
rect 19538 5107 19572 5126
rect 19538 5035 19572 5047
rect 19538 4963 19572 4979
rect 19538 4891 19572 4911
rect 19538 4819 19572 4843
rect 19538 4747 19572 4775
rect 19538 4675 19572 4707
rect 19538 4605 19572 4639
rect 19538 4537 19572 4569
rect 19538 4469 19572 4497
rect 19538 4401 19572 4425
rect 19538 4333 19572 4353
rect 19538 4265 19572 4281
rect 19538 4197 19572 4209
rect 19538 4060 19572 4137
rect 19634 5107 19668 5168
rect 19634 5035 19668 5047
rect 19634 4963 19668 4979
rect 19634 4891 19668 4911
rect 19634 4819 19668 4843
rect 19634 4747 19668 4775
rect 19634 4675 19668 4707
rect 19634 4605 19668 4639
rect 19634 4537 19668 4569
rect 19634 4469 19668 4497
rect 19634 4401 19668 4425
rect 19634 4333 19668 4353
rect 19634 4265 19668 4281
rect 19634 4197 19668 4209
rect 19634 4118 19668 4137
rect 19730 5107 19764 5126
rect 19730 5035 19764 5047
rect 19730 4963 19764 4979
rect 19730 4891 19764 4911
rect 19730 4819 19764 4843
rect 19730 4747 19764 4775
rect 19730 4675 19764 4707
rect 19730 4605 19764 4639
rect 19730 4537 19764 4569
rect 19730 4469 19764 4497
rect 19730 4401 19764 4425
rect 19730 4333 19764 4353
rect 19730 4265 19764 4281
rect 19730 4197 19764 4209
rect 19730 4060 19764 4137
rect 19826 5107 19860 5168
rect 19826 5035 19860 5047
rect 19826 4963 19860 4979
rect 19826 4891 19860 4911
rect 19826 4819 19860 4843
rect 19826 4747 19860 4775
rect 19826 4675 19860 4707
rect 19826 4605 19860 4639
rect 19826 4537 19860 4569
rect 19826 4469 19860 4497
rect 19826 4401 19860 4425
rect 19826 4333 19860 4353
rect 19826 4265 19860 4281
rect 19826 4197 19860 4209
rect 19826 4118 19860 4137
rect 19922 5107 19956 5126
rect 19922 5035 19956 5047
rect 19922 4963 19956 4979
rect 19922 4891 19956 4911
rect 19922 4819 19956 4843
rect 19922 4747 19956 4775
rect 19922 4675 19956 4707
rect 19922 4605 19956 4639
rect 19922 4537 19956 4569
rect 19922 4469 19956 4497
rect 19922 4401 19956 4425
rect 19922 4333 19956 4353
rect 19922 4265 19956 4281
rect 19922 4197 19956 4209
rect 19922 4060 19956 4137
rect 20018 5107 20052 5168
rect 20338 5174 22292 5196
rect 20018 5035 20052 5047
rect 20018 4963 20052 4979
rect 20018 4891 20052 4911
rect 20018 4819 20052 4843
rect 20018 4747 20052 4775
rect 20018 4675 20052 4707
rect 20018 4605 20052 4639
rect 20018 4537 20052 4569
rect 20018 4469 20052 4497
rect 20018 4401 20052 4425
rect 20018 4333 20052 4353
rect 20018 4265 20052 4281
rect 20018 4197 20052 4209
rect 20018 4118 20052 4137
rect 20114 5107 20148 5126
rect 20114 5035 20148 5047
rect 20114 4963 20148 4979
rect 20114 4891 20148 4911
rect 20114 4819 20148 4843
rect 20114 4747 20148 4775
rect 20114 4675 20148 4707
rect 20114 4605 20148 4639
rect 20114 4537 20148 4569
rect 20114 4469 20148 4497
rect 20114 4401 20148 4425
rect 20114 4333 20148 4353
rect 20114 4265 20148 4281
rect 20114 4197 20148 4209
rect 20114 4060 20148 4137
rect 20338 5101 20372 5174
rect 20338 5029 20372 5041
rect 20338 4957 20372 4973
rect 20338 4885 20372 4905
rect 20338 4813 20372 4837
rect 20338 4741 20372 4769
rect 20338 4669 20372 4701
rect 20338 4599 20372 4633
rect 20338 4531 20372 4563
rect 20338 4463 20372 4491
rect 20338 4395 20372 4419
rect 20338 4327 20372 4347
rect 20338 4259 20372 4275
rect 20338 4191 20372 4203
rect 20338 4112 20372 4131
rect 20434 5101 20468 5120
rect 20434 5029 20468 5041
rect 20434 4957 20468 4973
rect 20434 4885 20468 4905
rect 20434 4813 20468 4837
rect 20434 4741 20468 4769
rect 20434 4669 20468 4701
rect 20434 4599 20468 4633
rect 20434 4531 20468 4563
rect 20434 4463 20468 4491
rect 20434 4395 20468 4419
rect 20434 4327 20468 4347
rect 20434 4259 20468 4275
rect 20434 4191 20468 4203
rect 17502 3927 17518 3961
rect 17552 3927 17568 3961
rect 16814 3672 16830 3706
rect 16864 3672 16880 3706
rect -4814 3609 -4780 3625
rect 16974 3606 17008 3787
rect 17788 3819 17826 4032
rect 18770 4026 20148 4060
rect 20434 4066 20468 4131
rect 20530 5101 20564 5174
rect 20530 5029 20564 5041
rect 20530 4957 20564 4973
rect 20530 4885 20564 4905
rect 20530 4813 20564 4837
rect 20530 4741 20564 4769
rect 20530 4669 20564 4701
rect 20530 4599 20564 4633
rect 20530 4531 20564 4563
rect 20530 4463 20564 4491
rect 20530 4395 20564 4419
rect 20530 4327 20564 4347
rect 20530 4259 20564 4275
rect 20530 4191 20564 4203
rect 20530 4112 20564 4131
rect 20626 5101 20660 5120
rect 20626 5029 20660 5041
rect 20626 4957 20660 4973
rect 20626 4885 20660 4905
rect 20626 4813 20660 4837
rect 20626 4741 20660 4769
rect 20626 4669 20660 4701
rect 20626 4599 20660 4633
rect 20626 4531 20660 4563
rect 20626 4463 20660 4491
rect 20626 4395 20660 4419
rect 20626 4327 20660 4347
rect 20626 4259 20660 4275
rect 20626 4191 20660 4203
rect 20626 4066 20660 4131
rect 20722 5101 20756 5174
rect 20722 5029 20756 5041
rect 20722 4957 20756 4973
rect 20722 4885 20756 4905
rect 20722 4813 20756 4837
rect 20722 4741 20756 4769
rect 20722 4669 20756 4701
rect 20722 4599 20756 4633
rect 20722 4531 20756 4563
rect 20722 4463 20756 4491
rect 20722 4395 20756 4419
rect 20722 4327 20756 4347
rect 20722 4259 20756 4275
rect 20722 4191 20756 4203
rect 20722 4112 20756 4131
rect 20818 5101 20852 5120
rect 20818 5029 20852 5041
rect 20818 4957 20852 4973
rect 20818 4885 20852 4905
rect 20818 4813 20852 4837
rect 20818 4741 20852 4769
rect 20818 4669 20852 4701
rect 20818 4599 20852 4633
rect 20818 4531 20852 4563
rect 20818 4463 20852 4491
rect 20818 4395 20852 4419
rect 20818 4327 20852 4347
rect 20818 4259 20852 4275
rect 20818 4191 20852 4203
rect 20818 4066 20852 4131
rect 20914 5101 20948 5174
rect 20914 5029 20948 5041
rect 20914 4957 20948 4973
rect 20914 4885 20948 4905
rect 20914 4813 20948 4837
rect 20914 4741 20948 4769
rect 20914 4669 20948 4701
rect 20914 4599 20948 4633
rect 20914 4531 20948 4563
rect 20914 4463 20948 4491
rect 20914 4395 20948 4419
rect 20914 4327 20948 4347
rect 20914 4259 20948 4275
rect 20914 4191 20948 4203
rect 20914 4112 20948 4131
rect 21010 5101 21044 5120
rect 21010 5029 21044 5041
rect 21010 4957 21044 4973
rect 21010 4885 21044 4905
rect 21010 4813 21044 4837
rect 21010 4741 21044 4769
rect 21010 4669 21044 4701
rect 21010 4599 21044 4633
rect 21010 4531 21044 4563
rect 21010 4463 21044 4491
rect 21010 4395 21044 4419
rect 21010 4327 21044 4347
rect 21010 4259 21044 4275
rect 21010 4191 21044 4203
rect 21010 4066 21044 4131
rect 21106 5101 21140 5174
rect 21106 5029 21140 5041
rect 21106 4957 21140 4973
rect 21106 4885 21140 4905
rect 21106 4813 21140 4837
rect 21106 4741 21140 4769
rect 21106 4669 21140 4701
rect 21106 4599 21140 4633
rect 21106 4531 21140 4563
rect 21106 4463 21140 4491
rect 21106 4395 21140 4419
rect 21106 4327 21140 4347
rect 21106 4259 21140 4275
rect 21106 4191 21140 4203
rect 21106 4112 21140 4131
rect 21202 5101 21236 5120
rect 21202 5029 21236 5041
rect 21202 4957 21236 4973
rect 21202 4885 21236 4905
rect 21202 4813 21236 4837
rect 21202 4741 21236 4769
rect 21202 4669 21236 4701
rect 21202 4599 21236 4633
rect 21202 4531 21236 4563
rect 21202 4463 21236 4491
rect 21202 4395 21236 4419
rect 21202 4327 21236 4347
rect 21202 4259 21236 4275
rect 21202 4191 21236 4203
rect 21202 4066 21236 4131
rect 21298 5101 21332 5174
rect 21298 5029 21332 5041
rect 21298 4957 21332 4973
rect 21298 4885 21332 4905
rect 21298 4813 21332 4837
rect 21298 4741 21332 4769
rect 21298 4669 21332 4701
rect 21298 4599 21332 4633
rect 21298 4531 21332 4563
rect 21298 4463 21332 4491
rect 21298 4395 21332 4419
rect 21298 4327 21332 4347
rect 21298 4259 21332 4275
rect 21298 4191 21332 4203
rect 21298 4112 21332 4131
rect 21394 5101 21428 5120
rect 21394 5029 21428 5041
rect 21394 4957 21428 4973
rect 21394 4885 21428 4905
rect 21394 4813 21428 4837
rect 21394 4741 21428 4769
rect 21394 4669 21428 4701
rect 21394 4599 21428 4633
rect 21394 4531 21428 4563
rect 21394 4463 21428 4491
rect 21394 4395 21428 4419
rect 21394 4327 21428 4347
rect 21394 4259 21428 4275
rect 21394 4191 21428 4203
rect 21394 4066 21428 4131
rect 21490 5101 21524 5174
rect 21490 5029 21524 5041
rect 21490 4957 21524 4973
rect 21490 4885 21524 4905
rect 21490 4813 21524 4837
rect 21490 4741 21524 4769
rect 21490 4669 21524 4701
rect 21490 4599 21524 4633
rect 21490 4531 21524 4563
rect 21490 4463 21524 4491
rect 21490 4395 21524 4419
rect 21490 4327 21524 4347
rect 21490 4259 21524 4275
rect 21490 4191 21524 4203
rect 21490 4112 21524 4131
rect 21586 5101 21620 5120
rect 21586 5029 21620 5041
rect 21586 4957 21620 4973
rect 21586 4885 21620 4905
rect 21586 4813 21620 4837
rect 21586 4741 21620 4769
rect 21586 4669 21620 4701
rect 21586 4599 21620 4633
rect 21586 4531 21620 4563
rect 21586 4463 21620 4491
rect 21586 4395 21620 4419
rect 21586 4327 21620 4347
rect 21586 4259 21620 4275
rect 21586 4191 21620 4203
rect 21586 4066 21620 4131
rect 21682 5101 21716 5174
rect 21682 5029 21716 5041
rect 21682 4957 21716 4973
rect 21682 4885 21716 4905
rect 21682 4813 21716 4837
rect 21682 4741 21716 4769
rect 21682 4669 21716 4701
rect 21682 4599 21716 4633
rect 21682 4531 21716 4563
rect 21682 4463 21716 4491
rect 21682 4395 21716 4419
rect 21682 4327 21716 4347
rect 21682 4259 21716 4275
rect 21682 4191 21716 4203
rect 21682 4112 21716 4131
rect 21778 5101 21812 5120
rect 21778 5029 21812 5041
rect 21778 4957 21812 4973
rect 21778 4885 21812 4905
rect 21778 4813 21812 4837
rect 21778 4741 21812 4769
rect 21778 4669 21812 4701
rect 21778 4599 21812 4633
rect 21778 4531 21812 4563
rect 21778 4463 21812 4491
rect 21778 4395 21812 4419
rect 21778 4327 21812 4347
rect 21778 4259 21812 4275
rect 21778 4191 21812 4203
rect 21778 4066 21812 4131
rect 21874 5101 21908 5174
rect 21874 5029 21908 5041
rect 21874 4957 21908 4973
rect 21874 4885 21908 4905
rect 21874 4813 21908 4837
rect 21874 4741 21908 4769
rect 21874 4669 21908 4701
rect 21874 4599 21908 4633
rect 21874 4531 21908 4563
rect 21874 4463 21908 4491
rect 21874 4395 21908 4419
rect 21874 4327 21908 4347
rect 21874 4259 21908 4275
rect 21874 4191 21908 4203
rect 21874 4112 21908 4131
rect 21970 5101 22004 5120
rect 21970 5029 22004 5041
rect 21970 4957 22004 4973
rect 21970 4885 22004 4905
rect 21970 4813 22004 4837
rect 21970 4741 22004 4769
rect 21970 4669 22004 4701
rect 21970 4599 22004 4633
rect 21970 4531 22004 4563
rect 21970 4463 22004 4491
rect 21970 4395 22004 4419
rect 21970 4327 22004 4347
rect 21970 4259 22004 4275
rect 21970 4191 22004 4203
rect 21970 4066 22004 4131
rect 22066 5101 22100 5174
rect 22066 5029 22100 5041
rect 22066 4957 22100 4973
rect 22066 4885 22100 4905
rect 22066 4813 22100 4837
rect 22066 4741 22100 4769
rect 22066 4669 22100 4701
rect 22066 4599 22100 4633
rect 22066 4531 22100 4563
rect 22066 4463 22100 4491
rect 22066 4395 22100 4419
rect 22066 4327 22100 4347
rect 22066 4259 22100 4275
rect 22066 4191 22100 4203
rect 22066 4112 22100 4131
rect 22162 5101 22196 5120
rect 22162 5029 22196 5041
rect 22162 4957 22196 4973
rect 22162 4885 22196 4905
rect 22162 4813 22196 4837
rect 22162 4741 22196 4769
rect 22162 4669 22196 4701
rect 22162 4599 22196 4633
rect 22162 4531 22196 4563
rect 22162 4463 22196 4491
rect 22162 4395 22196 4419
rect 22162 4327 22196 4347
rect 22162 4259 22196 4275
rect 22162 4191 22196 4203
rect 22162 4066 22196 4131
rect 22258 5101 22292 5174
rect 22258 5029 22292 5041
rect 22258 4957 22292 4973
rect 22258 4885 22292 4905
rect 22258 4813 22292 4837
rect 22258 4741 22292 4769
rect 22258 4669 22292 4701
rect 22258 4599 22292 4633
rect 22258 4531 22292 4563
rect 22258 4463 22292 4491
rect 22258 4395 22292 4419
rect 22258 4327 22292 4347
rect 22258 4259 22292 4275
rect 22258 4191 22292 4203
rect 22258 4112 22292 4131
rect 23270 5194 28782 5206
rect 23270 5172 23688 5194
rect 23270 5113 23304 5172
rect 23270 5041 23304 5053
rect 23270 4969 23304 4985
rect 23270 4897 23304 4917
rect 23270 4825 23304 4849
rect 23270 4753 23304 4781
rect 23270 4681 23304 4713
rect 23270 4611 23304 4645
rect 23270 4543 23304 4575
rect 23270 4475 23304 4503
rect 23270 4407 23304 4431
rect 23270 4339 23304 4359
rect 23270 4271 23304 4287
rect 23270 4203 23304 4215
rect 23270 4124 23304 4143
rect 23366 5113 23400 5132
rect 23366 5041 23400 5053
rect 23366 4969 23400 4985
rect 23366 4897 23400 4917
rect 23366 4825 23400 4849
rect 23366 4753 23400 4781
rect 23366 4681 23400 4713
rect 23366 4611 23400 4645
rect 23366 4543 23400 4575
rect 23366 4475 23400 4503
rect 23366 4407 23400 4431
rect 23366 4339 23400 4359
rect 23366 4271 23400 4287
rect 23366 4203 23400 4215
rect 23366 4072 23400 4143
rect 23462 5113 23496 5172
rect 23462 5041 23496 5053
rect 23462 4969 23496 4985
rect 23462 4897 23496 4917
rect 23462 4825 23496 4849
rect 23462 4753 23496 4781
rect 23462 4681 23496 4713
rect 23462 4611 23496 4645
rect 23462 4543 23496 4575
rect 23462 4475 23496 4503
rect 23462 4407 23496 4431
rect 23462 4339 23496 4359
rect 23462 4271 23496 4287
rect 23462 4203 23496 4215
rect 23462 4124 23496 4143
rect 23558 5113 23592 5132
rect 23558 5041 23592 5053
rect 23558 4969 23592 4985
rect 23558 4897 23592 4917
rect 23558 4825 23592 4849
rect 23558 4753 23592 4781
rect 23558 4681 23592 4713
rect 23558 4611 23592 4645
rect 23558 4543 23592 4575
rect 23558 4475 23592 4503
rect 23558 4407 23592 4431
rect 23558 4339 23592 4359
rect 23558 4271 23592 4287
rect 23558 4203 23592 4215
rect 23558 4072 23592 4143
rect 23654 5113 23688 5172
rect 23958 5170 24952 5194
rect 23654 5041 23688 5053
rect 23654 4969 23688 4985
rect 23654 4897 23688 4917
rect 23654 4825 23688 4849
rect 23654 4753 23688 4781
rect 23654 4681 23688 4713
rect 23654 4611 23688 4645
rect 23654 4543 23688 4575
rect 23654 4475 23688 4503
rect 23654 4407 23688 4431
rect 23654 4339 23688 4359
rect 23654 4271 23688 4287
rect 23654 4203 23688 4215
rect 23654 4124 23688 4143
rect 23750 5113 23784 5132
rect 23750 5041 23784 5053
rect 23750 4969 23784 4985
rect 23750 4897 23784 4917
rect 23750 4825 23784 4849
rect 23750 4753 23784 4781
rect 23750 4681 23784 4713
rect 23750 4611 23784 4645
rect 23750 4543 23784 4575
rect 23750 4475 23784 4503
rect 23750 4407 23784 4431
rect 23750 4339 23784 4359
rect 23750 4271 23784 4287
rect 23750 4203 23784 4215
rect 23750 4072 23784 4143
rect 23958 5111 23992 5170
rect 23958 5039 23992 5051
rect 23958 4967 23992 4983
rect 23958 4895 23992 4915
rect 23958 4823 23992 4847
rect 23958 4751 23992 4779
rect 23958 4679 23992 4711
rect 23958 4609 23992 4643
rect 23958 4541 23992 4573
rect 23958 4473 23992 4501
rect 23958 4405 23992 4429
rect 23958 4337 23992 4357
rect 23958 4269 23992 4285
rect 23958 4201 23992 4213
rect 23958 4122 23992 4141
rect 24054 5111 24088 5130
rect 24054 5039 24088 5051
rect 24054 4967 24088 4983
rect 24054 4895 24088 4915
rect 24054 4823 24088 4847
rect 24054 4751 24088 4779
rect 24054 4679 24088 4711
rect 24054 4609 24088 4643
rect 24054 4541 24088 4573
rect 24054 4473 24088 4501
rect 24054 4405 24088 4429
rect 24054 4337 24088 4357
rect 24054 4269 24088 4285
rect 24054 4201 24088 4213
rect 20434 4032 22196 4066
rect 23364 4038 23784 4072
rect 24054 4064 24088 4141
rect 24150 5111 24184 5170
rect 24150 5039 24184 5051
rect 24150 4967 24184 4983
rect 24150 4895 24184 4915
rect 24150 4823 24184 4847
rect 24150 4751 24184 4779
rect 24150 4679 24184 4711
rect 24150 4609 24184 4643
rect 24150 4541 24184 4573
rect 24150 4473 24184 4501
rect 24150 4405 24184 4429
rect 24150 4337 24184 4357
rect 24150 4269 24184 4285
rect 24150 4201 24184 4213
rect 24150 4122 24184 4141
rect 24246 5111 24280 5130
rect 24246 5039 24280 5051
rect 24246 4967 24280 4983
rect 24246 4895 24280 4915
rect 24246 4823 24280 4847
rect 24246 4751 24280 4779
rect 24246 4679 24280 4711
rect 24246 4609 24280 4643
rect 24246 4541 24280 4573
rect 24246 4473 24280 4501
rect 24246 4405 24280 4429
rect 24246 4337 24280 4357
rect 24246 4269 24280 4285
rect 24246 4201 24280 4213
rect 24246 4064 24280 4141
rect 24342 5111 24376 5170
rect 24342 5039 24376 5051
rect 24342 4967 24376 4983
rect 24342 4895 24376 4915
rect 24342 4823 24376 4847
rect 24342 4751 24376 4779
rect 24342 4679 24376 4711
rect 24342 4609 24376 4643
rect 24342 4541 24376 4573
rect 24342 4473 24376 4501
rect 24342 4405 24376 4429
rect 24342 4337 24376 4357
rect 24342 4269 24376 4285
rect 24342 4201 24376 4213
rect 24342 4122 24376 4141
rect 24438 5111 24472 5130
rect 24438 5039 24472 5051
rect 24438 4967 24472 4983
rect 24438 4895 24472 4915
rect 24438 4823 24472 4847
rect 24438 4751 24472 4779
rect 24438 4679 24472 4711
rect 24438 4609 24472 4643
rect 24438 4541 24472 4573
rect 24438 4473 24472 4501
rect 24438 4405 24472 4429
rect 24438 4337 24472 4357
rect 24438 4269 24472 4285
rect 24438 4201 24472 4213
rect 24438 4064 24472 4141
rect 24534 5111 24568 5170
rect 24534 5039 24568 5051
rect 24534 4967 24568 4983
rect 24534 4895 24568 4915
rect 24534 4823 24568 4847
rect 24534 4751 24568 4779
rect 24534 4679 24568 4711
rect 24534 4609 24568 4643
rect 24534 4541 24568 4573
rect 24534 4473 24568 4501
rect 24534 4405 24568 4429
rect 24534 4337 24568 4357
rect 24534 4269 24568 4285
rect 24534 4201 24568 4213
rect 24534 4122 24568 4141
rect 24630 5111 24664 5130
rect 24630 5039 24664 5051
rect 24630 4967 24664 4983
rect 24630 4895 24664 4915
rect 24630 4823 24664 4847
rect 24630 4751 24664 4779
rect 24630 4679 24664 4711
rect 24630 4609 24664 4643
rect 24630 4541 24664 4573
rect 24630 4473 24664 4501
rect 24630 4405 24664 4429
rect 24630 4337 24664 4357
rect 24630 4269 24664 4285
rect 24630 4201 24664 4213
rect 24630 4064 24664 4141
rect 24726 5111 24760 5170
rect 24726 5039 24760 5051
rect 24726 4967 24760 4983
rect 24726 4895 24760 4915
rect 24726 4823 24760 4847
rect 24726 4751 24760 4779
rect 24726 4679 24760 4711
rect 24726 4609 24760 4643
rect 24726 4541 24760 4573
rect 24726 4473 24760 4501
rect 24726 4405 24760 4429
rect 24726 4337 24760 4357
rect 24726 4269 24760 4285
rect 24726 4201 24760 4213
rect 24726 4122 24760 4141
rect 24822 5111 24856 5130
rect 24822 5039 24856 5051
rect 24822 4967 24856 4983
rect 24822 4895 24856 4915
rect 24822 4823 24856 4847
rect 24822 4751 24856 4779
rect 24822 4679 24856 4711
rect 24822 4609 24856 4643
rect 24822 4541 24856 4573
rect 24822 4473 24856 4501
rect 24822 4405 24856 4429
rect 24822 4337 24856 4357
rect 24822 4269 24856 4285
rect 24822 4201 24856 4213
rect 24822 4064 24856 4141
rect 24918 5111 24952 5170
rect 24918 5039 24952 5051
rect 24918 4967 24952 4983
rect 24918 4895 24952 4915
rect 24918 4823 24952 4847
rect 24918 4751 24952 4779
rect 24918 4679 24952 4711
rect 24918 4609 24952 4643
rect 24918 4541 24952 4573
rect 24918 4473 24952 4501
rect 24918 4405 24952 4429
rect 24918 4337 24952 4357
rect 24918 4269 24952 4285
rect 24918 4201 24952 4213
rect 24918 4122 24952 4141
rect 25162 5166 26540 5194
rect 25162 5105 25196 5166
rect 25162 5033 25196 5045
rect 25162 4961 25196 4977
rect 25162 4889 25196 4909
rect 25162 4817 25196 4841
rect 25162 4745 25196 4773
rect 25162 4673 25196 4705
rect 25162 4603 25196 4637
rect 25162 4535 25196 4567
rect 25162 4467 25196 4495
rect 25162 4399 25196 4423
rect 25162 4331 25196 4351
rect 25162 4263 25196 4279
rect 25162 4195 25196 4207
rect 25162 4116 25196 4135
rect 25258 5105 25292 5124
rect 25258 5033 25292 5045
rect 25258 4961 25292 4977
rect 25258 4889 25292 4909
rect 25258 4817 25292 4841
rect 25258 4745 25292 4773
rect 25258 4673 25292 4705
rect 25258 4603 25292 4637
rect 25258 4535 25292 4567
rect 25258 4467 25292 4495
rect 25258 4399 25292 4423
rect 25258 4331 25292 4351
rect 25258 4263 25292 4279
rect 25258 4195 25292 4207
rect 18706 3921 18722 3955
rect 18756 3921 18772 3955
rect 17788 3785 17790 3819
rect 17824 3785 17826 3819
rect 17506 3702 17522 3736
rect 17556 3702 17572 3736
rect 17788 3616 17826 3785
rect 19440 3806 19480 4026
rect 20370 3915 20386 3949
rect 20420 3915 20436 3949
rect 19440 3772 19443 3806
rect 19477 3772 19480 3806
rect 18704 3658 18720 3692
rect 18754 3658 18770 3692
rect -4814 3541 -4780 3553
rect 16782 3572 17200 3606
rect -4814 3462 -4780 3481
rect 16686 3519 16720 3538
rect 16686 3447 16720 3459
rect -5294 3376 -4874 3410
rect -1606 3394 -1590 3428
rect -1556 3394 -1540 3428
rect -8434 3251 -8418 3285
rect -8384 3251 -8368 3285
rect -9684 3106 -9678 3140
rect -9644 3106 -9638 3140
rect -11344 3010 -11328 3044
rect -11294 3010 -11278 3044
rect -13170 2771 -13136 2783
rect -13170 2699 -13136 2715
rect -13170 2627 -13136 2647
rect -13170 2555 -13136 2579
rect -13170 2483 -13136 2511
rect -13170 2411 -13136 2443
rect -13170 2341 -13136 2375
rect -13170 2273 -13136 2305
rect -13170 2205 -13136 2233
rect -13170 2137 -13136 2161
rect -13170 2069 -13136 2089
rect -13170 2001 -13136 2017
rect -13170 1933 -13136 1945
rect -13170 1854 -13136 1873
rect -13074 2843 -13040 2862
rect -13074 2771 -13040 2783
rect -13074 2699 -13040 2715
rect -13074 2627 -13040 2647
rect -13074 2555 -13040 2579
rect -13074 2483 -13040 2511
rect -13074 2411 -13040 2443
rect -13074 2341 -13040 2375
rect -13074 2273 -13040 2305
rect -13074 2205 -13040 2233
rect -13074 2137 -13040 2161
rect -13074 2069 -13040 2089
rect -13074 2001 -13040 2017
rect -13074 1933 -13040 1945
rect -13074 1812 -13040 1873
rect -14430 1798 -13040 1812
rect -12836 2847 -12802 2866
rect -12836 2775 -12802 2787
rect -12836 2703 -12802 2719
rect -12836 2631 -12802 2651
rect -12836 2559 -12802 2583
rect -12836 2487 -12802 2515
rect -12836 2415 -12802 2447
rect -12836 2345 -12802 2379
rect -12836 2277 -12802 2309
rect -12836 2209 -12802 2237
rect -12836 2141 -12802 2165
rect -12836 2073 -12802 2093
rect -12836 2005 -12802 2021
rect -12836 1937 -12802 1949
rect -12836 1824 -12802 1877
rect -12740 2847 -12706 2920
rect -12740 2775 -12706 2787
rect -12740 2703 -12706 2719
rect -12740 2631 -12706 2651
rect -12740 2559 -12706 2583
rect -12740 2487 -12706 2515
rect -12740 2415 -12706 2447
rect -12740 2345 -12706 2379
rect -12740 2277 -12706 2309
rect -12740 2209 -12706 2237
rect -12740 2141 -12706 2165
rect -12740 2073 -12706 2093
rect -12740 2005 -12706 2021
rect -12740 1937 -12706 1949
rect -12740 1858 -12706 1877
rect -12644 2847 -12610 2866
rect -12644 2775 -12610 2787
rect -12644 2703 -12610 2719
rect -12644 2631 -12610 2651
rect -12644 2559 -12610 2583
rect -12644 2487 -12610 2515
rect -12644 2415 -12610 2447
rect -12644 2345 -12610 2379
rect -12644 2277 -12610 2309
rect -12644 2209 -12610 2237
rect -12644 2141 -12610 2165
rect -12644 2073 -12610 2093
rect -12644 2005 -12610 2021
rect -12644 1937 -12610 1949
rect -12644 1824 -12610 1877
rect -12548 2847 -12514 2920
rect -12548 2775 -12514 2787
rect -12548 2703 -12514 2719
rect -12548 2631 -12514 2651
rect -12548 2559 -12514 2583
rect -12548 2487 -12514 2515
rect -12548 2415 -12514 2447
rect -12548 2345 -12514 2379
rect -12548 2277 -12514 2309
rect -12548 2209 -12514 2237
rect -12548 2141 -12514 2165
rect -12548 2073 -12514 2093
rect -12548 2005 -12514 2021
rect -12548 1937 -12514 1949
rect -12548 1858 -12514 1877
rect -12452 2847 -12418 2866
rect -12452 2775 -12418 2787
rect -12452 2703 -12418 2719
rect -12452 2631 -12418 2651
rect -12452 2559 -12418 2583
rect -12452 2487 -12418 2515
rect -12452 2415 -12418 2447
rect -12452 2345 -12418 2379
rect -12452 2277 -12418 2309
rect -12452 2209 -12418 2237
rect -12452 2141 -12418 2165
rect -12452 2073 -12418 2093
rect -12452 2005 -12418 2021
rect -12452 1937 -12418 1949
rect -12452 1824 -12418 1877
rect -12356 2847 -12322 2920
rect -12356 2775 -12322 2787
rect -12356 2703 -12322 2719
rect -12356 2631 -12322 2651
rect -12356 2559 -12322 2583
rect -12356 2487 -12322 2515
rect -12356 2415 -12322 2447
rect -12356 2345 -12322 2379
rect -12356 2277 -12322 2309
rect -12356 2209 -12322 2237
rect -12356 2141 -12322 2165
rect -12356 2073 -12322 2093
rect -12356 2005 -12322 2021
rect -12356 1937 -12322 1949
rect -12356 1858 -12322 1877
rect -12260 2847 -12226 2866
rect -12260 2775 -12226 2787
rect -12260 2703 -12226 2719
rect -12260 2631 -12226 2651
rect -12260 2559 -12226 2583
rect -12260 2487 -12226 2515
rect -12260 2415 -12226 2447
rect -12260 2345 -12226 2379
rect -12260 2277 -12226 2309
rect -12260 2209 -12226 2237
rect -12260 2141 -12226 2165
rect -12260 2073 -12226 2093
rect -12260 2005 -12226 2021
rect -12260 1937 -12226 1949
rect -12260 1824 -12226 1877
rect -12164 2847 -12130 2920
rect -12164 2775 -12130 2787
rect -12164 2703 -12130 2719
rect -12164 2631 -12130 2651
rect -12164 2559 -12130 2583
rect -12164 2487 -12130 2515
rect -12164 2415 -12130 2447
rect -12164 2345 -12130 2379
rect -12164 2277 -12130 2309
rect -12164 2209 -12130 2237
rect -12164 2141 -12130 2165
rect -12164 2073 -12130 2093
rect -12164 2005 -12130 2021
rect -12164 1937 -12130 1949
rect -12164 1858 -12130 1877
rect -12068 2847 -12034 2866
rect -12068 2775 -12034 2787
rect -12068 2703 -12034 2719
rect -12068 2631 -12034 2651
rect -12068 2559 -12034 2583
rect -12068 2487 -12034 2515
rect -12068 2415 -12034 2447
rect -12068 2345 -12034 2379
rect -12068 2277 -12034 2309
rect -12068 2209 -12034 2237
rect -12068 2141 -12034 2165
rect -12068 2073 -12034 2093
rect -12068 2005 -12034 2021
rect -12068 1937 -12034 1949
rect -12068 1824 -12034 1877
rect -11972 2847 -11938 2920
rect -11664 2910 -11246 2944
rect -9684 2940 -9638 3106
rect -7478 3142 -7438 3362
rect -6770 3257 -6754 3291
rect -6720 3257 -6704 3291
rect -7478 3108 -7475 3142
rect -7441 3108 -7438 3142
rect -8436 2992 -8420 3026
rect -8386 2992 -8370 3026
rect -7478 2944 -7438 3108
rect -5824 3155 -5786 3368
rect -5566 3263 -5550 3297
rect -5516 3263 -5500 3297
rect -5824 3121 -5822 3155
rect -5788 3121 -5786 3155
rect -6768 2994 -6752 3028
rect -6718 2994 -6702 3028
rect -5824 2952 -5786 3121
rect -5006 3157 -4972 3376
rect 16686 3375 16720 3391
rect -1590 3290 -1110 3324
rect -1076 3290 -980 3324
rect -4878 3245 -4862 3279
rect -4828 3245 -4812 3279
rect -5570 3038 -5554 3072
rect -5520 3038 -5504 3072
rect -11972 2775 -11938 2787
rect -11972 2703 -11938 2719
rect -11972 2631 -11938 2651
rect -11972 2559 -11938 2583
rect -11972 2487 -11938 2515
rect -11972 2415 -11938 2447
rect -11972 2345 -11938 2379
rect -11972 2277 -11938 2309
rect -11972 2209 -11938 2237
rect -11972 2141 -11938 2165
rect -11972 2073 -11938 2093
rect -11972 2005 -11938 2021
rect -11972 1937 -11938 1949
rect -11972 1858 -11938 1877
rect -11876 2847 -11842 2866
rect -11876 2775 -11842 2787
rect -11876 2703 -11842 2719
rect -11876 2631 -11842 2651
rect -11876 2559 -11842 2583
rect -11876 2487 -11842 2515
rect -11876 2415 -11842 2447
rect -11876 2345 -11842 2379
rect -11876 2277 -11842 2309
rect -11876 2209 -11842 2237
rect -11876 2141 -11842 2165
rect -11876 2073 -11842 2093
rect -11876 2005 -11842 2021
rect -11876 1937 -11842 1949
rect -11876 1824 -11842 1877
rect -11664 2857 -11630 2910
rect -11664 2785 -11630 2797
rect -11664 2713 -11630 2729
rect -11664 2641 -11630 2661
rect -11664 2569 -11630 2593
rect -11664 2497 -11630 2525
rect -11664 2425 -11630 2457
rect -11664 2355 -11630 2389
rect -11664 2287 -11630 2319
rect -11664 2219 -11630 2247
rect -11664 2151 -11630 2175
rect -11664 2083 -11630 2103
rect -11664 2015 -11630 2031
rect -11664 1947 -11630 1959
rect -11664 1868 -11630 1887
rect -11568 2857 -11534 2876
rect -11568 2785 -11534 2797
rect -11568 2713 -11534 2729
rect -11568 2641 -11534 2661
rect -11568 2569 -11534 2593
rect -11568 2497 -11534 2525
rect -11568 2425 -11534 2457
rect -11568 2355 -11534 2389
rect -11568 2287 -11534 2319
rect -11568 2219 -11534 2247
rect -11568 2151 -11534 2175
rect -11568 2083 -11534 2103
rect -11568 2015 -11534 2031
rect -11568 1947 -11534 1959
rect -12836 1798 -11842 1824
rect -11568 1820 -11534 1887
rect -11472 2857 -11438 2910
rect -11472 2785 -11438 2797
rect -11472 2713 -11438 2729
rect -11472 2641 -11438 2661
rect -11472 2569 -11438 2593
rect -11472 2497 -11438 2525
rect -11472 2425 -11438 2457
rect -11472 2355 -11438 2389
rect -11472 2287 -11438 2319
rect -11472 2219 -11438 2247
rect -11472 2151 -11438 2175
rect -11472 2083 -11438 2103
rect -11472 2015 -11438 2031
rect -11472 1947 -11438 1959
rect -11472 1868 -11438 1887
rect -11376 2857 -11342 2876
rect -11376 2785 -11342 2797
rect -11376 2713 -11342 2729
rect -11376 2641 -11342 2661
rect -11376 2569 -11342 2593
rect -11376 2497 -11342 2525
rect -11376 2425 -11342 2457
rect -11376 2355 -11342 2389
rect -11376 2287 -11342 2319
rect -11376 2219 -11342 2247
rect -11376 2151 -11342 2175
rect -11376 2083 -11342 2103
rect -11376 2015 -11342 2031
rect -11376 1947 -11342 1959
rect -11376 1820 -11342 1887
rect -11280 2857 -11246 2910
rect -10102 2906 -8338 2940
rect -11280 2785 -11246 2797
rect -11280 2713 -11246 2729
rect -11280 2641 -11246 2661
rect -11280 2569 -11246 2593
rect -11280 2497 -11246 2525
rect -11280 2425 -11246 2457
rect -11280 2355 -11246 2389
rect -11280 2287 -11246 2319
rect -11280 2219 -11246 2247
rect -11280 2151 -11246 2175
rect -11280 2083 -11246 2103
rect -11280 2015 -11246 2031
rect -11280 1947 -11246 1959
rect -11280 1868 -11246 1887
rect -11184 2857 -11150 2876
rect -11184 2785 -11150 2797
rect -11184 2713 -11150 2729
rect -11184 2641 -11150 2661
rect -11184 2569 -11150 2593
rect -11184 2497 -11150 2525
rect -11184 2425 -11150 2457
rect -11184 2355 -11150 2389
rect -11184 2287 -11150 2319
rect -11184 2219 -11150 2247
rect -11184 2151 -11150 2175
rect -11184 2083 -11150 2103
rect -11184 2015 -11150 2031
rect -11184 1947 -11150 1959
rect -11184 1820 -11150 1887
rect -11568 1798 -11150 1820
rect -16662 1786 -11150 1798
rect -10196 2849 -10162 2868
rect -10196 2777 -10162 2789
rect -10196 2705 -10162 2721
rect -10196 2633 -10162 2653
rect -10196 2561 -10162 2585
rect -10196 2489 -10162 2517
rect -10196 2417 -10162 2449
rect -10196 2347 -10162 2381
rect -10196 2279 -10162 2311
rect -10196 2211 -10162 2239
rect -10196 2143 -10162 2167
rect -10196 2075 -10162 2095
rect -10196 2007 -10162 2023
rect -10196 1939 -10162 1951
rect -10196 1818 -10162 1879
rect -10100 2849 -10066 2906
rect -10100 2777 -10066 2789
rect -10100 2705 -10066 2721
rect -10100 2633 -10066 2653
rect -10100 2561 -10066 2585
rect -10100 2489 -10066 2517
rect -10100 2417 -10066 2449
rect -10100 2347 -10066 2381
rect -10100 2279 -10066 2311
rect -10100 2211 -10066 2239
rect -10100 2143 -10066 2167
rect -10100 2075 -10066 2095
rect -10100 2007 -10066 2023
rect -10100 1939 -10066 1951
rect -10100 1860 -10066 1879
rect -10004 2849 -9970 2868
rect -10004 2777 -9970 2789
rect -10004 2705 -9970 2721
rect -10004 2633 -9970 2653
rect -10004 2561 -9970 2585
rect -10004 2489 -9970 2517
rect -10004 2417 -9970 2449
rect -10004 2347 -9970 2381
rect -10004 2279 -9970 2311
rect -10004 2211 -9970 2239
rect -10004 2143 -9970 2167
rect -10004 2075 -9970 2095
rect -10004 2007 -9970 2023
rect -10004 1939 -9970 1951
rect -10004 1818 -9970 1879
rect -9908 2849 -9874 2906
rect -9908 2777 -9874 2789
rect -9908 2705 -9874 2721
rect -9908 2633 -9874 2653
rect -9908 2561 -9874 2585
rect -9908 2489 -9874 2517
rect -9908 2417 -9874 2449
rect -9908 2347 -9874 2381
rect -9908 2279 -9874 2311
rect -9908 2211 -9874 2239
rect -9908 2143 -9874 2167
rect -9908 2075 -9874 2095
rect -9908 2007 -9874 2023
rect -9908 1939 -9874 1951
rect -9908 1860 -9874 1879
rect -9812 2849 -9778 2868
rect -9812 2777 -9778 2789
rect -9812 2705 -9778 2721
rect -9812 2633 -9778 2653
rect -9812 2561 -9778 2585
rect -9812 2489 -9778 2517
rect -9812 2417 -9778 2449
rect -9812 2347 -9778 2381
rect -9812 2279 -9778 2311
rect -9812 2211 -9778 2239
rect -9812 2143 -9778 2167
rect -9812 2075 -9778 2095
rect -9812 2007 -9778 2023
rect -9812 1939 -9778 1951
rect -9812 1818 -9778 1879
rect -9716 2849 -9682 2906
rect -9716 2777 -9682 2789
rect -9716 2705 -9682 2721
rect -9716 2633 -9682 2653
rect -9716 2561 -9682 2585
rect -9716 2489 -9682 2517
rect -9716 2417 -9682 2449
rect -9716 2347 -9682 2381
rect -9716 2279 -9682 2311
rect -9716 2211 -9682 2239
rect -9716 2143 -9682 2167
rect -9716 2075 -9682 2095
rect -9716 2007 -9682 2023
rect -9716 1939 -9682 1951
rect -9716 1860 -9682 1879
rect -9620 2849 -9586 2868
rect -9620 2777 -9586 2789
rect -9620 2705 -9586 2721
rect -9620 2633 -9586 2653
rect -9620 2561 -9586 2585
rect -9620 2489 -9586 2517
rect -9620 2417 -9586 2449
rect -9620 2347 -9586 2381
rect -9620 2279 -9586 2311
rect -9620 2211 -9586 2239
rect -9620 2143 -9586 2167
rect -9620 2075 -9586 2095
rect -9620 2007 -9586 2023
rect -9620 1939 -9586 1951
rect -9620 1818 -9586 1879
rect -9524 2849 -9490 2906
rect -9524 2777 -9490 2789
rect -9524 2705 -9490 2721
rect -9524 2633 -9490 2653
rect -9524 2561 -9490 2585
rect -9524 2489 -9490 2517
rect -9524 2417 -9490 2449
rect -9524 2347 -9490 2381
rect -9524 2279 -9490 2311
rect -9524 2211 -9490 2239
rect -9524 2143 -9490 2167
rect -9524 2075 -9490 2095
rect -9524 2007 -9490 2023
rect -9524 1939 -9490 1951
rect -9524 1860 -9490 1879
rect -9428 2849 -9394 2868
rect -9428 2777 -9394 2789
rect -9428 2705 -9394 2721
rect -9428 2633 -9394 2653
rect -9428 2561 -9394 2585
rect -9428 2489 -9394 2517
rect -9428 2417 -9394 2449
rect -9428 2347 -9394 2381
rect -9428 2279 -9394 2311
rect -9428 2211 -9394 2239
rect -9428 2143 -9394 2167
rect -9428 2075 -9394 2095
rect -9428 2007 -9394 2023
rect -9428 1939 -9394 1951
rect -9428 1818 -9394 1879
rect -9332 2849 -9298 2906
rect -9332 2777 -9298 2789
rect -9332 2705 -9298 2721
rect -9332 2633 -9298 2653
rect -9332 2561 -9298 2585
rect -9332 2489 -9298 2517
rect -9332 2417 -9298 2449
rect -9332 2347 -9298 2381
rect -9332 2279 -9298 2311
rect -9332 2211 -9298 2239
rect -9332 2143 -9298 2167
rect -9332 2075 -9298 2095
rect -9332 2007 -9298 2023
rect -9332 1939 -9298 1951
rect -9332 1860 -9298 1879
rect -9236 2849 -9202 2868
rect -9236 2777 -9202 2789
rect -9236 2705 -9202 2721
rect -9236 2633 -9202 2653
rect -9236 2561 -9202 2585
rect -9236 2489 -9202 2517
rect -9236 2417 -9202 2449
rect -9236 2347 -9202 2381
rect -9236 2279 -9202 2311
rect -9236 2211 -9202 2239
rect -9236 2143 -9202 2167
rect -9236 2075 -9202 2095
rect -9236 2007 -9202 2023
rect -9236 1939 -9202 1951
rect -9236 1818 -9202 1879
rect -9140 2849 -9106 2906
rect -9140 2777 -9106 2789
rect -9140 2705 -9106 2721
rect -9140 2633 -9106 2653
rect -9140 2561 -9106 2585
rect -9140 2489 -9106 2517
rect -9140 2417 -9106 2449
rect -9140 2347 -9106 2381
rect -9140 2279 -9106 2311
rect -9140 2211 -9106 2239
rect -9140 2143 -9106 2167
rect -9140 2075 -9106 2095
rect -9140 2007 -9106 2023
rect -9140 1939 -9106 1951
rect -9140 1860 -9106 1879
rect -9044 2849 -9010 2868
rect -9044 2777 -9010 2789
rect -9044 2705 -9010 2721
rect -9044 2633 -9010 2653
rect -9044 2561 -9010 2585
rect -9044 2489 -9010 2517
rect -9044 2417 -9010 2449
rect -9044 2347 -9010 2381
rect -9044 2279 -9010 2311
rect -9044 2211 -9010 2239
rect -9044 2143 -9010 2167
rect -9044 2075 -9010 2095
rect -9044 2007 -9010 2023
rect -9044 1939 -9010 1951
rect -9044 1818 -9010 1879
rect -8948 2849 -8914 2906
rect -8948 2777 -8914 2789
rect -8948 2705 -8914 2721
rect -8948 2633 -8914 2653
rect -8948 2561 -8914 2585
rect -8948 2489 -8914 2517
rect -8948 2417 -8914 2449
rect -8948 2347 -8914 2381
rect -8948 2279 -8914 2311
rect -8948 2211 -8914 2239
rect -8948 2143 -8914 2167
rect -8948 2075 -8914 2095
rect -8948 2007 -8914 2023
rect -8948 1939 -8914 1951
rect -8948 1860 -8914 1879
rect -8852 2849 -8818 2868
rect -8852 2777 -8818 2789
rect -8852 2705 -8818 2721
rect -8852 2633 -8818 2653
rect -8852 2561 -8818 2585
rect -8852 2489 -8818 2517
rect -8852 2417 -8818 2449
rect -8852 2347 -8818 2381
rect -8852 2279 -8818 2311
rect -8852 2211 -8818 2239
rect -8852 2143 -8818 2167
rect -8852 2075 -8818 2095
rect -8852 2007 -8818 2023
rect -8852 1939 -8818 1951
rect -8852 1818 -8818 1879
rect -8756 2849 -8722 2906
rect -8756 2777 -8722 2789
rect -8756 2705 -8722 2721
rect -8756 2633 -8722 2653
rect -8756 2561 -8722 2585
rect -8756 2489 -8722 2517
rect -8756 2417 -8722 2449
rect -8756 2347 -8722 2381
rect -8756 2279 -8722 2311
rect -8756 2211 -8722 2239
rect -8756 2143 -8722 2167
rect -8756 2075 -8722 2095
rect -8756 2007 -8722 2023
rect -8756 1939 -8722 1951
rect -8756 1860 -8722 1879
rect -8660 2849 -8626 2868
rect -8660 2777 -8626 2789
rect -8660 2705 -8626 2721
rect -8660 2633 -8626 2653
rect -8660 2561 -8626 2585
rect -8660 2489 -8626 2517
rect -8660 2417 -8626 2449
rect -8660 2347 -8626 2381
rect -8660 2279 -8626 2311
rect -8660 2211 -8626 2239
rect -8660 2143 -8626 2167
rect -8660 2075 -8626 2095
rect -8660 2007 -8626 2023
rect -8660 1939 -8626 1951
rect -8660 1818 -8626 1879
rect -8564 2849 -8530 2906
rect -8564 2777 -8530 2789
rect -8564 2705 -8530 2721
rect -8564 2633 -8530 2653
rect -8564 2561 -8530 2585
rect -8564 2489 -8530 2517
rect -8564 2417 -8530 2449
rect -8564 2347 -8530 2381
rect -8564 2279 -8530 2311
rect -8564 2211 -8530 2239
rect -8564 2143 -8530 2167
rect -8564 2075 -8530 2095
rect -8564 2007 -8530 2023
rect -8564 1939 -8530 1951
rect -8564 1860 -8530 1879
rect -8468 2849 -8434 2868
rect -8468 2777 -8434 2789
rect -8468 2705 -8434 2721
rect -8468 2633 -8434 2653
rect -8468 2561 -8434 2585
rect -8468 2489 -8434 2517
rect -8468 2417 -8434 2449
rect -8468 2347 -8434 2381
rect -8468 2279 -8434 2311
rect -8468 2211 -8434 2239
rect -8468 2143 -8434 2167
rect -8468 2075 -8434 2095
rect -8468 2007 -8434 2023
rect -8468 1939 -8434 1951
rect -8468 1818 -8434 1879
rect -8372 2849 -8338 2906
rect -8048 2910 -6670 2944
rect -8372 2777 -8338 2789
rect -8372 2705 -8338 2721
rect -8372 2633 -8338 2653
rect -8372 2561 -8338 2585
rect -8372 2489 -8338 2517
rect -8372 2417 -8338 2449
rect -8372 2347 -8338 2381
rect -8372 2279 -8338 2311
rect -8372 2211 -8338 2239
rect -8372 2143 -8338 2167
rect -8372 2075 -8338 2095
rect -8372 2007 -8338 2023
rect -8372 1939 -8338 1951
rect -8372 1860 -8338 1879
rect -8276 2849 -8242 2868
rect -8276 2777 -8242 2789
rect -8276 2705 -8242 2721
rect -8276 2633 -8242 2653
rect -8276 2561 -8242 2585
rect -8276 2489 -8242 2517
rect -8276 2417 -8242 2449
rect -8276 2347 -8242 2381
rect -8276 2279 -8242 2311
rect -8276 2211 -8242 2239
rect -8276 2143 -8242 2167
rect -8276 2075 -8242 2095
rect -8276 2007 -8242 2023
rect -8276 1939 -8242 1951
rect -8276 1818 -8242 1879
rect -8048 2841 -8014 2910
rect -8048 2769 -8014 2781
rect -8048 2697 -8014 2713
rect -8048 2625 -8014 2645
rect -8048 2553 -8014 2577
rect -8048 2481 -8014 2509
rect -8048 2409 -8014 2441
rect -8048 2339 -8014 2373
rect -8048 2271 -8014 2303
rect -8048 2203 -8014 2231
rect -8048 2135 -8014 2159
rect -8048 2067 -8014 2087
rect -8048 1999 -8014 2015
rect -8048 1931 -8014 1943
rect -8048 1852 -8014 1871
rect -7952 2841 -7918 2860
rect -7952 2769 -7918 2781
rect -7952 2697 -7918 2713
rect -7952 2625 -7918 2645
rect -7952 2553 -7918 2577
rect -7952 2481 -7918 2509
rect -7952 2409 -7918 2441
rect -7952 2339 -7918 2373
rect -7952 2271 -7918 2303
rect -7952 2203 -7918 2231
rect -7952 2135 -7918 2159
rect -7952 2067 -7918 2087
rect -7952 1999 -7918 2015
rect -7952 1931 -7918 1943
rect -10196 1802 -8242 1818
rect -7952 1810 -7918 1871
rect -7856 2841 -7822 2910
rect -7856 2769 -7822 2781
rect -7856 2697 -7822 2713
rect -7856 2625 -7822 2645
rect -7856 2553 -7822 2577
rect -7856 2481 -7822 2509
rect -7856 2409 -7822 2441
rect -7856 2339 -7822 2373
rect -7856 2271 -7822 2303
rect -7856 2203 -7822 2231
rect -7856 2135 -7822 2159
rect -7856 2067 -7822 2087
rect -7856 1999 -7822 2015
rect -7856 1931 -7822 1943
rect -7856 1852 -7822 1871
rect -7760 2841 -7726 2860
rect -7760 2769 -7726 2781
rect -7760 2697 -7726 2713
rect -7760 2625 -7726 2645
rect -7760 2553 -7726 2577
rect -7760 2481 -7726 2509
rect -7760 2409 -7726 2441
rect -7760 2339 -7726 2373
rect -7760 2271 -7726 2303
rect -7760 2203 -7726 2231
rect -7760 2135 -7726 2159
rect -7760 2067 -7726 2087
rect -7760 1999 -7726 2015
rect -7760 1931 -7726 1943
rect -7760 1810 -7726 1871
rect -7664 2841 -7630 2910
rect -7664 2769 -7630 2781
rect -7664 2697 -7630 2713
rect -7664 2625 -7630 2645
rect -7664 2553 -7630 2577
rect -7664 2481 -7630 2509
rect -7664 2409 -7630 2441
rect -7664 2339 -7630 2373
rect -7664 2271 -7630 2303
rect -7664 2203 -7630 2231
rect -7664 2135 -7630 2159
rect -7664 2067 -7630 2087
rect -7664 1999 -7630 2015
rect -7664 1931 -7630 1943
rect -7664 1852 -7630 1871
rect -7568 2841 -7534 2860
rect -7568 2769 -7534 2781
rect -7568 2697 -7534 2713
rect -7568 2625 -7534 2645
rect -7568 2553 -7534 2577
rect -7568 2481 -7534 2509
rect -7568 2409 -7534 2441
rect -7568 2339 -7534 2373
rect -7568 2271 -7534 2303
rect -7568 2203 -7534 2231
rect -7568 2135 -7534 2159
rect -7568 2067 -7534 2087
rect -7568 1999 -7534 2015
rect -7568 1931 -7534 1943
rect -7568 1810 -7534 1871
rect -7472 2841 -7438 2910
rect -7472 2769 -7438 2781
rect -7472 2697 -7438 2713
rect -7472 2625 -7438 2645
rect -7472 2553 -7438 2577
rect -7472 2481 -7438 2509
rect -7472 2409 -7438 2441
rect -7472 2339 -7438 2373
rect -7472 2271 -7438 2303
rect -7472 2203 -7438 2231
rect -7472 2135 -7438 2159
rect -7472 2067 -7438 2087
rect -7472 1999 -7438 2015
rect -7472 1931 -7438 1943
rect -7472 1852 -7438 1871
rect -7376 2841 -7342 2860
rect -7376 2769 -7342 2781
rect -7376 2697 -7342 2713
rect -7376 2625 -7342 2645
rect -7376 2553 -7342 2577
rect -7376 2481 -7342 2509
rect -7376 2409 -7342 2441
rect -7376 2339 -7342 2373
rect -7376 2271 -7342 2303
rect -7376 2203 -7342 2231
rect -7376 2135 -7342 2159
rect -7376 2067 -7342 2087
rect -7376 1999 -7342 2015
rect -7376 1931 -7342 1943
rect -7376 1810 -7342 1871
rect -7280 2841 -7246 2910
rect -7280 2769 -7246 2781
rect -7280 2697 -7246 2713
rect -7280 2625 -7246 2645
rect -7280 2553 -7246 2577
rect -7280 2481 -7246 2509
rect -7280 2409 -7246 2441
rect -7280 2339 -7246 2373
rect -7280 2271 -7246 2303
rect -7280 2203 -7246 2231
rect -7280 2135 -7246 2159
rect -7280 2067 -7246 2087
rect -7280 1999 -7246 2015
rect -7280 1931 -7246 1943
rect -7280 1852 -7246 1871
rect -7184 2841 -7150 2860
rect -7184 2769 -7150 2781
rect -7184 2697 -7150 2713
rect -7184 2625 -7150 2645
rect -7184 2553 -7150 2577
rect -7184 2481 -7150 2509
rect -7184 2409 -7150 2441
rect -7184 2339 -7150 2373
rect -7184 2271 -7150 2303
rect -7184 2203 -7150 2231
rect -7184 2135 -7150 2159
rect -7184 2067 -7150 2087
rect -7184 1999 -7150 2015
rect -7184 1931 -7150 1943
rect -7184 1810 -7150 1871
rect -7088 2841 -7054 2910
rect -7088 2769 -7054 2781
rect -7088 2697 -7054 2713
rect -7088 2625 -7054 2645
rect -7088 2553 -7054 2577
rect -7088 2481 -7054 2509
rect -7088 2409 -7054 2441
rect -7088 2339 -7054 2373
rect -7088 2271 -7054 2303
rect -7088 2203 -7054 2231
rect -7088 2135 -7054 2159
rect -7088 2067 -7054 2087
rect -7088 1999 -7054 2015
rect -7088 1931 -7054 1943
rect -7088 1852 -7054 1871
rect -6992 2841 -6958 2860
rect -6992 2769 -6958 2781
rect -6992 2697 -6958 2713
rect -6992 2625 -6958 2645
rect -6992 2553 -6958 2577
rect -6992 2481 -6958 2509
rect -6992 2409 -6958 2441
rect -6992 2339 -6958 2373
rect -6992 2271 -6958 2303
rect -6992 2203 -6958 2231
rect -6992 2135 -6958 2159
rect -6992 2067 -6958 2087
rect -6992 1999 -6958 2015
rect -6992 1931 -6958 1943
rect -6992 1810 -6958 1871
rect -6896 2841 -6862 2910
rect -6896 2769 -6862 2781
rect -6896 2697 -6862 2713
rect -6896 2625 -6862 2645
rect -6896 2553 -6862 2577
rect -6896 2481 -6862 2509
rect -6896 2409 -6862 2441
rect -6896 2339 -6862 2373
rect -6896 2271 -6862 2303
rect -6896 2203 -6862 2231
rect -6896 2135 -6862 2159
rect -6896 2067 -6862 2087
rect -6896 1999 -6862 2015
rect -6896 1931 -6862 1943
rect -6896 1852 -6862 1871
rect -6800 2841 -6766 2860
rect -6800 2769 -6766 2781
rect -6800 2697 -6766 2713
rect -6800 2625 -6766 2645
rect -6800 2553 -6766 2577
rect -6800 2481 -6766 2509
rect -6800 2409 -6766 2441
rect -6800 2339 -6766 2373
rect -6800 2271 -6766 2303
rect -6800 2203 -6766 2231
rect -6800 2135 -6766 2159
rect -6800 2067 -6766 2087
rect -6800 1999 -6766 2015
rect -6800 1931 -6766 1943
rect -6800 1810 -6766 1871
rect -6704 2841 -6670 2910
rect -6274 2918 -5472 2952
rect -5006 2942 -4972 3123
rect -1686 3221 -1652 3240
rect -1686 3149 -1652 3161
rect -1686 3077 -1652 3093
rect -4878 3008 -4862 3042
rect -4828 3008 -4812 3042
rect -1686 3005 -1652 3025
rect -6704 2769 -6670 2781
rect -6704 2697 -6670 2713
rect -6704 2625 -6670 2645
rect -6704 2553 -6670 2577
rect -6704 2481 -6670 2509
rect -6704 2409 -6670 2441
rect -6704 2339 -6670 2373
rect -6704 2271 -6670 2303
rect -6704 2203 -6670 2231
rect -6704 2135 -6670 2159
rect -6704 2067 -6670 2087
rect -6704 1999 -6670 2015
rect -6704 1931 -6670 1943
rect -6704 1852 -6670 1871
rect -6608 2841 -6574 2860
rect -6608 2769 -6574 2781
rect -6608 2697 -6574 2713
rect -6608 2625 -6574 2645
rect -6608 2553 -6574 2577
rect -6608 2481 -6574 2509
rect -6608 2409 -6574 2441
rect -6608 2339 -6574 2373
rect -6608 2271 -6574 2303
rect -6608 2203 -6574 2231
rect -6608 2135 -6574 2159
rect -6608 2067 -6574 2087
rect -6608 1999 -6574 2015
rect -6608 1931 -6574 1943
rect -6608 1810 -6574 1871
rect -7964 1802 -6574 1810
rect -6370 2845 -6336 2864
rect -6370 2773 -6336 2785
rect -6370 2701 -6336 2717
rect -6370 2629 -6336 2649
rect -6370 2557 -6336 2581
rect -6370 2485 -6336 2513
rect -6370 2413 -6336 2445
rect -6370 2343 -6336 2377
rect -6370 2275 -6336 2307
rect -6370 2207 -6336 2235
rect -6370 2139 -6336 2163
rect -6370 2071 -6336 2091
rect -6370 2003 -6336 2019
rect -6370 1935 -6336 1947
rect -6370 1822 -6336 1875
rect -6274 2845 -6240 2918
rect -6274 2773 -6240 2785
rect -6274 2701 -6240 2717
rect -6274 2629 -6240 2649
rect -6274 2557 -6240 2581
rect -6274 2485 -6240 2513
rect -6274 2413 -6240 2445
rect -6274 2343 -6240 2377
rect -6274 2275 -6240 2307
rect -6274 2207 -6240 2235
rect -6274 2139 -6240 2163
rect -6274 2071 -6240 2091
rect -6274 2003 -6240 2019
rect -6274 1935 -6240 1947
rect -6274 1856 -6240 1875
rect -6178 2845 -6144 2864
rect -6178 2773 -6144 2785
rect -6178 2701 -6144 2717
rect -6178 2629 -6144 2649
rect -6178 2557 -6144 2581
rect -6178 2485 -6144 2513
rect -6178 2413 -6144 2445
rect -6178 2343 -6144 2377
rect -6178 2275 -6144 2307
rect -6178 2207 -6144 2235
rect -6178 2139 -6144 2163
rect -6178 2071 -6144 2091
rect -6178 2003 -6144 2019
rect -6178 1935 -6144 1947
rect -6178 1822 -6144 1875
rect -6082 2845 -6048 2918
rect -6082 2773 -6048 2785
rect -6082 2701 -6048 2717
rect -6082 2629 -6048 2649
rect -6082 2557 -6048 2581
rect -6082 2485 -6048 2513
rect -6082 2413 -6048 2445
rect -6082 2343 -6048 2377
rect -6082 2275 -6048 2307
rect -6082 2207 -6048 2235
rect -6082 2139 -6048 2163
rect -6082 2071 -6048 2091
rect -6082 2003 -6048 2019
rect -6082 1935 -6048 1947
rect -6082 1856 -6048 1875
rect -5986 2845 -5952 2864
rect -5986 2773 -5952 2785
rect -5986 2701 -5952 2717
rect -5986 2629 -5952 2649
rect -5986 2557 -5952 2581
rect -5986 2485 -5952 2513
rect -5986 2413 -5952 2445
rect -5986 2343 -5952 2377
rect -5986 2275 -5952 2307
rect -5986 2207 -5952 2235
rect -5986 2139 -5952 2163
rect -5986 2071 -5952 2091
rect -5986 2003 -5952 2019
rect -5986 1935 -5952 1947
rect -5986 1822 -5952 1875
rect -5890 2845 -5856 2918
rect -5890 2773 -5856 2785
rect -5890 2701 -5856 2717
rect -5890 2629 -5856 2649
rect -5890 2557 -5856 2581
rect -5890 2485 -5856 2513
rect -5890 2413 -5856 2445
rect -5890 2343 -5856 2377
rect -5890 2275 -5856 2307
rect -5890 2207 -5856 2235
rect -5890 2139 -5856 2163
rect -5890 2071 -5856 2091
rect -5890 2003 -5856 2019
rect -5890 1935 -5856 1947
rect -5890 1856 -5856 1875
rect -5794 2845 -5760 2864
rect -5794 2773 -5760 2785
rect -5794 2701 -5760 2717
rect -5794 2629 -5760 2649
rect -5794 2557 -5760 2581
rect -5794 2485 -5760 2513
rect -5794 2413 -5760 2445
rect -5794 2343 -5760 2377
rect -5794 2275 -5760 2307
rect -5794 2207 -5760 2235
rect -5794 2139 -5760 2163
rect -5794 2071 -5760 2091
rect -5794 2003 -5760 2019
rect -5794 1935 -5760 1947
rect -5794 1822 -5760 1875
rect -5698 2845 -5664 2918
rect -5698 2773 -5664 2785
rect -5698 2701 -5664 2717
rect -5698 2629 -5664 2649
rect -5698 2557 -5664 2581
rect -5698 2485 -5664 2513
rect -5698 2413 -5664 2445
rect -5698 2343 -5664 2377
rect -5698 2275 -5664 2307
rect -5698 2207 -5664 2235
rect -5698 2139 -5664 2163
rect -5698 2071 -5664 2091
rect -5698 2003 -5664 2019
rect -5698 1935 -5664 1947
rect -5698 1856 -5664 1875
rect -5602 2845 -5568 2864
rect -5602 2773 -5568 2785
rect -5602 2701 -5568 2717
rect -5602 2629 -5568 2649
rect -5602 2557 -5568 2581
rect -5602 2485 -5568 2513
rect -5602 2413 -5568 2445
rect -5602 2343 -5568 2377
rect -5602 2275 -5568 2307
rect -5602 2207 -5568 2235
rect -5602 2139 -5568 2163
rect -5602 2071 -5568 2091
rect -5602 2003 -5568 2019
rect -5602 1935 -5568 1947
rect -5602 1822 -5568 1875
rect -5506 2845 -5472 2918
rect -5198 2908 -4780 2942
rect -5506 2773 -5472 2785
rect -5506 2701 -5472 2717
rect -5506 2629 -5472 2649
rect -5506 2557 -5472 2581
rect -5506 2485 -5472 2513
rect -5506 2413 -5472 2445
rect -5506 2343 -5472 2377
rect -5506 2275 -5472 2307
rect -5506 2207 -5472 2235
rect -5506 2139 -5472 2163
rect -5506 2071 -5472 2091
rect -5506 2003 -5472 2019
rect -5506 1935 -5472 1947
rect -5506 1856 -5472 1875
rect -5410 2845 -5376 2864
rect -5410 2773 -5376 2785
rect -5410 2701 -5376 2717
rect -5410 2629 -5376 2649
rect -5410 2557 -5376 2581
rect -5410 2485 -5376 2513
rect -5410 2413 -5376 2445
rect -5410 2343 -5376 2377
rect -5410 2275 -5376 2307
rect -5410 2207 -5376 2235
rect -5410 2139 -5376 2163
rect -5410 2071 -5376 2091
rect -5410 2003 -5376 2019
rect -5410 1935 -5376 1947
rect -5410 1822 -5376 1875
rect -5198 2855 -5164 2908
rect -5198 2783 -5164 2795
rect -5198 2711 -5164 2727
rect -5198 2639 -5164 2659
rect -5198 2567 -5164 2591
rect -5198 2495 -5164 2523
rect -5198 2423 -5164 2455
rect -5198 2353 -5164 2387
rect -5198 2285 -5164 2317
rect -5198 2217 -5164 2245
rect -5198 2149 -5164 2173
rect -5198 2081 -5164 2101
rect -5198 2013 -5164 2029
rect -5198 1945 -5164 1957
rect -5198 1866 -5164 1885
rect -5102 2855 -5068 2874
rect -5102 2783 -5068 2795
rect -5102 2711 -5068 2727
rect -5102 2639 -5068 2659
rect -5102 2567 -5068 2591
rect -5102 2495 -5068 2523
rect -5102 2423 -5068 2455
rect -5102 2353 -5068 2387
rect -5102 2285 -5068 2317
rect -5102 2217 -5068 2245
rect -5102 2149 -5068 2173
rect -5102 2081 -5068 2101
rect -5102 2013 -5068 2029
rect -5102 1945 -5068 1957
rect -6370 1802 -5376 1822
rect -5102 1818 -5068 1885
rect -5006 2855 -4972 2908
rect -5006 2783 -4972 2795
rect -5006 2711 -4972 2727
rect -5006 2639 -4972 2659
rect -5006 2567 -4972 2591
rect -5006 2495 -4972 2523
rect -5006 2423 -4972 2455
rect -5006 2353 -4972 2387
rect -5006 2285 -4972 2317
rect -5006 2217 -4972 2245
rect -5006 2149 -4972 2173
rect -5006 2081 -4972 2101
rect -5006 2013 -4972 2029
rect -5006 1945 -4972 1957
rect -5006 1866 -4972 1885
rect -4910 2855 -4876 2874
rect -4910 2783 -4876 2795
rect -4910 2711 -4876 2727
rect -4910 2639 -4876 2659
rect -4910 2567 -4876 2591
rect -4910 2495 -4876 2523
rect -4910 2423 -4876 2455
rect -4910 2353 -4876 2387
rect -4910 2285 -4876 2317
rect -4910 2217 -4876 2245
rect -4910 2149 -4876 2173
rect -4910 2081 -4876 2101
rect -4910 2013 -4876 2029
rect -4910 1945 -4876 1957
rect -4910 1818 -4876 1885
rect -4814 2855 -4780 2908
rect -1686 2933 -1652 2957
rect -4814 2783 -4780 2795
rect -4814 2711 -4780 2727
rect -4814 2639 -4780 2659
rect -4814 2567 -4780 2591
rect -4814 2495 -4780 2523
rect -4814 2423 -4780 2455
rect -4814 2353 -4780 2387
rect -4814 2285 -4780 2317
rect -4814 2217 -4780 2245
rect -4814 2149 -4780 2173
rect -4814 2081 -4780 2101
rect -4814 2013 -4780 2029
rect -4814 1945 -4780 1957
rect -4814 1866 -4780 1885
rect -4718 2855 -4684 2874
rect -4718 2783 -4684 2795
rect -4718 2711 -4684 2727
rect -4718 2639 -4684 2659
rect -4718 2567 -4684 2591
rect -4718 2495 -4684 2523
rect -4718 2423 -4684 2455
rect -4718 2353 -4684 2387
rect -4718 2285 -4684 2317
rect -4718 2217 -4684 2245
rect -4718 2149 -4684 2173
rect -1686 2861 -1652 2889
rect -1686 2789 -1652 2821
rect -1686 2719 -1652 2753
rect -1686 2651 -1652 2683
rect -1686 2583 -1652 2611
rect -1686 2515 -1652 2539
rect -1686 2447 -1652 2467
rect -1686 2379 -1652 2395
rect -1686 2311 -1652 2323
rect -1686 2172 -1652 2251
rect -1590 3221 -1556 3290
rect -1590 3149 -1556 3161
rect -1590 3077 -1556 3093
rect -1590 3005 -1556 3025
rect -1590 2933 -1556 2957
rect -1590 2861 -1556 2889
rect -1590 2789 -1556 2821
rect -1590 2719 -1556 2753
rect -1590 2651 -1556 2683
rect -1590 2583 -1556 2611
rect -1590 2515 -1556 2539
rect -1590 2447 -1556 2467
rect -1590 2379 -1556 2395
rect -1590 2311 -1556 2323
rect -1590 2232 -1556 2251
rect -1494 3221 -1460 3240
rect -1494 3149 -1460 3161
rect -1494 3077 -1460 3093
rect -1494 3005 -1460 3025
rect -1494 2933 -1460 2957
rect -1494 2861 -1460 2889
rect -1494 2789 -1460 2821
rect -1494 2719 -1460 2753
rect -1494 2651 -1460 2683
rect -1494 2583 -1460 2611
rect -1494 2515 -1460 2539
rect -1494 2447 -1460 2467
rect -1494 2379 -1460 2395
rect -1494 2311 -1460 2323
rect -1494 2172 -1460 2251
rect -1398 3221 -1364 3290
rect -1398 3149 -1364 3161
rect -1398 3077 -1364 3093
rect -1398 3005 -1364 3025
rect -1398 2933 -1364 2957
rect -1398 2861 -1364 2889
rect -1398 2789 -1364 2821
rect -1398 2719 -1364 2753
rect -1398 2651 -1364 2683
rect -1398 2583 -1364 2611
rect -1398 2515 -1364 2539
rect -1398 2447 -1364 2467
rect -1398 2379 -1364 2395
rect -1398 2311 -1364 2323
rect -1398 2232 -1364 2251
rect -1302 3221 -1268 3240
rect -1302 3149 -1268 3161
rect -1302 3077 -1268 3093
rect -1302 3005 -1268 3025
rect -1302 2933 -1268 2957
rect -1302 2861 -1268 2889
rect -1302 2789 -1268 2821
rect -1302 2719 -1268 2753
rect -1302 2651 -1268 2683
rect -1302 2583 -1268 2611
rect -1302 2515 -1268 2539
rect -1302 2447 -1268 2467
rect -1302 2379 -1268 2395
rect -1302 2311 -1268 2323
rect -1302 2172 -1268 2251
rect -1206 3221 -1172 3290
rect -1206 3149 -1172 3161
rect -1206 3077 -1172 3093
rect -1206 3005 -1172 3025
rect -1206 2933 -1172 2957
rect -1206 2861 -1172 2889
rect -1206 2789 -1172 2821
rect -1206 2719 -1172 2753
rect -1206 2651 -1172 2683
rect -1206 2583 -1172 2611
rect -1206 2515 -1172 2539
rect -1206 2447 -1172 2467
rect -1206 2379 -1172 2395
rect -1206 2311 -1172 2323
rect -1206 2232 -1172 2251
rect -1110 3221 -1076 3240
rect -1110 3149 -1076 3161
rect -1110 3077 -1076 3093
rect -1110 3005 -1076 3025
rect -1110 2933 -1076 2957
rect -1110 2861 -1076 2889
rect -1110 2789 -1076 2821
rect -1110 2719 -1076 2753
rect -1110 2651 -1076 2683
rect -1110 2583 -1076 2611
rect -1110 2515 -1076 2539
rect -1110 2447 -1076 2467
rect -1110 2379 -1076 2395
rect -1110 2311 -1076 2323
rect -1110 2172 -1076 2251
rect -1014 3221 -980 3290
rect 16686 3303 16720 3323
rect -1014 3149 -980 3161
rect -1014 3077 -980 3093
rect -1014 3005 -980 3025
rect -1014 2933 -980 2957
rect -1014 2861 -980 2889
rect -1014 2789 -980 2821
rect -1014 2719 -980 2753
rect -1014 2651 -980 2683
rect -1014 2583 -980 2611
rect -1014 2515 -980 2539
rect -1014 2447 -980 2467
rect -1014 2379 -980 2395
rect -1014 2311 -980 2323
rect -1014 2232 -980 2251
rect -918 3221 -884 3240
rect -918 3149 -884 3161
rect -918 3077 -884 3093
rect -918 3005 -884 3025
rect 16686 3231 16720 3255
rect 16686 3159 16720 3187
rect 16686 3087 16720 3119
rect 16686 3017 16720 3051
rect 1562 2968 1578 3002
rect 1612 2968 1628 3002
rect -918 2933 -884 2957
rect 1674 2906 1708 2960
rect 4518 2952 4534 2986
rect 4568 2952 4584 2986
rect 7548 2952 7564 2986
rect 7598 2952 7614 2986
rect -918 2861 -884 2889
rect 1578 2872 1804 2906
rect 4630 2890 4664 2944
rect 10636 2950 10652 2984
rect 10686 2950 10702 2984
rect 7660 2890 7694 2944
rect -918 2789 -884 2821
rect -918 2719 -884 2753
rect -918 2651 -884 2683
rect -918 2583 -884 2611
rect -918 2515 -884 2539
rect -918 2447 -884 2467
rect -918 2379 -884 2395
rect -918 2311 -884 2323
rect -918 2172 -884 2251
rect -1686 2138 -1097 2172
rect -1063 2138 -884 2172
rect 1482 2815 1516 2832
rect 1482 2743 1516 2755
rect 1482 2671 1516 2687
rect 1482 2599 1516 2619
rect 1482 2527 1516 2551
rect 1482 2455 1516 2483
rect 1482 2383 1516 2415
rect 1482 2313 1516 2347
rect 1482 2245 1516 2277
rect 1482 2177 1516 2205
rect -4718 2081 -4684 2101
rect -4718 2013 -4684 2029
rect -4718 1945 -4684 1957
rect -4718 1818 -4684 1885
rect -5102 1802 -4684 1818
rect -23492 1668 -18012 1774
rect -16662 1680 -11182 1786
rect -10196 1784 -4684 1802
rect 1482 2109 1516 2133
rect 1482 2041 1516 2061
rect 1482 1973 1516 1989
rect 1482 1905 1516 1917
rect -16732 1672 -11114 1680
rect -10196 1678 -4716 1784
rect 1482 1780 1516 1845
rect 1578 2815 1612 2872
rect 1674 2868 1708 2872
rect 1578 2743 1612 2755
rect 1578 2671 1612 2687
rect 1578 2599 1612 2619
rect 1578 2527 1612 2551
rect 1578 2455 1612 2483
rect 1578 2383 1612 2415
rect 1578 2313 1612 2347
rect 1578 2245 1612 2277
rect 1578 2177 1612 2205
rect 1578 2109 1612 2133
rect 1578 2041 1612 2061
rect 1578 1973 1612 1989
rect 1578 1905 1612 1917
rect 1578 1826 1612 1845
rect 1674 2815 1708 2832
rect 1674 2743 1708 2755
rect 1674 2671 1708 2687
rect 1674 2599 1708 2619
rect 1674 2527 1708 2551
rect 1674 2455 1708 2483
rect 1674 2383 1708 2415
rect 1674 2313 1708 2347
rect 1674 2245 1708 2277
rect 1674 2177 1708 2205
rect 1674 2109 1708 2133
rect 1674 2041 1708 2061
rect 1674 1973 1708 1989
rect 1674 1905 1708 1917
rect 1674 1780 1708 1845
rect 1770 2815 1804 2872
rect 4534 2856 4760 2890
rect 1770 2743 1804 2755
rect 1770 2671 1804 2687
rect 1770 2599 1804 2619
rect 1770 2527 1804 2551
rect 1770 2455 1804 2483
rect 1770 2383 1804 2415
rect 1770 2313 1804 2347
rect 1770 2245 1804 2277
rect 1770 2177 1804 2205
rect 1770 2109 1804 2133
rect 1770 2041 1804 2061
rect 1770 1973 1804 1989
rect 1770 1905 1804 1917
rect 1770 1828 1804 1845
rect 1866 2815 1900 2832
rect 1866 2743 1900 2755
rect 1866 2671 1900 2687
rect 1866 2599 1900 2619
rect 1866 2527 1900 2551
rect 1866 2455 1900 2483
rect 4438 2799 4472 2816
rect 4438 2727 4472 2739
rect 4438 2655 4472 2671
rect 4438 2583 4472 2603
rect 4438 2511 4472 2535
rect 4438 2439 4472 2467
rect 1866 2383 1900 2415
rect 2546 2394 2579 2428
rect 2613 2394 2646 2428
rect 4438 2367 4472 2399
rect 1866 2313 1900 2347
rect 2426 2316 2692 2350
rect 1866 2245 1900 2277
rect 1866 2177 1900 2205
rect 1866 2109 1900 2133
rect 1866 2041 1900 2061
rect 1866 1973 1900 1989
rect 1866 1905 1900 1917
rect 2500 2261 2534 2280
rect 2500 2193 2534 2195
rect 2500 2157 2534 2159
rect 2500 1912 2534 2091
rect 2658 2261 2692 2316
rect 2658 2193 2692 2195
rect 2658 2157 2692 2159
rect 2658 2072 2692 2091
rect 4438 2297 4472 2331
rect 4438 2229 4472 2261
rect 4438 2161 4472 2189
rect 4438 2093 4472 2117
rect 1866 1780 1900 1845
rect 1482 1746 1900 1780
rect 2102 1878 2534 1912
rect 4438 2025 4472 2045
rect 4438 1957 4472 1973
rect 4438 1889 4472 1901
rect 1578 1696 1612 1746
rect -23562 1660 -17944 1668
rect -23562 1490 -23524 1660
rect -17982 1490 -17944 1660
rect -16732 1502 -16694 1672
rect -11152 1502 -11114 1672
rect -16732 1494 -11114 1502
rect -10266 1670 -4648 1678
rect -10266 1500 -10228 1670
rect -4686 1500 -4648 1670
rect 2102 1522 2136 1878
rect 4438 1764 4472 1829
rect 4534 2799 4568 2856
rect 4630 2852 4664 2856
rect 4534 2727 4568 2739
rect 4534 2655 4568 2671
rect 4534 2583 4568 2603
rect 4534 2511 4568 2535
rect 4534 2439 4568 2467
rect 4534 2367 4568 2399
rect 4534 2297 4568 2331
rect 4534 2229 4568 2261
rect 4534 2161 4568 2189
rect 4534 2093 4568 2117
rect 4534 2025 4568 2045
rect 4534 1957 4568 1973
rect 4534 1889 4568 1901
rect 4534 1810 4568 1829
rect 4630 2799 4664 2816
rect 4630 2727 4664 2739
rect 4630 2655 4664 2671
rect 4630 2583 4664 2603
rect 4630 2511 4664 2535
rect 4630 2439 4664 2467
rect 4630 2367 4664 2399
rect 4630 2297 4664 2331
rect 4630 2229 4664 2261
rect 4630 2161 4664 2189
rect 4630 2093 4664 2117
rect 4630 2025 4664 2045
rect 4630 1957 4664 1973
rect 4630 1889 4664 1901
rect 4630 1764 4664 1829
rect 4726 2799 4760 2856
rect 7564 2856 7790 2890
rect 10748 2888 10782 2942
rect 13792 2924 13808 2958
rect 13842 2924 13858 2958
rect 4726 2727 4760 2739
rect 4726 2655 4760 2671
rect 4726 2583 4760 2603
rect 4726 2511 4760 2535
rect 4726 2439 4760 2467
rect 4726 2367 4760 2399
rect 4726 2297 4760 2331
rect 4726 2229 4760 2261
rect 4726 2161 4760 2189
rect 4726 2093 4760 2117
rect 4726 2025 4760 2045
rect 4726 1957 4760 1973
rect 4726 1889 4760 1901
rect 4726 1812 4760 1829
rect 4822 2799 4856 2816
rect 4822 2727 4856 2739
rect 4822 2655 4856 2671
rect 4822 2583 4856 2603
rect 4822 2511 4856 2535
rect 4822 2439 4856 2467
rect 7468 2799 7502 2816
rect 7468 2727 7502 2739
rect 7468 2655 7502 2671
rect 7468 2583 7502 2603
rect 7468 2511 7502 2535
rect 7468 2439 7502 2467
rect 4822 2367 4856 2399
rect 5546 2394 5579 2428
rect 5613 2394 5646 2428
rect 7468 2367 7502 2399
rect 4822 2297 4856 2331
rect 5426 2316 5692 2350
rect 4822 2229 4856 2261
rect 4822 2161 4856 2189
rect 4822 2093 4856 2117
rect 4822 2025 4856 2045
rect 4822 1957 4856 1973
rect 4822 1889 4856 1901
rect 4822 1764 4856 1829
rect 5500 2261 5534 2280
rect 5500 2193 5534 2195
rect 5500 2157 5534 2159
rect 5500 1788 5534 2091
rect 5658 2261 5692 2316
rect 5658 2193 5692 2195
rect 5658 2157 5692 2159
rect 5658 2070 5692 2091
rect 7468 2297 7502 2331
rect 7468 2229 7502 2261
rect 7468 2161 7502 2189
rect 7468 2093 7502 2117
rect 4438 1730 4856 1764
rect 4974 1754 5534 1788
rect 7468 2025 7502 2045
rect 7468 1957 7502 1973
rect 7468 1889 7502 1901
rect 7468 1764 7502 1829
rect 7564 2799 7598 2856
rect 7660 2852 7694 2856
rect 7564 2727 7598 2739
rect 7564 2655 7598 2671
rect 7564 2583 7598 2603
rect 7564 2511 7598 2535
rect 7564 2439 7598 2467
rect 7564 2367 7598 2399
rect 7564 2297 7598 2331
rect 7564 2229 7598 2261
rect 7564 2161 7598 2189
rect 7564 2093 7598 2117
rect 7564 2025 7598 2045
rect 7564 1957 7598 1973
rect 7564 1889 7598 1901
rect 7564 1810 7598 1829
rect 7660 2799 7694 2816
rect 7660 2727 7694 2739
rect 7660 2655 7694 2671
rect 7660 2583 7694 2603
rect 7660 2511 7694 2535
rect 7660 2439 7694 2467
rect 7660 2367 7694 2399
rect 7660 2297 7694 2331
rect 7660 2229 7694 2261
rect 7660 2161 7694 2189
rect 7660 2093 7694 2117
rect 7660 2025 7694 2045
rect 7660 1957 7694 1973
rect 7660 1889 7694 1901
rect 7660 1764 7694 1829
rect 7756 2799 7790 2856
rect 10652 2854 10878 2888
rect 13904 2862 13938 2916
rect 16686 2949 16720 2981
rect 16686 2881 16720 2909
rect 7756 2727 7790 2739
rect 7756 2655 7790 2671
rect 7756 2583 7790 2603
rect 7756 2511 7790 2535
rect 7756 2439 7790 2467
rect 7756 2367 7790 2399
rect 7756 2297 7790 2331
rect 7756 2229 7790 2261
rect 7756 2161 7790 2189
rect 7756 2093 7790 2117
rect 7756 2025 7790 2045
rect 7756 1957 7790 1973
rect 7756 1889 7790 1901
rect 7756 1812 7790 1829
rect 7852 2799 7886 2816
rect 7852 2727 7886 2739
rect 7852 2655 7886 2671
rect 7852 2583 7886 2603
rect 7852 2511 7886 2535
rect 7852 2439 7886 2467
rect 10556 2797 10590 2814
rect 10556 2725 10590 2737
rect 10556 2653 10590 2669
rect 10556 2581 10590 2601
rect 10556 2509 10590 2533
rect 10556 2437 10590 2465
rect 7852 2367 7886 2399
rect 8546 2394 8579 2428
rect 8613 2394 8646 2428
rect 10556 2365 10590 2397
rect 7852 2297 7886 2331
rect 8426 2316 8692 2350
rect 7852 2229 7886 2261
rect 7852 2161 7886 2189
rect 7852 2093 7886 2117
rect 7852 2025 7886 2045
rect 7852 1957 7886 1973
rect 7852 1889 7886 1901
rect 7852 1764 7886 1829
rect 8500 2261 8534 2280
rect 8500 2193 8534 2195
rect 8500 2157 8534 2159
rect 8500 1802 8534 2091
rect 8658 2261 8692 2316
rect 8658 2193 8692 2195
rect 8658 2157 8692 2159
rect 8658 2070 8692 2091
rect 10556 2295 10590 2329
rect 10556 2227 10590 2259
rect 10556 2159 10590 2187
rect 10556 2091 10590 2115
rect 4534 1680 4568 1730
rect -10266 1492 -4648 1500
rect -23562 1482 -17944 1490
rect 1484 1488 2136 1522
rect 4974 1490 5008 1754
rect 7468 1730 7886 1764
rect 8002 1768 8534 1802
rect 10556 2023 10590 2043
rect 10556 1955 10590 1971
rect 10556 1887 10590 1899
rect 7564 1680 7598 1730
rect 8002 1496 8036 1768
rect 10556 1762 10590 1827
rect 10652 2797 10686 2854
rect 10748 2850 10782 2854
rect 10652 2725 10686 2737
rect 10652 2653 10686 2669
rect 10652 2581 10686 2601
rect 10652 2509 10686 2533
rect 10652 2437 10686 2465
rect 10652 2365 10686 2397
rect 10652 2295 10686 2329
rect 10652 2227 10686 2259
rect 10652 2159 10686 2187
rect 10652 2091 10686 2115
rect 10652 2023 10686 2043
rect 10652 1955 10686 1971
rect 10652 1887 10686 1899
rect 10652 1808 10686 1827
rect 10748 2797 10782 2814
rect 10748 2725 10782 2737
rect 10748 2653 10782 2669
rect 10748 2581 10782 2601
rect 10748 2509 10782 2533
rect 10748 2437 10782 2465
rect 10748 2365 10782 2397
rect 10748 2295 10782 2329
rect 10748 2227 10782 2259
rect 10748 2159 10782 2187
rect 10748 2091 10782 2115
rect 10748 2023 10782 2043
rect 10748 1955 10782 1971
rect 10748 1887 10782 1899
rect 10748 1762 10782 1827
rect 10844 2797 10878 2854
rect 13808 2828 14034 2862
rect 10844 2725 10878 2737
rect 10844 2653 10878 2669
rect 10844 2581 10878 2601
rect 10844 2509 10878 2533
rect 10844 2437 10878 2465
rect 10844 2365 10878 2397
rect 10844 2295 10878 2329
rect 10844 2227 10878 2259
rect 10844 2159 10878 2187
rect 10844 2091 10878 2115
rect 10844 2023 10878 2043
rect 10844 1955 10878 1971
rect 10844 1887 10878 1899
rect 10844 1810 10878 1827
rect 10940 2797 10974 2814
rect 10940 2725 10974 2737
rect 10940 2653 10974 2669
rect 10940 2581 10974 2601
rect 10940 2509 10974 2533
rect 10940 2437 10974 2465
rect 13712 2771 13746 2788
rect 13712 2699 13746 2711
rect 13712 2627 13746 2643
rect 13712 2555 13746 2575
rect 13712 2483 13746 2507
rect 10940 2365 10974 2397
rect 11546 2394 11579 2428
rect 11613 2394 11646 2428
rect 13712 2411 13746 2439
rect 10940 2295 10974 2329
rect 11426 2316 11692 2350
rect 10940 2227 10974 2259
rect 10940 2159 10974 2187
rect 10940 2091 10974 2115
rect 10940 2023 10974 2043
rect 10940 1955 10974 1971
rect 10940 1887 10974 1899
rect 10940 1762 10974 1827
rect 10556 1728 10974 1762
rect 11500 2261 11534 2280
rect 11500 2193 11534 2195
rect 11500 2157 11534 2159
rect 10652 1678 10686 1728
rect 11500 1690 11534 2091
rect 11658 2261 11692 2316
rect 11658 2193 11692 2195
rect 11658 2157 11692 2159
rect 11658 2068 11692 2091
rect 13712 2339 13746 2371
rect 13712 2269 13746 2303
rect 13712 2201 13746 2233
rect 13712 2133 13746 2161
rect 13712 2065 13746 2089
rect 13712 1997 13746 2017
rect 13712 1929 13746 1945
rect 13712 1861 13746 1873
rect 13712 1736 13746 1801
rect 13808 2771 13842 2828
rect 13904 2824 13938 2828
rect 13808 2699 13842 2711
rect 13808 2627 13842 2643
rect 13808 2555 13842 2575
rect 13808 2483 13842 2507
rect 13808 2411 13842 2439
rect 13808 2339 13842 2371
rect 13808 2269 13842 2303
rect 13808 2201 13842 2233
rect 13808 2133 13842 2161
rect 13808 2065 13842 2089
rect 13808 1997 13842 2017
rect 13808 1929 13842 1945
rect 13808 1861 13842 1873
rect 13808 1782 13842 1801
rect 13904 2771 13938 2788
rect 13904 2699 13938 2711
rect 13904 2627 13938 2643
rect 13904 2555 13938 2575
rect 13904 2483 13938 2507
rect 13904 2411 13938 2439
rect 13904 2339 13938 2371
rect 13904 2269 13938 2303
rect 13904 2201 13938 2233
rect 13904 2133 13938 2161
rect 13904 2065 13938 2089
rect 13904 1997 13938 2017
rect 13904 1929 13938 1945
rect 13904 1861 13938 1873
rect 13904 1736 13938 1801
rect 14000 2771 14034 2828
rect 16686 2813 16720 2837
rect 14000 2699 14034 2711
rect 14000 2627 14034 2643
rect 14000 2555 14034 2575
rect 14000 2483 14034 2507
rect 14000 2411 14034 2439
rect 14000 2339 14034 2371
rect 14000 2269 14034 2303
rect 14000 2201 14034 2233
rect 14000 2133 14034 2161
rect 14000 2065 14034 2089
rect 14000 1997 14034 2017
rect 14000 1929 14034 1945
rect 14000 1861 14034 1873
rect 14000 1784 14034 1801
rect 14096 2771 14130 2788
rect 14096 2699 14130 2711
rect 14096 2627 14130 2643
rect 14096 2555 14130 2575
rect 14096 2483 14130 2507
rect 14096 2411 14130 2439
rect 16686 2745 16720 2765
rect 16686 2677 16720 2693
rect 16686 2609 16720 2621
rect 16686 2482 16720 2549
rect 16782 3519 16816 3572
rect 16782 3447 16816 3459
rect 16782 3375 16816 3391
rect 16782 3303 16816 3323
rect 16782 3231 16816 3255
rect 16782 3159 16816 3187
rect 16782 3087 16816 3119
rect 16782 3017 16816 3051
rect 16782 2949 16816 2981
rect 16782 2881 16816 2909
rect 16782 2813 16816 2837
rect 16782 2745 16816 2765
rect 16782 2677 16816 2693
rect 16782 2609 16816 2621
rect 16782 2530 16816 2549
rect 16878 3519 16912 3538
rect 16878 3447 16912 3459
rect 16878 3375 16912 3391
rect 16878 3303 16912 3323
rect 16878 3231 16912 3255
rect 16878 3159 16912 3187
rect 16878 3087 16912 3119
rect 16878 3017 16912 3051
rect 16878 2949 16912 2981
rect 16878 2881 16912 2909
rect 16878 2813 16912 2837
rect 16878 2745 16912 2765
rect 16878 2677 16912 2693
rect 16878 2609 16912 2621
rect 16878 2482 16912 2549
rect 16974 3519 17008 3572
rect 16974 3447 17008 3459
rect 16974 3375 17008 3391
rect 16974 3303 17008 3323
rect 16974 3231 17008 3255
rect 16974 3159 17008 3187
rect 16974 3087 17008 3119
rect 16974 3017 17008 3051
rect 16974 2949 17008 2981
rect 16974 2881 17008 2909
rect 16974 2813 17008 2837
rect 16974 2745 17008 2765
rect 16974 2677 17008 2693
rect 16974 2609 17008 2621
rect 16974 2530 17008 2549
rect 17070 3519 17104 3538
rect 17070 3447 17104 3459
rect 17070 3375 17104 3391
rect 17070 3303 17104 3323
rect 17070 3231 17104 3255
rect 17070 3159 17104 3187
rect 17070 3087 17104 3119
rect 17070 3017 17104 3051
rect 17070 2949 17104 2981
rect 17070 2881 17104 2909
rect 17070 2813 17104 2837
rect 17070 2745 17104 2765
rect 17070 2677 17104 2693
rect 17070 2609 17104 2621
rect 17070 2482 17104 2549
rect 17166 3519 17200 3572
rect 17474 3582 18276 3616
rect 19440 3608 19480 3772
rect 21640 3804 21686 4032
rect 23302 3907 23318 3941
rect 23352 3907 23368 3941
rect 21640 3770 21646 3804
rect 21680 3770 21686 3804
rect 20372 3656 20388 3690
rect 20422 3656 20438 3690
rect 17166 3447 17200 3459
rect 17166 3375 17200 3391
rect 17166 3303 17200 3323
rect 17166 3231 17200 3255
rect 17166 3159 17200 3187
rect 17166 3087 17200 3119
rect 17166 3017 17200 3051
rect 17166 2949 17200 2981
rect 17166 2881 17200 2909
rect 17166 2813 17200 2837
rect 17166 2745 17200 2765
rect 17166 2677 17200 2693
rect 17166 2609 17200 2621
rect 17166 2530 17200 2549
rect 17378 3509 17412 3528
rect 17378 3437 17412 3449
rect 17378 3365 17412 3381
rect 17378 3293 17412 3313
rect 17378 3221 17412 3245
rect 17378 3149 17412 3177
rect 17378 3077 17412 3109
rect 17378 3007 17412 3041
rect 17378 2939 17412 2971
rect 17378 2871 17412 2899
rect 17378 2803 17412 2827
rect 17378 2735 17412 2755
rect 17378 2667 17412 2683
rect 17378 2599 17412 2611
rect 16686 2460 17104 2482
rect 17378 2486 17412 2539
rect 17474 3509 17508 3582
rect 17474 3437 17508 3449
rect 17474 3365 17508 3381
rect 17474 3293 17508 3313
rect 17474 3221 17508 3245
rect 17474 3149 17508 3177
rect 17474 3077 17508 3109
rect 17474 3007 17508 3041
rect 17474 2939 17508 2971
rect 17474 2871 17508 2899
rect 17474 2803 17508 2827
rect 17474 2735 17508 2755
rect 17474 2667 17508 2683
rect 17474 2599 17508 2611
rect 17474 2520 17508 2539
rect 17570 3509 17604 3528
rect 17570 3437 17604 3449
rect 17570 3365 17604 3381
rect 17570 3293 17604 3313
rect 17570 3221 17604 3245
rect 17570 3149 17604 3177
rect 17570 3077 17604 3109
rect 17570 3007 17604 3041
rect 17570 2939 17604 2971
rect 17570 2871 17604 2899
rect 17570 2803 17604 2827
rect 17570 2735 17604 2755
rect 17570 2667 17604 2683
rect 17570 2599 17604 2611
rect 17570 2486 17604 2539
rect 17666 3509 17700 3582
rect 17666 3437 17700 3449
rect 17666 3365 17700 3381
rect 17666 3293 17700 3313
rect 17666 3221 17700 3245
rect 17666 3149 17700 3177
rect 17666 3077 17700 3109
rect 17666 3007 17700 3041
rect 17666 2939 17700 2971
rect 17666 2871 17700 2899
rect 17666 2803 17700 2827
rect 17666 2735 17700 2755
rect 17666 2667 17700 2683
rect 17666 2599 17700 2611
rect 17666 2520 17700 2539
rect 17762 3509 17796 3528
rect 17762 3437 17796 3449
rect 17762 3365 17796 3381
rect 17762 3293 17796 3313
rect 17762 3221 17796 3245
rect 17762 3149 17796 3177
rect 17762 3077 17796 3109
rect 17762 3007 17796 3041
rect 17762 2939 17796 2971
rect 17762 2871 17796 2899
rect 17762 2803 17796 2827
rect 17762 2735 17796 2755
rect 17762 2667 17796 2683
rect 17762 2599 17796 2611
rect 17762 2486 17796 2539
rect 17858 3509 17892 3582
rect 17858 3437 17892 3449
rect 17858 3365 17892 3381
rect 17858 3293 17892 3313
rect 17858 3221 17892 3245
rect 17858 3149 17892 3177
rect 17858 3077 17892 3109
rect 17858 3007 17892 3041
rect 17858 2939 17892 2971
rect 17858 2871 17892 2899
rect 17858 2803 17892 2827
rect 17858 2735 17892 2755
rect 17858 2667 17892 2683
rect 17858 2599 17892 2611
rect 17858 2520 17892 2539
rect 17954 3509 17988 3528
rect 17954 3437 17988 3449
rect 17954 3365 17988 3381
rect 17954 3293 17988 3313
rect 17954 3221 17988 3245
rect 17954 3149 17988 3177
rect 17954 3077 17988 3109
rect 17954 3007 17988 3041
rect 17954 2939 17988 2971
rect 17954 2871 17988 2899
rect 17954 2803 17988 2827
rect 17954 2735 17988 2755
rect 17954 2667 17988 2683
rect 17954 2599 17988 2611
rect 17954 2486 17988 2539
rect 18050 3509 18084 3582
rect 18050 3437 18084 3449
rect 18050 3365 18084 3381
rect 18050 3293 18084 3313
rect 18050 3221 18084 3245
rect 18050 3149 18084 3177
rect 18050 3077 18084 3109
rect 18050 3007 18084 3041
rect 18050 2939 18084 2971
rect 18050 2871 18084 2899
rect 18050 2803 18084 2827
rect 18050 2735 18084 2755
rect 18050 2667 18084 2683
rect 18050 2599 18084 2611
rect 18050 2520 18084 2539
rect 18146 3509 18180 3528
rect 18146 3437 18180 3449
rect 18146 3365 18180 3381
rect 18146 3293 18180 3313
rect 18146 3221 18180 3245
rect 18146 3149 18180 3177
rect 18146 3077 18180 3109
rect 18146 3007 18180 3041
rect 18146 2939 18180 2971
rect 18146 2871 18180 2899
rect 18146 2803 18180 2827
rect 18146 2735 18180 2755
rect 18146 2667 18180 2683
rect 18146 2599 18180 2611
rect 18146 2486 18180 2539
rect 18242 3509 18276 3582
rect 18672 3574 20050 3608
rect 21640 3604 21686 3770
rect 23462 3819 23496 4038
rect 24054 4030 24856 4064
rect 25258 4058 25292 4135
rect 25354 5105 25388 5166
rect 25354 5033 25388 5045
rect 25354 4961 25388 4977
rect 25354 4889 25388 4909
rect 25354 4817 25388 4841
rect 25354 4745 25388 4773
rect 25354 4673 25388 4705
rect 25354 4603 25388 4637
rect 25354 4535 25388 4567
rect 25354 4467 25388 4495
rect 25354 4399 25388 4423
rect 25354 4331 25388 4351
rect 25354 4263 25388 4279
rect 25354 4195 25388 4207
rect 25354 4116 25388 4135
rect 25450 5105 25484 5124
rect 25450 5033 25484 5045
rect 25450 4961 25484 4977
rect 25450 4889 25484 4909
rect 25450 4817 25484 4841
rect 25450 4745 25484 4773
rect 25450 4673 25484 4705
rect 25450 4603 25484 4637
rect 25450 4535 25484 4567
rect 25450 4467 25484 4495
rect 25450 4399 25484 4423
rect 25450 4331 25484 4351
rect 25450 4263 25484 4279
rect 25450 4195 25484 4207
rect 25450 4058 25484 4135
rect 25546 5105 25580 5166
rect 25546 5033 25580 5045
rect 25546 4961 25580 4977
rect 25546 4889 25580 4909
rect 25546 4817 25580 4841
rect 25546 4745 25580 4773
rect 25546 4673 25580 4705
rect 25546 4603 25580 4637
rect 25546 4535 25580 4567
rect 25546 4467 25580 4495
rect 25546 4399 25580 4423
rect 25546 4331 25580 4351
rect 25546 4263 25580 4279
rect 25546 4195 25580 4207
rect 25546 4116 25580 4135
rect 25642 5105 25676 5124
rect 25642 5033 25676 5045
rect 25642 4961 25676 4977
rect 25642 4889 25676 4909
rect 25642 4817 25676 4841
rect 25642 4745 25676 4773
rect 25642 4673 25676 4705
rect 25642 4603 25676 4637
rect 25642 4535 25676 4567
rect 25642 4467 25676 4495
rect 25642 4399 25676 4423
rect 25642 4331 25676 4351
rect 25642 4263 25676 4279
rect 25642 4195 25676 4207
rect 25642 4058 25676 4135
rect 25738 5105 25772 5166
rect 25738 5033 25772 5045
rect 25738 4961 25772 4977
rect 25738 4889 25772 4909
rect 25738 4817 25772 4841
rect 25738 4745 25772 4773
rect 25738 4673 25772 4705
rect 25738 4603 25772 4637
rect 25738 4535 25772 4567
rect 25738 4467 25772 4495
rect 25738 4399 25772 4423
rect 25738 4331 25772 4351
rect 25738 4263 25772 4279
rect 25738 4195 25772 4207
rect 25738 4116 25772 4135
rect 25834 5105 25868 5124
rect 25834 5033 25868 5045
rect 25834 4961 25868 4977
rect 25834 4889 25868 4909
rect 25834 4817 25868 4841
rect 25834 4745 25868 4773
rect 25834 4673 25868 4705
rect 25834 4603 25868 4637
rect 25834 4535 25868 4567
rect 25834 4467 25868 4495
rect 25834 4399 25868 4423
rect 25834 4331 25868 4351
rect 25834 4263 25868 4279
rect 25834 4195 25868 4207
rect 25834 4058 25868 4135
rect 25930 5105 25964 5166
rect 25930 5033 25964 5045
rect 25930 4961 25964 4977
rect 25930 4889 25964 4909
rect 25930 4817 25964 4841
rect 25930 4745 25964 4773
rect 25930 4673 25964 4705
rect 25930 4603 25964 4637
rect 25930 4535 25964 4567
rect 25930 4467 25964 4495
rect 25930 4399 25964 4423
rect 25930 4331 25964 4351
rect 25930 4263 25964 4279
rect 25930 4195 25964 4207
rect 25930 4116 25964 4135
rect 26026 5105 26060 5124
rect 26026 5033 26060 5045
rect 26026 4961 26060 4977
rect 26026 4889 26060 4909
rect 26026 4817 26060 4841
rect 26026 4745 26060 4773
rect 26026 4673 26060 4705
rect 26026 4603 26060 4637
rect 26026 4535 26060 4567
rect 26026 4467 26060 4495
rect 26026 4399 26060 4423
rect 26026 4331 26060 4351
rect 26026 4263 26060 4279
rect 26026 4195 26060 4207
rect 26026 4058 26060 4135
rect 26122 5105 26156 5166
rect 26122 5033 26156 5045
rect 26122 4961 26156 4977
rect 26122 4889 26156 4909
rect 26122 4817 26156 4841
rect 26122 4745 26156 4773
rect 26122 4673 26156 4705
rect 26122 4603 26156 4637
rect 26122 4535 26156 4567
rect 26122 4467 26156 4495
rect 26122 4399 26156 4423
rect 26122 4331 26156 4351
rect 26122 4263 26156 4279
rect 26122 4195 26156 4207
rect 26122 4116 26156 4135
rect 26218 5105 26252 5124
rect 26218 5033 26252 5045
rect 26218 4961 26252 4977
rect 26218 4889 26252 4909
rect 26218 4817 26252 4841
rect 26218 4745 26252 4773
rect 26218 4673 26252 4705
rect 26218 4603 26252 4637
rect 26218 4535 26252 4567
rect 26218 4467 26252 4495
rect 26218 4399 26252 4423
rect 26218 4331 26252 4351
rect 26218 4263 26252 4279
rect 26218 4195 26252 4207
rect 26218 4058 26252 4135
rect 26314 5105 26348 5166
rect 26314 5033 26348 5045
rect 26314 4961 26348 4977
rect 26314 4889 26348 4909
rect 26314 4817 26348 4841
rect 26314 4745 26348 4773
rect 26314 4673 26348 4705
rect 26314 4603 26348 4637
rect 26314 4535 26348 4567
rect 26314 4467 26348 4495
rect 26314 4399 26348 4423
rect 26314 4331 26348 4351
rect 26314 4263 26348 4279
rect 26314 4195 26348 4207
rect 26314 4116 26348 4135
rect 26410 5105 26444 5124
rect 26410 5033 26444 5045
rect 26410 4961 26444 4977
rect 26410 4889 26444 4909
rect 26410 4817 26444 4841
rect 26410 4745 26444 4773
rect 26410 4673 26444 4705
rect 26410 4603 26444 4637
rect 26410 4535 26444 4567
rect 26410 4467 26444 4495
rect 26410 4399 26444 4423
rect 26410 4331 26444 4351
rect 26410 4263 26444 4279
rect 26410 4195 26444 4207
rect 26410 4058 26444 4135
rect 26506 5105 26540 5166
rect 26826 5172 28780 5194
rect 26506 5033 26540 5045
rect 26506 4961 26540 4977
rect 26506 4889 26540 4909
rect 26506 4817 26540 4841
rect 26506 4745 26540 4773
rect 26506 4673 26540 4705
rect 26506 4603 26540 4637
rect 26506 4535 26540 4567
rect 26506 4467 26540 4495
rect 26506 4399 26540 4423
rect 26506 4331 26540 4351
rect 26506 4263 26540 4279
rect 26506 4195 26540 4207
rect 26506 4116 26540 4135
rect 26602 5105 26636 5124
rect 26602 5033 26636 5045
rect 26602 4961 26636 4977
rect 26602 4889 26636 4909
rect 26602 4817 26636 4841
rect 26602 4745 26636 4773
rect 26602 4673 26636 4705
rect 26602 4603 26636 4637
rect 26602 4535 26636 4567
rect 26602 4467 26636 4495
rect 26602 4399 26636 4423
rect 26602 4331 26636 4351
rect 26602 4263 26636 4279
rect 26602 4195 26636 4207
rect 26602 4058 26636 4135
rect 26826 5099 26860 5172
rect 26826 5027 26860 5039
rect 26826 4955 26860 4971
rect 26826 4883 26860 4903
rect 26826 4811 26860 4835
rect 26826 4739 26860 4767
rect 26826 4667 26860 4699
rect 26826 4597 26860 4631
rect 26826 4529 26860 4561
rect 26826 4461 26860 4489
rect 26826 4393 26860 4417
rect 26826 4325 26860 4345
rect 26826 4257 26860 4273
rect 26826 4189 26860 4201
rect 26826 4110 26860 4129
rect 26922 5099 26956 5118
rect 26922 5027 26956 5039
rect 26922 4955 26956 4971
rect 26922 4883 26956 4903
rect 26922 4811 26956 4835
rect 26922 4739 26956 4767
rect 26922 4667 26956 4699
rect 26922 4597 26956 4631
rect 26922 4529 26956 4561
rect 26922 4461 26956 4489
rect 26922 4393 26956 4417
rect 26922 4325 26956 4345
rect 26922 4257 26956 4273
rect 26922 4189 26956 4201
rect 23990 3925 24006 3959
rect 24040 3925 24056 3959
rect 23302 3670 23318 3704
rect 23352 3670 23368 3704
rect 23462 3604 23496 3785
rect 24276 3817 24314 4030
rect 25258 4024 26636 4058
rect 26922 4064 26956 4129
rect 27018 5099 27052 5172
rect 27018 5027 27052 5039
rect 27018 4955 27052 4971
rect 27018 4883 27052 4903
rect 27018 4811 27052 4835
rect 27018 4739 27052 4767
rect 27018 4667 27052 4699
rect 27018 4597 27052 4631
rect 27018 4529 27052 4561
rect 27018 4461 27052 4489
rect 27018 4393 27052 4417
rect 27018 4325 27052 4345
rect 27018 4257 27052 4273
rect 27018 4189 27052 4201
rect 27018 4110 27052 4129
rect 27114 5099 27148 5118
rect 27114 5027 27148 5039
rect 27114 4955 27148 4971
rect 27114 4883 27148 4903
rect 27114 4811 27148 4835
rect 27114 4739 27148 4767
rect 27114 4667 27148 4699
rect 27114 4597 27148 4631
rect 27114 4529 27148 4561
rect 27114 4461 27148 4489
rect 27114 4393 27148 4417
rect 27114 4325 27148 4345
rect 27114 4257 27148 4273
rect 27114 4189 27148 4201
rect 27114 4064 27148 4129
rect 27210 5099 27244 5172
rect 27210 5027 27244 5039
rect 27210 4955 27244 4971
rect 27210 4883 27244 4903
rect 27210 4811 27244 4835
rect 27210 4739 27244 4767
rect 27210 4667 27244 4699
rect 27210 4597 27244 4631
rect 27210 4529 27244 4561
rect 27210 4461 27244 4489
rect 27210 4393 27244 4417
rect 27210 4325 27244 4345
rect 27210 4257 27244 4273
rect 27210 4189 27244 4201
rect 27210 4110 27244 4129
rect 27306 5099 27340 5118
rect 27306 5027 27340 5039
rect 27306 4955 27340 4971
rect 27306 4883 27340 4903
rect 27306 4811 27340 4835
rect 27306 4739 27340 4767
rect 27306 4667 27340 4699
rect 27306 4597 27340 4631
rect 27306 4529 27340 4561
rect 27306 4461 27340 4489
rect 27306 4393 27340 4417
rect 27306 4325 27340 4345
rect 27306 4257 27340 4273
rect 27306 4189 27340 4201
rect 27306 4064 27340 4129
rect 27402 5099 27436 5172
rect 27402 5027 27436 5039
rect 27402 4955 27436 4971
rect 27402 4883 27436 4903
rect 27402 4811 27436 4835
rect 27402 4739 27436 4767
rect 27402 4667 27436 4699
rect 27402 4597 27436 4631
rect 27402 4529 27436 4561
rect 27402 4461 27436 4489
rect 27402 4393 27436 4417
rect 27402 4325 27436 4345
rect 27402 4257 27436 4273
rect 27402 4189 27436 4201
rect 27402 4110 27436 4129
rect 27498 5099 27532 5118
rect 27498 5027 27532 5039
rect 27498 4955 27532 4971
rect 27498 4883 27532 4903
rect 27498 4811 27532 4835
rect 27498 4739 27532 4767
rect 27498 4667 27532 4699
rect 27498 4597 27532 4631
rect 27498 4529 27532 4561
rect 27498 4461 27532 4489
rect 27498 4393 27532 4417
rect 27498 4325 27532 4345
rect 27498 4257 27532 4273
rect 27498 4189 27532 4201
rect 27498 4064 27532 4129
rect 27594 5099 27628 5172
rect 27594 5027 27628 5039
rect 27594 4955 27628 4971
rect 27594 4883 27628 4903
rect 27594 4811 27628 4835
rect 27594 4739 27628 4767
rect 27594 4667 27628 4699
rect 27594 4597 27628 4631
rect 27594 4529 27628 4561
rect 27594 4461 27628 4489
rect 27594 4393 27628 4417
rect 27594 4325 27628 4345
rect 27594 4257 27628 4273
rect 27594 4189 27628 4201
rect 27594 4110 27628 4129
rect 27690 5099 27724 5118
rect 27690 5027 27724 5039
rect 27690 4955 27724 4971
rect 27690 4883 27724 4903
rect 27690 4811 27724 4835
rect 27690 4739 27724 4767
rect 27690 4667 27724 4699
rect 27690 4597 27724 4631
rect 27690 4529 27724 4561
rect 27690 4461 27724 4489
rect 27690 4393 27724 4417
rect 27690 4325 27724 4345
rect 27690 4257 27724 4273
rect 27690 4189 27724 4201
rect 27690 4064 27724 4129
rect 27786 5099 27820 5172
rect 27786 5027 27820 5039
rect 27786 4955 27820 4971
rect 27786 4883 27820 4903
rect 27786 4811 27820 4835
rect 27786 4739 27820 4767
rect 27786 4667 27820 4699
rect 27786 4597 27820 4631
rect 27786 4529 27820 4561
rect 27786 4461 27820 4489
rect 27786 4393 27820 4417
rect 27786 4325 27820 4345
rect 27786 4257 27820 4273
rect 27786 4189 27820 4201
rect 27786 4110 27820 4129
rect 27882 5099 27916 5118
rect 27882 5027 27916 5039
rect 27882 4955 27916 4971
rect 27882 4883 27916 4903
rect 27882 4811 27916 4835
rect 27882 4739 27916 4767
rect 27882 4667 27916 4699
rect 27882 4597 27916 4631
rect 27882 4529 27916 4561
rect 27882 4461 27916 4489
rect 27882 4393 27916 4417
rect 27882 4325 27916 4345
rect 27882 4257 27916 4273
rect 27882 4189 27916 4201
rect 27882 4064 27916 4129
rect 27978 5099 28012 5172
rect 27978 5027 28012 5039
rect 27978 4955 28012 4971
rect 27978 4883 28012 4903
rect 27978 4811 28012 4835
rect 27978 4739 28012 4767
rect 27978 4667 28012 4699
rect 27978 4597 28012 4631
rect 27978 4529 28012 4561
rect 27978 4461 28012 4489
rect 27978 4393 28012 4417
rect 27978 4325 28012 4345
rect 27978 4257 28012 4273
rect 27978 4189 28012 4201
rect 27978 4110 28012 4129
rect 28074 5099 28108 5118
rect 28074 5027 28108 5039
rect 28074 4955 28108 4971
rect 28074 4883 28108 4903
rect 28074 4811 28108 4835
rect 28074 4739 28108 4767
rect 28074 4667 28108 4699
rect 28074 4597 28108 4631
rect 28074 4529 28108 4561
rect 28074 4461 28108 4489
rect 28074 4393 28108 4417
rect 28074 4325 28108 4345
rect 28074 4257 28108 4273
rect 28074 4189 28108 4201
rect 28074 4064 28108 4129
rect 28170 5099 28204 5172
rect 28170 5027 28204 5039
rect 28170 4955 28204 4971
rect 28170 4883 28204 4903
rect 28170 4811 28204 4835
rect 28170 4739 28204 4767
rect 28170 4667 28204 4699
rect 28170 4597 28204 4631
rect 28170 4529 28204 4561
rect 28170 4461 28204 4489
rect 28170 4393 28204 4417
rect 28170 4325 28204 4345
rect 28170 4257 28204 4273
rect 28170 4189 28204 4201
rect 28170 4110 28204 4129
rect 28266 5099 28300 5118
rect 28266 5027 28300 5039
rect 28266 4955 28300 4971
rect 28266 4883 28300 4903
rect 28266 4811 28300 4835
rect 28266 4739 28300 4767
rect 28266 4667 28300 4699
rect 28266 4597 28300 4631
rect 28266 4529 28300 4561
rect 28266 4461 28300 4489
rect 28266 4393 28300 4417
rect 28266 4325 28300 4345
rect 28266 4257 28300 4273
rect 28266 4189 28300 4201
rect 28266 4064 28300 4129
rect 28362 5099 28396 5172
rect 28362 5027 28396 5039
rect 28362 4955 28396 4971
rect 28362 4883 28396 4903
rect 28362 4811 28396 4835
rect 28362 4739 28396 4767
rect 28362 4667 28396 4699
rect 28362 4597 28396 4631
rect 28362 4529 28396 4561
rect 28362 4461 28396 4489
rect 28362 4393 28396 4417
rect 28362 4325 28396 4345
rect 28362 4257 28396 4273
rect 28362 4189 28396 4201
rect 28362 4110 28396 4129
rect 28458 5099 28492 5118
rect 28458 5027 28492 5039
rect 28458 4955 28492 4971
rect 28458 4883 28492 4903
rect 28458 4811 28492 4835
rect 28458 4739 28492 4767
rect 28458 4667 28492 4699
rect 28458 4597 28492 4631
rect 28458 4529 28492 4561
rect 28458 4461 28492 4489
rect 28458 4393 28492 4417
rect 28458 4325 28492 4345
rect 28458 4257 28492 4273
rect 28458 4189 28492 4201
rect 28458 4064 28492 4129
rect 28554 5099 28588 5172
rect 28554 5027 28588 5039
rect 28554 4955 28588 4971
rect 28554 4883 28588 4903
rect 28554 4811 28588 4835
rect 28554 4739 28588 4767
rect 28554 4667 28588 4699
rect 28554 4597 28588 4631
rect 28554 4529 28588 4561
rect 28554 4461 28588 4489
rect 28554 4393 28588 4417
rect 28554 4325 28588 4345
rect 28554 4257 28588 4273
rect 28554 4189 28588 4201
rect 28554 4110 28588 4129
rect 28650 5099 28684 5118
rect 28650 5027 28684 5039
rect 28650 4955 28684 4971
rect 28650 4883 28684 4903
rect 28650 4811 28684 4835
rect 28650 4739 28684 4767
rect 28650 4667 28684 4699
rect 28650 4597 28684 4631
rect 28650 4529 28684 4561
rect 28650 4461 28684 4489
rect 28650 4393 28684 4417
rect 28650 4325 28684 4345
rect 28650 4257 28684 4273
rect 28650 4189 28684 4201
rect 28650 4064 28684 4129
rect 28746 5099 28780 5172
rect 28746 5027 28780 5039
rect 28746 4955 28780 4971
rect 28746 4883 28780 4903
rect 28746 4811 28780 4835
rect 28746 4739 28780 4767
rect 28746 4667 28780 4699
rect 28746 4597 28780 4631
rect 28746 4529 28780 4561
rect 28746 4461 28780 4489
rect 28746 4393 28780 4417
rect 28746 4325 28780 4345
rect 28746 4257 28780 4273
rect 28746 4189 28780 4201
rect 28746 4110 28780 4129
rect 26922 4030 28684 4064
rect 25194 3919 25210 3953
rect 25244 3919 25260 3953
rect 24276 3783 24278 3817
rect 24312 3783 24314 3817
rect 23994 3700 24010 3734
rect 24044 3700 24060 3734
rect 24276 3614 24314 3783
rect 25928 3804 25968 4024
rect 26858 3913 26874 3947
rect 26908 3913 26924 3947
rect 25928 3770 25931 3804
rect 25965 3770 25968 3804
rect 25192 3656 25208 3690
rect 25242 3656 25258 3690
rect 18242 3437 18276 3449
rect 18242 3365 18276 3381
rect 18242 3293 18276 3313
rect 18242 3221 18276 3245
rect 18242 3149 18276 3177
rect 18242 3077 18276 3109
rect 18242 3007 18276 3041
rect 18242 2939 18276 2971
rect 18242 2871 18276 2899
rect 18242 2803 18276 2827
rect 18242 2735 18276 2755
rect 18242 2667 18276 2683
rect 18242 2599 18276 2611
rect 18242 2520 18276 2539
rect 18338 3509 18372 3528
rect 18338 3437 18372 3449
rect 18338 3365 18372 3381
rect 18338 3293 18372 3313
rect 18338 3221 18372 3245
rect 18338 3149 18372 3177
rect 18338 3077 18372 3109
rect 18338 3007 18372 3041
rect 18338 2939 18372 2971
rect 18338 2871 18372 2899
rect 18338 2803 18372 2827
rect 18338 2735 18372 2755
rect 18338 2667 18372 2683
rect 18338 2599 18372 2611
rect 18338 2486 18372 2539
rect 17378 2460 18372 2486
rect 18576 3505 18610 3524
rect 18576 3433 18610 3445
rect 18576 3361 18610 3377
rect 18576 3289 18610 3309
rect 18576 3217 18610 3241
rect 18576 3145 18610 3173
rect 18576 3073 18610 3105
rect 18576 3003 18610 3037
rect 18576 2935 18610 2967
rect 18576 2867 18610 2895
rect 18576 2799 18610 2823
rect 18576 2731 18610 2751
rect 18576 2663 18610 2679
rect 18576 2595 18610 2607
rect 18576 2474 18610 2535
rect 18672 3505 18706 3574
rect 18672 3433 18706 3445
rect 18672 3361 18706 3377
rect 18672 3289 18706 3309
rect 18672 3217 18706 3241
rect 18672 3145 18706 3173
rect 18672 3073 18706 3105
rect 18672 3003 18706 3037
rect 18672 2935 18706 2967
rect 18672 2867 18706 2895
rect 18672 2799 18706 2823
rect 18672 2731 18706 2751
rect 18672 2663 18706 2679
rect 18672 2595 18706 2607
rect 18672 2516 18706 2535
rect 18768 3505 18802 3524
rect 18768 3433 18802 3445
rect 18768 3361 18802 3377
rect 18768 3289 18802 3309
rect 18768 3217 18802 3241
rect 18768 3145 18802 3173
rect 18768 3073 18802 3105
rect 18768 3003 18802 3037
rect 18768 2935 18802 2967
rect 18768 2867 18802 2895
rect 18768 2799 18802 2823
rect 18768 2731 18802 2751
rect 18768 2663 18802 2679
rect 18768 2595 18802 2607
rect 18768 2474 18802 2535
rect 18864 3505 18898 3574
rect 18864 3433 18898 3445
rect 18864 3361 18898 3377
rect 18864 3289 18898 3309
rect 18864 3217 18898 3241
rect 18864 3145 18898 3173
rect 18864 3073 18898 3105
rect 18864 3003 18898 3037
rect 18864 2935 18898 2967
rect 18864 2867 18898 2895
rect 18864 2799 18898 2823
rect 18864 2731 18898 2751
rect 18864 2663 18898 2679
rect 18864 2595 18898 2607
rect 18864 2516 18898 2535
rect 18960 3505 18994 3524
rect 18960 3433 18994 3445
rect 18960 3361 18994 3377
rect 18960 3289 18994 3309
rect 18960 3217 18994 3241
rect 18960 3145 18994 3173
rect 18960 3073 18994 3105
rect 18960 3003 18994 3037
rect 18960 2935 18994 2967
rect 18960 2867 18994 2895
rect 18960 2799 18994 2823
rect 18960 2731 18994 2751
rect 18960 2663 18994 2679
rect 18960 2595 18994 2607
rect 18960 2474 18994 2535
rect 19056 3505 19090 3574
rect 19056 3433 19090 3445
rect 19056 3361 19090 3377
rect 19056 3289 19090 3309
rect 19056 3217 19090 3241
rect 19056 3145 19090 3173
rect 19056 3073 19090 3105
rect 19056 3003 19090 3037
rect 19056 2935 19090 2967
rect 19056 2867 19090 2895
rect 19056 2799 19090 2823
rect 19056 2731 19090 2751
rect 19056 2663 19090 2679
rect 19056 2595 19090 2607
rect 19056 2516 19090 2535
rect 19152 3505 19186 3524
rect 19152 3433 19186 3445
rect 19152 3361 19186 3377
rect 19152 3289 19186 3309
rect 19152 3217 19186 3241
rect 19152 3145 19186 3173
rect 19152 3073 19186 3105
rect 19152 3003 19186 3037
rect 19152 2935 19186 2967
rect 19152 2867 19186 2895
rect 19152 2799 19186 2823
rect 19152 2731 19186 2751
rect 19152 2663 19186 2679
rect 19152 2595 19186 2607
rect 19152 2474 19186 2535
rect 19248 3505 19282 3574
rect 19248 3433 19282 3445
rect 19248 3361 19282 3377
rect 19248 3289 19282 3309
rect 19248 3217 19282 3241
rect 19248 3145 19282 3173
rect 19248 3073 19282 3105
rect 19248 3003 19282 3037
rect 19248 2935 19282 2967
rect 19248 2867 19282 2895
rect 19248 2799 19282 2823
rect 19248 2731 19282 2751
rect 19248 2663 19282 2679
rect 19248 2595 19282 2607
rect 19248 2516 19282 2535
rect 19344 3505 19378 3524
rect 19344 3433 19378 3445
rect 19344 3361 19378 3377
rect 19344 3289 19378 3309
rect 19344 3217 19378 3241
rect 19344 3145 19378 3173
rect 19344 3073 19378 3105
rect 19344 3003 19378 3037
rect 19344 2935 19378 2967
rect 19344 2867 19378 2895
rect 19344 2799 19378 2823
rect 19344 2731 19378 2751
rect 19344 2663 19378 2679
rect 19344 2595 19378 2607
rect 19344 2474 19378 2535
rect 19440 3505 19474 3574
rect 19440 3433 19474 3445
rect 19440 3361 19474 3377
rect 19440 3289 19474 3309
rect 19440 3217 19474 3241
rect 19440 3145 19474 3173
rect 19440 3073 19474 3105
rect 19440 3003 19474 3037
rect 19440 2935 19474 2967
rect 19440 2867 19474 2895
rect 19440 2799 19474 2823
rect 19440 2731 19474 2751
rect 19440 2663 19474 2679
rect 19440 2595 19474 2607
rect 19440 2516 19474 2535
rect 19536 3505 19570 3524
rect 19536 3433 19570 3445
rect 19536 3361 19570 3377
rect 19536 3289 19570 3309
rect 19536 3217 19570 3241
rect 19536 3145 19570 3173
rect 19536 3073 19570 3105
rect 19536 3003 19570 3037
rect 19536 2935 19570 2967
rect 19536 2867 19570 2895
rect 19536 2799 19570 2823
rect 19536 2731 19570 2751
rect 19536 2663 19570 2679
rect 19536 2595 19570 2607
rect 19536 2474 19570 2535
rect 19632 3505 19666 3574
rect 19632 3433 19666 3445
rect 19632 3361 19666 3377
rect 19632 3289 19666 3309
rect 19632 3217 19666 3241
rect 19632 3145 19666 3173
rect 19632 3073 19666 3105
rect 19632 3003 19666 3037
rect 19632 2935 19666 2967
rect 19632 2867 19666 2895
rect 19632 2799 19666 2823
rect 19632 2731 19666 2751
rect 19632 2663 19666 2679
rect 19632 2595 19666 2607
rect 19632 2516 19666 2535
rect 19728 3505 19762 3524
rect 19728 3433 19762 3445
rect 19728 3361 19762 3377
rect 19728 3289 19762 3309
rect 19728 3217 19762 3241
rect 19728 3145 19762 3173
rect 19728 3073 19762 3105
rect 19728 3003 19762 3037
rect 19728 2935 19762 2967
rect 19728 2867 19762 2895
rect 19728 2799 19762 2823
rect 19728 2731 19762 2751
rect 19728 2663 19762 2679
rect 19728 2595 19762 2607
rect 19728 2474 19762 2535
rect 19824 3505 19858 3574
rect 19824 3433 19858 3445
rect 19824 3361 19858 3377
rect 19824 3289 19858 3309
rect 19824 3217 19858 3241
rect 19824 3145 19858 3173
rect 19824 3073 19858 3105
rect 19824 3003 19858 3037
rect 19824 2935 19858 2967
rect 19824 2867 19858 2895
rect 19824 2799 19858 2823
rect 19824 2731 19858 2751
rect 19824 2663 19858 2679
rect 19824 2595 19858 2607
rect 19824 2516 19858 2535
rect 19920 3505 19954 3524
rect 19920 3433 19954 3445
rect 19920 3361 19954 3377
rect 19920 3289 19954 3309
rect 19920 3217 19954 3241
rect 19920 3145 19954 3173
rect 19920 3073 19954 3105
rect 19920 3003 19954 3037
rect 19920 2935 19954 2967
rect 19920 2867 19954 2895
rect 19920 2799 19954 2823
rect 19920 2731 19954 2751
rect 19920 2663 19954 2679
rect 19920 2595 19954 2607
rect 19920 2474 19954 2535
rect 20016 3505 20050 3574
rect 20340 3570 22104 3604
rect 23270 3570 23688 3604
rect 20016 3433 20050 3445
rect 20016 3361 20050 3377
rect 20016 3289 20050 3309
rect 20016 3217 20050 3241
rect 20016 3145 20050 3173
rect 20016 3073 20050 3105
rect 20016 3003 20050 3037
rect 20016 2935 20050 2967
rect 20016 2867 20050 2895
rect 20016 2799 20050 2823
rect 20016 2731 20050 2751
rect 20016 2663 20050 2679
rect 20016 2595 20050 2607
rect 20016 2516 20050 2535
rect 20244 3513 20278 3532
rect 20244 3441 20278 3453
rect 20244 3369 20278 3385
rect 20244 3297 20278 3317
rect 20244 3225 20278 3249
rect 20244 3153 20278 3181
rect 20244 3081 20278 3113
rect 20244 3011 20278 3045
rect 20244 2943 20278 2975
rect 20244 2875 20278 2903
rect 20244 2807 20278 2831
rect 20244 2739 20278 2759
rect 20244 2671 20278 2687
rect 20244 2603 20278 2615
rect 20244 2482 20278 2543
rect 20340 3513 20374 3570
rect 20340 3441 20374 3453
rect 20340 3369 20374 3385
rect 20340 3297 20374 3317
rect 20340 3225 20374 3249
rect 20340 3153 20374 3181
rect 20340 3081 20374 3113
rect 20340 3011 20374 3045
rect 20340 2943 20374 2975
rect 20340 2875 20374 2903
rect 20340 2807 20374 2831
rect 20340 2739 20374 2759
rect 20340 2671 20374 2687
rect 20340 2603 20374 2615
rect 20340 2524 20374 2543
rect 20436 3513 20470 3532
rect 20436 3441 20470 3453
rect 20436 3369 20470 3385
rect 20436 3297 20470 3317
rect 20436 3225 20470 3249
rect 20436 3153 20470 3181
rect 20436 3081 20470 3113
rect 20436 3011 20470 3045
rect 20436 2943 20470 2975
rect 20436 2875 20470 2903
rect 20436 2807 20470 2831
rect 20436 2739 20470 2759
rect 20436 2671 20470 2687
rect 20436 2603 20470 2615
rect 20436 2482 20470 2543
rect 20532 3513 20566 3570
rect 20532 3441 20566 3453
rect 20532 3369 20566 3385
rect 20532 3297 20566 3317
rect 20532 3225 20566 3249
rect 20532 3153 20566 3181
rect 20532 3081 20566 3113
rect 20532 3011 20566 3045
rect 20532 2943 20566 2975
rect 20532 2875 20566 2903
rect 20532 2807 20566 2831
rect 20532 2739 20566 2759
rect 20532 2671 20566 2687
rect 20532 2603 20566 2615
rect 20532 2524 20566 2543
rect 20628 3513 20662 3532
rect 20628 3441 20662 3453
rect 20628 3369 20662 3385
rect 20628 3297 20662 3317
rect 20628 3225 20662 3249
rect 20628 3153 20662 3181
rect 20628 3081 20662 3113
rect 20628 3011 20662 3045
rect 20628 2943 20662 2975
rect 20628 2875 20662 2903
rect 20628 2807 20662 2831
rect 20628 2739 20662 2759
rect 20628 2671 20662 2687
rect 20628 2603 20662 2615
rect 20628 2482 20662 2543
rect 20724 3513 20758 3570
rect 20724 3441 20758 3453
rect 20724 3369 20758 3385
rect 20724 3297 20758 3317
rect 20724 3225 20758 3249
rect 20724 3153 20758 3181
rect 20724 3081 20758 3113
rect 20724 3011 20758 3045
rect 20724 2943 20758 2975
rect 20724 2875 20758 2903
rect 20724 2807 20758 2831
rect 20724 2739 20758 2759
rect 20724 2671 20758 2687
rect 20724 2603 20758 2615
rect 20724 2524 20758 2543
rect 20820 3513 20854 3532
rect 20820 3441 20854 3453
rect 20820 3369 20854 3385
rect 20820 3297 20854 3317
rect 20820 3225 20854 3249
rect 20820 3153 20854 3181
rect 20820 3081 20854 3113
rect 20820 3011 20854 3045
rect 20820 2943 20854 2975
rect 20820 2875 20854 2903
rect 20820 2807 20854 2831
rect 20820 2739 20854 2759
rect 20820 2671 20854 2687
rect 20820 2603 20854 2615
rect 20820 2482 20854 2543
rect 20916 3513 20950 3570
rect 20916 3441 20950 3453
rect 20916 3369 20950 3385
rect 20916 3297 20950 3317
rect 20916 3225 20950 3249
rect 20916 3153 20950 3181
rect 20916 3081 20950 3113
rect 20916 3011 20950 3045
rect 20916 2943 20950 2975
rect 20916 2875 20950 2903
rect 20916 2807 20950 2831
rect 20916 2739 20950 2759
rect 20916 2671 20950 2687
rect 20916 2603 20950 2615
rect 20916 2524 20950 2543
rect 21012 3513 21046 3532
rect 21012 3441 21046 3453
rect 21012 3369 21046 3385
rect 21012 3297 21046 3317
rect 21012 3225 21046 3249
rect 21012 3153 21046 3181
rect 21012 3081 21046 3113
rect 21012 3011 21046 3045
rect 21012 2943 21046 2975
rect 21012 2875 21046 2903
rect 21012 2807 21046 2831
rect 21012 2739 21046 2759
rect 21012 2671 21046 2687
rect 21012 2603 21046 2615
rect 21012 2482 21046 2543
rect 21108 3513 21142 3570
rect 21108 3441 21142 3453
rect 21108 3369 21142 3385
rect 21108 3297 21142 3317
rect 21108 3225 21142 3249
rect 21108 3153 21142 3181
rect 21108 3081 21142 3113
rect 21108 3011 21142 3045
rect 21108 2943 21142 2975
rect 21108 2875 21142 2903
rect 21108 2807 21142 2831
rect 21108 2739 21142 2759
rect 21108 2671 21142 2687
rect 21108 2603 21142 2615
rect 21108 2524 21142 2543
rect 21204 3513 21238 3532
rect 21204 3441 21238 3453
rect 21204 3369 21238 3385
rect 21204 3297 21238 3317
rect 21204 3225 21238 3249
rect 21204 3153 21238 3181
rect 21204 3081 21238 3113
rect 21204 3011 21238 3045
rect 21204 2943 21238 2975
rect 21204 2875 21238 2903
rect 21204 2807 21238 2831
rect 21204 2739 21238 2759
rect 21204 2671 21238 2687
rect 21204 2603 21238 2615
rect 21204 2482 21238 2543
rect 21300 3513 21334 3570
rect 21300 3441 21334 3453
rect 21300 3369 21334 3385
rect 21300 3297 21334 3317
rect 21300 3225 21334 3249
rect 21300 3153 21334 3181
rect 21300 3081 21334 3113
rect 21300 3011 21334 3045
rect 21300 2943 21334 2975
rect 21300 2875 21334 2903
rect 21300 2807 21334 2831
rect 21300 2739 21334 2759
rect 21300 2671 21334 2687
rect 21300 2603 21334 2615
rect 21300 2524 21334 2543
rect 21396 3513 21430 3532
rect 21396 3441 21430 3453
rect 21396 3369 21430 3385
rect 21396 3297 21430 3317
rect 21396 3225 21430 3249
rect 21396 3153 21430 3181
rect 21396 3081 21430 3113
rect 21396 3011 21430 3045
rect 21396 2943 21430 2975
rect 21396 2875 21430 2903
rect 21396 2807 21430 2831
rect 21396 2739 21430 2759
rect 21396 2671 21430 2687
rect 21396 2603 21430 2615
rect 21396 2482 21430 2543
rect 21492 3513 21526 3570
rect 21492 3441 21526 3453
rect 21492 3369 21526 3385
rect 21492 3297 21526 3317
rect 21492 3225 21526 3249
rect 21492 3153 21526 3181
rect 21492 3081 21526 3113
rect 21492 3011 21526 3045
rect 21492 2943 21526 2975
rect 21492 2875 21526 2903
rect 21492 2807 21526 2831
rect 21492 2739 21526 2759
rect 21492 2671 21526 2687
rect 21492 2603 21526 2615
rect 21492 2524 21526 2543
rect 21588 3513 21622 3532
rect 21588 3441 21622 3453
rect 21588 3369 21622 3385
rect 21588 3297 21622 3317
rect 21588 3225 21622 3249
rect 21588 3153 21622 3181
rect 21588 3081 21622 3113
rect 21588 3011 21622 3045
rect 21588 2943 21622 2975
rect 21588 2875 21622 2903
rect 21588 2807 21622 2831
rect 21588 2739 21622 2759
rect 21588 2671 21622 2687
rect 21588 2603 21622 2615
rect 21588 2482 21622 2543
rect 21684 3513 21718 3570
rect 21684 3441 21718 3453
rect 21684 3369 21718 3385
rect 21684 3297 21718 3317
rect 21684 3225 21718 3249
rect 21684 3153 21718 3181
rect 21684 3081 21718 3113
rect 21684 3011 21718 3045
rect 21684 2943 21718 2975
rect 21684 2875 21718 2903
rect 21684 2807 21718 2831
rect 21684 2739 21718 2759
rect 21684 2671 21718 2687
rect 21684 2603 21718 2615
rect 21684 2524 21718 2543
rect 21780 3513 21814 3532
rect 21780 3441 21814 3453
rect 21780 3369 21814 3385
rect 21780 3297 21814 3317
rect 21780 3225 21814 3249
rect 21780 3153 21814 3181
rect 21780 3081 21814 3113
rect 21780 3011 21814 3045
rect 21780 2943 21814 2975
rect 21780 2875 21814 2903
rect 21780 2807 21814 2831
rect 21780 2739 21814 2759
rect 21780 2671 21814 2687
rect 21780 2603 21814 2615
rect 21780 2482 21814 2543
rect 21876 3513 21910 3570
rect 21876 3441 21910 3453
rect 21876 3369 21910 3385
rect 21876 3297 21910 3317
rect 21876 3225 21910 3249
rect 21876 3153 21910 3181
rect 21876 3081 21910 3113
rect 21876 3011 21910 3045
rect 21876 2943 21910 2975
rect 21876 2875 21910 2903
rect 21876 2807 21910 2831
rect 21876 2739 21910 2759
rect 21876 2671 21910 2687
rect 21876 2603 21910 2615
rect 21876 2524 21910 2543
rect 21972 3513 22006 3532
rect 21972 3441 22006 3453
rect 21972 3369 22006 3385
rect 21972 3297 22006 3317
rect 21972 3225 22006 3249
rect 21972 3153 22006 3181
rect 21972 3081 22006 3113
rect 21972 3011 22006 3045
rect 21972 2943 22006 2975
rect 21972 2875 22006 2903
rect 21972 2807 22006 2831
rect 21972 2739 22006 2759
rect 21972 2671 22006 2687
rect 21972 2603 22006 2615
rect 21972 2482 22006 2543
rect 22068 3513 22102 3570
rect 22068 3441 22102 3453
rect 22068 3369 22102 3385
rect 22068 3297 22102 3317
rect 22068 3225 22102 3249
rect 22068 3153 22102 3181
rect 22068 3081 22102 3113
rect 22068 3011 22102 3045
rect 22068 2943 22102 2975
rect 22068 2875 22102 2903
rect 22068 2807 22102 2831
rect 22068 2739 22102 2759
rect 22068 2671 22102 2687
rect 22068 2603 22102 2615
rect 22068 2524 22102 2543
rect 22164 3513 22198 3532
rect 22164 3441 22198 3453
rect 22164 3369 22198 3385
rect 22164 3297 22198 3317
rect 22164 3225 22198 3249
rect 22164 3153 22198 3181
rect 22164 3081 22198 3113
rect 22164 3011 22198 3045
rect 22164 2943 22198 2975
rect 22164 2875 22198 2903
rect 22164 2807 22198 2831
rect 22164 2739 22198 2759
rect 22164 2671 22198 2687
rect 22164 2603 22198 2615
rect 22164 2482 22198 2543
rect 18576 2460 19966 2474
rect 20244 2460 22198 2482
rect 23174 3517 23208 3536
rect 23174 3445 23208 3457
rect 23174 3373 23208 3389
rect 23174 3301 23208 3321
rect 23174 3229 23208 3253
rect 23174 3157 23208 3185
rect 23174 3085 23208 3117
rect 23174 3015 23208 3049
rect 23174 2947 23208 2979
rect 23174 2879 23208 2907
rect 23174 2811 23208 2835
rect 23174 2743 23208 2763
rect 23174 2675 23208 2691
rect 23174 2607 23208 2619
rect 23174 2480 23208 2547
rect 23270 3517 23304 3570
rect 23270 3445 23304 3457
rect 23270 3373 23304 3389
rect 23270 3301 23304 3321
rect 23270 3229 23304 3253
rect 23270 3157 23304 3185
rect 23270 3085 23304 3117
rect 23270 3015 23304 3049
rect 23270 2947 23304 2979
rect 23270 2879 23304 2907
rect 23270 2811 23304 2835
rect 23270 2743 23304 2763
rect 23270 2675 23304 2691
rect 23270 2607 23304 2619
rect 23270 2528 23304 2547
rect 23366 3517 23400 3536
rect 23366 3445 23400 3457
rect 23366 3373 23400 3389
rect 23366 3301 23400 3321
rect 23366 3229 23400 3253
rect 23366 3157 23400 3185
rect 23366 3085 23400 3117
rect 23366 3015 23400 3049
rect 23366 2947 23400 2979
rect 23366 2879 23400 2907
rect 23366 2811 23400 2835
rect 23366 2743 23400 2763
rect 23366 2675 23400 2691
rect 23366 2607 23400 2619
rect 23366 2480 23400 2547
rect 23462 3517 23496 3570
rect 23462 3445 23496 3457
rect 23462 3373 23496 3389
rect 23462 3301 23496 3321
rect 23462 3229 23496 3253
rect 23462 3157 23496 3185
rect 23462 3085 23496 3117
rect 23462 3015 23496 3049
rect 23462 2947 23496 2979
rect 23462 2879 23496 2907
rect 23462 2811 23496 2835
rect 23462 2743 23496 2763
rect 23462 2675 23496 2691
rect 23462 2607 23496 2619
rect 23462 2528 23496 2547
rect 23558 3517 23592 3536
rect 23558 3445 23592 3457
rect 23558 3373 23592 3389
rect 23558 3301 23592 3321
rect 23558 3229 23592 3253
rect 23558 3157 23592 3185
rect 23558 3085 23592 3117
rect 23558 3015 23592 3049
rect 23558 2947 23592 2979
rect 23558 2879 23592 2907
rect 23558 2811 23592 2835
rect 23558 2743 23592 2763
rect 23558 2675 23592 2691
rect 23558 2607 23592 2619
rect 23558 2480 23592 2547
rect 23654 3517 23688 3570
rect 23962 3580 24764 3614
rect 25928 3606 25968 3770
rect 28128 3802 28174 4030
rect 28128 3768 28134 3802
rect 28168 3768 28174 3802
rect 26860 3654 26876 3688
rect 26910 3654 26926 3688
rect 23654 3445 23688 3457
rect 23654 3373 23688 3389
rect 23654 3301 23688 3321
rect 23654 3229 23688 3253
rect 23654 3157 23688 3185
rect 23654 3085 23688 3117
rect 23654 3015 23688 3049
rect 23654 2947 23688 2979
rect 23654 2879 23688 2907
rect 23654 2811 23688 2835
rect 23654 2743 23688 2763
rect 23654 2675 23688 2691
rect 23654 2607 23688 2619
rect 23654 2528 23688 2547
rect 23866 3507 23900 3526
rect 23866 3435 23900 3447
rect 23866 3363 23900 3379
rect 23866 3291 23900 3311
rect 23866 3219 23900 3243
rect 23866 3147 23900 3175
rect 23866 3075 23900 3107
rect 23866 3005 23900 3039
rect 23866 2937 23900 2969
rect 23866 2869 23900 2897
rect 23866 2801 23900 2825
rect 23866 2733 23900 2753
rect 23866 2665 23900 2681
rect 23866 2597 23900 2609
rect 23174 2468 23592 2480
rect 23866 2484 23900 2537
rect 23962 3507 23996 3580
rect 23962 3435 23996 3447
rect 23962 3363 23996 3379
rect 23962 3291 23996 3311
rect 23962 3219 23996 3243
rect 23962 3147 23996 3175
rect 23962 3075 23996 3107
rect 23962 3005 23996 3039
rect 23962 2937 23996 2969
rect 23962 2869 23996 2897
rect 23962 2801 23996 2825
rect 23962 2733 23996 2753
rect 23962 2665 23996 2681
rect 23962 2597 23996 2609
rect 23962 2518 23996 2537
rect 24058 3507 24092 3526
rect 24058 3435 24092 3447
rect 24058 3363 24092 3379
rect 24058 3291 24092 3311
rect 24058 3219 24092 3243
rect 24058 3147 24092 3175
rect 24058 3075 24092 3107
rect 24058 3005 24092 3039
rect 24058 2937 24092 2969
rect 24058 2869 24092 2897
rect 24058 2801 24092 2825
rect 24058 2733 24092 2753
rect 24058 2665 24092 2681
rect 24058 2597 24092 2609
rect 24058 2484 24092 2537
rect 24154 3507 24188 3580
rect 24154 3435 24188 3447
rect 24154 3363 24188 3379
rect 24154 3291 24188 3311
rect 24154 3219 24188 3243
rect 24154 3147 24188 3175
rect 24154 3075 24188 3107
rect 24154 3005 24188 3039
rect 24154 2937 24188 2969
rect 24154 2869 24188 2897
rect 24154 2801 24188 2825
rect 24154 2733 24188 2753
rect 24154 2665 24188 2681
rect 24154 2597 24188 2609
rect 24154 2518 24188 2537
rect 24250 3507 24284 3526
rect 24250 3435 24284 3447
rect 24250 3363 24284 3379
rect 24250 3291 24284 3311
rect 24250 3219 24284 3243
rect 24250 3147 24284 3175
rect 24250 3075 24284 3107
rect 24250 3005 24284 3039
rect 24250 2937 24284 2969
rect 24250 2869 24284 2897
rect 24250 2801 24284 2825
rect 24250 2733 24284 2753
rect 24250 2665 24284 2681
rect 24250 2597 24284 2609
rect 24250 2484 24284 2537
rect 24346 3507 24380 3580
rect 24346 3435 24380 3447
rect 24346 3363 24380 3379
rect 24346 3291 24380 3311
rect 24346 3219 24380 3243
rect 24346 3147 24380 3175
rect 24346 3075 24380 3107
rect 24346 3005 24380 3039
rect 24346 2937 24380 2969
rect 24346 2869 24380 2897
rect 24346 2801 24380 2825
rect 24346 2733 24380 2753
rect 24346 2665 24380 2681
rect 24346 2597 24380 2609
rect 24346 2518 24380 2537
rect 24442 3507 24476 3526
rect 24442 3435 24476 3447
rect 24442 3363 24476 3379
rect 24442 3291 24476 3311
rect 24442 3219 24476 3243
rect 24442 3147 24476 3175
rect 24442 3075 24476 3107
rect 24442 3005 24476 3039
rect 24442 2937 24476 2969
rect 24442 2869 24476 2897
rect 24442 2801 24476 2825
rect 24442 2733 24476 2753
rect 24442 2665 24476 2681
rect 24442 2597 24476 2609
rect 24442 2484 24476 2537
rect 24538 3507 24572 3580
rect 24538 3435 24572 3447
rect 24538 3363 24572 3379
rect 24538 3291 24572 3311
rect 24538 3219 24572 3243
rect 24538 3147 24572 3175
rect 24538 3075 24572 3107
rect 24538 3005 24572 3039
rect 24538 2937 24572 2969
rect 24538 2869 24572 2897
rect 24538 2801 24572 2825
rect 24538 2733 24572 2753
rect 24538 2665 24572 2681
rect 24538 2597 24572 2609
rect 24538 2518 24572 2537
rect 24634 3507 24668 3526
rect 24634 3435 24668 3447
rect 24634 3363 24668 3379
rect 24634 3291 24668 3311
rect 24634 3219 24668 3243
rect 24634 3147 24668 3175
rect 24634 3075 24668 3107
rect 24634 3005 24668 3039
rect 24634 2937 24668 2969
rect 24634 2869 24668 2897
rect 24634 2801 24668 2825
rect 24634 2733 24668 2753
rect 24634 2665 24668 2681
rect 24634 2597 24668 2609
rect 24634 2484 24668 2537
rect 24730 3507 24764 3580
rect 25160 3572 26538 3606
rect 28128 3602 28174 3768
rect 24730 3435 24764 3447
rect 24730 3363 24764 3379
rect 24730 3291 24764 3311
rect 24730 3219 24764 3243
rect 24730 3147 24764 3175
rect 24730 3075 24764 3107
rect 24730 3005 24764 3039
rect 24730 2937 24764 2969
rect 24730 2869 24764 2897
rect 24730 2801 24764 2825
rect 24730 2733 24764 2753
rect 24730 2665 24764 2681
rect 24730 2597 24764 2609
rect 24730 2518 24764 2537
rect 24826 3507 24860 3526
rect 24826 3435 24860 3447
rect 24826 3363 24860 3379
rect 24826 3291 24860 3311
rect 24826 3219 24860 3243
rect 24826 3147 24860 3175
rect 24826 3075 24860 3107
rect 24826 3005 24860 3039
rect 24826 2937 24860 2969
rect 24826 2869 24860 2897
rect 24826 2801 24860 2825
rect 24826 2733 24860 2753
rect 24826 2665 24860 2681
rect 24826 2597 24860 2609
rect 24826 2484 24860 2537
rect 23866 2468 24860 2484
rect 25064 3503 25098 3522
rect 25064 3431 25098 3443
rect 25064 3359 25098 3375
rect 25064 3287 25098 3307
rect 25064 3215 25098 3239
rect 25064 3143 25098 3171
rect 25064 3071 25098 3103
rect 25064 3001 25098 3035
rect 25064 2933 25098 2965
rect 25064 2865 25098 2893
rect 25064 2797 25098 2821
rect 25064 2729 25098 2749
rect 25064 2661 25098 2677
rect 25064 2593 25098 2605
rect 25064 2472 25098 2533
rect 25160 3503 25194 3572
rect 25160 3431 25194 3443
rect 25160 3359 25194 3375
rect 25160 3287 25194 3307
rect 25160 3215 25194 3239
rect 25160 3143 25194 3171
rect 25160 3071 25194 3103
rect 25160 3001 25194 3035
rect 25160 2933 25194 2965
rect 25160 2865 25194 2893
rect 25160 2797 25194 2821
rect 25160 2729 25194 2749
rect 25160 2661 25194 2677
rect 25160 2593 25194 2605
rect 25160 2514 25194 2533
rect 25256 3503 25290 3522
rect 25256 3431 25290 3443
rect 25256 3359 25290 3375
rect 25256 3287 25290 3307
rect 25256 3215 25290 3239
rect 25256 3143 25290 3171
rect 25256 3071 25290 3103
rect 25256 3001 25290 3035
rect 25256 2933 25290 2965
rect 25256 2865 25290 2893
rect 25256 2797 25290 2821
rect 25256 2729 25290 2749
rect 25256 2661 25290 2677
rect 25256 2593 25290 2605
rect 25256 2472 25290 2533
rect 25352 3503 25386 3572
rect 25352 3431 25386 3443
rect 25352 3359 25386 3375
rect 25352 3287 25386 3307
rect 25352 3215 25386 3239
rect 25352 3143 25386 3171
rect 25352 3071 25386 3103
rect 25352 3001 25386 3035
rect 25352 2933 25386 2965
rect 25352 2865 25386 2893
rect 25352 2797 25386 2821
rect 25352 2729 25386 2749
rect 25352 2661 25386 2677
rect 25352 2593 25386 2605
rect 25352 2514 25386 2533
rect 25448 3503 25482 3522
rect 25448 3431 25482 3443
rect 25448 3359 25482 3375
rect 25448 3287 25482 3307
rect 25448 3215 25482 3239
rect 25448 3143 25482 3171
rect 25448 3071 25482 3103
rect 25448 3001 25482 3035
rect 25448 2933 25482 2965
rect 25448 2865 25482 2893
rect 25448 2797 25482 2821
rect 25448 2729 25482 2749
rect 25448 2661 25482 2677
rect 25448 2593 25482 2605
rect 25448 2472 25482 2533
rect 25544 3503 25578 3572
rect 25544 3431 25578 3443
rect 25544 3359 25578 3375
rect 25544 3287 25578 3307
rect 25544 3215 25578 3239
rect 25544 3143 25578 3171
rect 25544 3071 25578 3103
rect 25544 3001 25578 3035
rect 25544 2933 25578 2965
rect 25544 2865 25578 2893
rect 25544 2797 25578 2821
rect 25544 2729 25578 2749
rect 25544 2661 25578 2677
rect 25544 2593 25578 2605
rect 25544 2514 25578 2533
rect 25640 3503 25674 3522
rect 25640 3431 25674 3443
rect 25640 3359 25674 3375
rect 25640 3287 25674 3307
rect 25640 3215 25674 3239
rect 25640 3143 25674 3171
rect 25640 3071 25674 3103
rect 25640 3001 25674 3035
rect 25640 2933 25674 2965
rect 25640 2865 25674 2893
rect 25640 2797 25674 2821
rect 25640 2729 25674 2749
rect 25640 2661 25674 2677
rect 25640 2593 25674 2605
rect 25640 2472 25674 2533
rect 25736 3503 25770 3572
rect 25736 3431 25770 3443
rect 25736 3359 25770 3375
rect 25736 3287 25770 3307
rect 25736 3215 25770 3239
rect 25736 3143 25770 3171
rect 25736 3071 25770 3103
rect 25736 3001 25770 3035
rect 25736 2933 25770 2965
rect 25736 2865 25770 2893
rect 25736 2797 25770 2821
rect 25736 2729 25770 2749
rect 25736 2661 25770 2677
rect 25736 2593 25770 2605
rect 25736 2514 25770 2533
rect 25832 3503 25866 3522
rect 25832 3431 25866 3443
rect 25832 3359 25866 3375
rect 25832 3287 25866 3307
rect 25832 3215 25866 3239
rect 25832 3143 25866 3171
rect 25832 3071 25866 3103
rect 25832 3001 25866 3035
rect 25832 2933 25866 2965
rect 25832 2865 25866 2893
rect 25832 2797 25866 2821
rect 25832 2729 25866 2749
rect 25832 2661 25866 2677
rect 25832 2593 25866 2605
rect 25832 2472 25866 2533
rect 25928 3503 25962 3572
rect 25928 3431 25962 3443
rect 25928 3359 25962 3375
rect 25928 3287 25962 3307
rect 25928 3215 25962 3239
rect 25928 3143 25962 3171
rect 25928 3071 25962 3103
rect 25928 3001 25962 3035
rect 25928 2933 25962 2965
rect 25928 2865 25962 2893
rect 25928 2797 25962 2821
rect 25928 2729 25962 2749
rect 25928 2661 25962 2677
rect 25928 2593 25962 2605
rect 25928 2514 25962 2533
rect 26024 3503 26058 3522
rect 26024 3431 26058 3443
rect 26024 3359 26058 3375
rect 26024 3287 26058 3307
rect 26024 3215 26058 3239
rect 26024 3143 26058 3171
rect 26024 3071 26058 3103
rect 26024 3001 26058 3035
rect 26024 2933 26058 2965
rect 26024 2865 26058 2893
rect 26024 2797 26058 2821
rect 26024 2729 26058 2749
rect 26024 2661 26058 2677
rect 26024 2593 26058 2605
rect 26024 2472 26058 2533
rect 26120 3503 26154 3572
rect 26120 3431 26154 3443
rect 26120 3359 26154 3375
rect 26120 3287 26154 3307
rect 26120 3215 26154 3239
rect 26120 3143 26154 3171
rect 26120 3071 26154 3103
rect 26120 3001 26154 3035
rect 26120 2933 26154 2965
rect 26120 2865 26154 2893
rect 26120 2797 26154 2821
rect 26120 2729 26154 2749
rect 26120 2661 26154 2677
rect 26120 2593 26154 2605
rect 26120 2514 26154 2533
rect 26216 3503 26250 3522
rect 26216 3431 26250 3443
rect 26216 3359 26250 3375
rect 26216 3287 26250 3307
rect 26216 3215 26250 3239
rect 26216 3143 26250 3171
rect 26216 3071 26250 3103
rect 26216 3001 26250 3035
rect 26216 2933 26250 2965
rect 26216 2865 26250 2893
rect 26216 2797 26250 2821
rect 26216 2729 26250 2749
rect 26216 2661 26250 2677
rect 26216 2593 26250 2605
rect 26216 2472 26250 2533
rect 26312 3503 26346 3572
rect 26312 3431 26346 3443
rect 26312 3359 26346 3375
rect 26312 3287 26346 3307
rect 26312 3215 26346 3239
rect 26312 3143 26346 3171
rect 26312 3071 26346 3103
rect 26312 3001 26346 3035
rect 26312 2933 26346 2965
rect 26312 2865 26346 2893
rect 26312 2797 26346 2821
rect 26312 2729 26346 2749
rect 26312 2661 26346 2677
rect 26312 2593 26346 2605
rect 26312 2514 26346 2533
rect 26408 3503 26442 3522
rect 26408 3431 26442 3443
rect 26408 3359 26442 3375
rect 26408 3287 26442 3307
rect 26408 3215 26442 3239
rect 26408 3143 26442 3171
rect 26408 3071 26442 3103
rect 26408 3001 26442 3035
rect 26408 2933 26442 2965
rect 26408 2865 26442 2893
rect 26408 2797 26442 2821
rect 26408 2729 26442 2749
rect 26408 2661 26442 2677
rect 26408 2593 26442 2605
rect 26408 2472 26442 2533
rect 26504 3503 26538 3572
rect 26828 3568 28592 3602
rect 26504 3431 26538 3443
rect 26504 3359 26538 3375
rect 26504 3287 26538 3307
rect 26504 3215 26538 3239
rect 26504 3143 26538 3171
rect 26504 3071 26538 3103
rect 26504 3001 26538 3035
rect 26504 2933 26538 2965
rect 26504 2865 26538 2893
rect 26504 2797 26538 2821
rect 26504 2729 26538 2749
rect 26504 2661 26538 2677
rect 26504 2593 26538 2605
rect 26504 2514 26538 2533
rect 26732 3511 26766 3530
rect 26732 3439 26766 3451
rect 26732 3367 26766 3383
rect 26732 3295 26766 3315
rect 26732 3223 26766 3247
rect 26732 3151 26766 3179
rect 26732 3079 26766 3111
rect 26732 3009 26766 3043
rect 26732 2941 26766 2973
rect 26732 2873 26766 2901
rect 26732 2805 26766 2829
rect 26732 2737 26766 2757
rect 26732 2669 26766 2685
rect 26732 2601 26766 2613
rect 26732 2480 26766 2541
rect 26828 3511 26862 3568
rect 26828 3439 26862 3451
rect 26828 3367 26862 3383
rect 26828 3295 26862 3315
rect 26828 3223 26862 3247
rect 26828 3151 26862 3179
rect 26828 3079 26862 3111
rect 26828 3009 26862 3043
rect 26828 2941 26862 2973
rect 26828 2873 26862 2901
rect 26828 2805 26862 2829
rect 26828 2737 26862 2757
rect 26828 2669 26862 2685
rect 26828 2601 26862 2613
rect 26828 2522 26862 2541
rect 26924 3511 26958 3530
rect 26924 3439 26958 3451
rect 26924 3367 26958 3383
rect 26924 3295 26958 3315
rect 26924 3223 26958 3247
rect 26924 3151 26958 3179
rect 26924 3079 26958 3111
rect 26924 3009 26958 3043
rect 26924 2941 26958 2973
rect 26924 2873 26958 2901
rect 26924 2805 26958 2829
rect 26924 2737 26958 2757
rect 26924 2669 26958 2685
rect 26924 2601 26958 2613
rect 26924 2480 26958 2541
rect 27020 3511 27054 3568
rect 27020 3439 27054 3451
rect 27020 3367 27054 3383
rect 27020 3295 27054 3315
rect 27020 3223 27054 3247
rect 27020 3151 27054 3179
rect 27020 3079 27054 3111
rect 27020 3009 27054 3043
rect 27020 2941 27054 2973
rect 27020 2873 27054 2901
rect 27020 2805 27054 2829
rect 27020 2737 27054 2757
rect 27020 2669 27054 2685
rect 27020 2601 27054 2613
rect 27020 2522 27054 2541
rect 27116 3511 27150 3530
rect 27116 3439 27150 3451
rect 27116 3367 27150 3383
rect 27116 3295 27150 3315
rect 27116 3223 27150 3247
rect 27116 3151 27150 3179
rect 27116 3079 27150 3111
rect 27116 3009 27150 3043
rect 27116 2941 27150 2973
rect 27116 2873 27150 2901
rect 27116 2805 27150 2829
rect 27116 2737 27150 2757
rect 27116 2669 27150 2685
rect 27116 2601 27150 2613
rect 27116 2480 27150 2541
rect 27212 3511 27246 3568
rect 27212 3439 27246 3451
rect 27212 3367 27246 3383
rect 27212 3295 27246 3315
rect 27212 3223 27246 3247
rect 27212 3151 27246 3179
rect 27212 3079 27246 3111
rect 27212 3009 27246 3043
rect 27212 2941 27246 2973
rect 27212 2873 27246 2901
rect 27212 2805 27246 2829
rect 27212 2737 27246 2757
rect 27212 2669 27246 2685
rect 27212 2601 27246 2613
rect 27212 2522 27246 2541
rect 27308 3511 27342 3530
rect 27308 3439 27342 3451
rect 27308 3367 27342 3383
rect 27308 3295 27342 3315
rect 27308 3223 27342 3247
rect 27308 3151 27342 3179
rect 27308 3079 27342 3111
rect 27308 3009 27342 3043
rect 27308 2941 27342 2973
rect 27308 2873 27342 2901
rect 27308 2805 27342 2829
rect 27308 2737 27342 2757
rect 27308 2669 27342 2685
rect 27308 2601 27342 2613
rect 27308 2480 27342 2541
rect 27404 3511 27438 3568
rect 27404 3439 27438 3451
rect 27404 3367 27438 3383
rect 27404 3295 27438 3315
rect 27404 3223 27438 3247
rect 27404 3151 27438 3179
rect 27404 3079 27438 3111
rect 27404 3009 27438 3043
rect 27404 2941 27438 2973
rect 27404 2873 27438 2901
rect 27404 2805 27438 2829
rect 27404 2737 27438 2757
rect 27404 2669 27438 2685
rect 27404 2601 27438 2613
rect 27404 2522 27438 2541
rect 27500 3511 27534 3530
rect 27500 3439 27534 3451
rect 27500 3367 27534 3383
rect 27500 3295 27534 3315
rect 27500 3223 27534 3247
rect 27500 3151 27534 3179
rect 27500 3079 27534 3111
rect 27500 3009 27534 3043
rect 27500 2941 27534 2973
rect 27500 2873 27534 2901
rect 27500 2805 27534 2829
rect 27500 2737 27534 2757
rect 27500 2669 27534 2685
rect 27500 2601 27534 2613
rect 27500 2480 27534 2541
rect 27596 3511 27630 3568
rect 27596 3439 27630 3451
rect 27596 3367 27630 3383
rect 27596 3295 27630 3315
rect 27596 3223 27630 3247
rect 27596 3151 27630 3179
rect 27596 3079 27630 3111
rect 27596 3009 27630 3043
rect 27596 2941 27630 2973
rect 27596 2873 27630 2901
rect 27596 2805 27630 2829
rect 27596 2737 27630 2757
rect 27596 2669 27630 2685
rect 27596 2601 27630 2613
rect 27596 2522 27630 2541
rect 27692 3511 27726 3530
rect 27692 3439 27726 3451
rect 27692 3367 27726 3383
rect 27692 3295 27726 3315
rect 27692 3223 27726 3247
rect 27692 3151 27726 3179
rect 27692 3079 27726 3111
rect 27692 3009 27726 3043
rect 27692 2941 27726 2973
rect 27692 2873 27726 2901
rect 27692 2805 27726 2829
rect 27692 2737 27726 2757
rect 27692 2669 27726 2685
rect 27692 2601 27726 2613
rect 27692 2480 27726 2541
rect 27788 3511 27822 3568
rect 27788 3439 27822 3451
rect 27788 3367 27822 3383
rect 27788 3295 27822 3315
rect 27788 3223 27822 3247
rect 27788 3151 27822 3179
rect 27788 3079 27822 3111
rect 27788 3009 27822 3043
rect 27788 2941 27822 2973
rect 27788 2873 27822 2901
rect 27788 2805 27822 2829
rect 27788 2737 27822 2757
rect 27788 2669 27822 2685
rect 27788 2601 27822 2613
rect 27788 2522 27822 2541
rect 27884 3511 27918 3530
rect 27884 3439 27918 3451
rect 27884 3367 27918 3383
rect 27884 3295 27918 3315
rect 27884 3223 27918 3247
rect 27884 3151 27918 3179
rect 27884 3079 27918 3111
rect 27884 3009 27918 3043
rect 27884 2941 27918 2973
rect 27884 2873 27918 2901
rect 27884 2805 27918 2829
rect 27884 2737 27918 2757
rect 27884 2669 27918 2685
rect 27884 2601 27918 2613
rect 27884 2480 27918 2541
rect 27980 3511 28014 3568
rect 27980 3439 28014 3451
rect 27980 3367 28014 3383
rect 27980 3295 28014 3315
rect 27980 3223 28014 3247
rect 27980 3151 28014 3179
rect 27980 3079 28014 3111
rect 27980 3009 28014 3043
rect 27980 2941 28014 2973
rect 27980 2873 28014 2901
rect 27980 2805 28014 2829
rect 27980 2737 28014 2757
rect 27980 2669 28014 2685
rect 27980 2601 28014 2613
rect 27980 2522 28014 2541
rect 28076 3511 28110 3530
rect 28076 3439 28110 3451
rect 28076 3367 28110 3383
rect 28076 3295 28110 3315
rect 28076 3223 28110 3247
rect 28076 3151 28110 3179
rect 28076 3079 28110 3111
rect 28076 3009 28110 3043
rect 28076 2941 28110 2973
rect 28076 2873 28110 2901
rect 28076 2805 28110 2829
rect 28076 2737 28110 2757
rect 28076 2669 28110 2685
rect 28076 2601 28110 2613
rect 28076 2480 28110 2541
rect 28172 3511 28206 3568
rect 28172 3439 28206 3451
rect 28172 3367 28206 3383
rect 28172 3295 28206 3315
rect 28172 3223 28206 3247
rect 28172 3151 28206 3179
rect 28172 3079 28206 3111
rect 28172 3009 28206 3043
rect 28172 2941 28206 2973
rect 28172 2873 28206 2901
rect 28172 2805 28206 2829
rect 28172 2737 28206 2757
rect 28172 2669 28206 2685
rect 28172 2601 28206 2613
rect 28172 2522 28206 2541
rect 28268 3511 28302 3530
rect 28268 3439 28302 3451
rect 28268 3367 28302 3383
rect 28268 3295 28302 3315
rect 28268 3223 28302 3247
rect 28268 3151 28302 3179
rect 28268 3079 28302 3111
rect 28268 3009 28302 3043
rect 28268 2941 28302 2973
rect 28268 2873 28302 2901
rect 28268 2805 28302 2829
rect 28268 2737 28302 2757
rect 28268 2669 28302 2685
rect 28268 2601 28302 2613
rect 28268 2480 28302 2541
rect 28364 3511 28398 3568
rect 28364 3439 28398 3451
rect 28364 3367 28398 3383
rect 28364 3295 28398 3315
rect 28364 3223 28398 3247
rect 28364 3151 28398 3179
rect 28364 3079 28398 3111
rect 28364 3009 28398 3043
rect 28364 2941 28398 2973
rect 28364 2873 28398 2901
rect 28364 2805 28398 2829
rect 28364 2737 28398 2757
rect 28364 2669 28398 2685
rect 28364 2601 28398 2613
rect 28364 2522 28398 2541
rect 28460 3511 28494 3530
rect 28460 3439 28494 3451
rect 28460 3367 28494 3383
rect 28460 3295 28494 3315
rect 28460 3223 28494 3247
rect 28460 3151 28494 3179
rect 28460 3079 28494 3111
rect 28460 3009 28494 3043
rect 28460 2941 28494 2973
rect 28460 2873 28494 2901
rect 28460 2805 28494 2829
rect 28460 2737 28494 2757
rect 28460 2669 28494 2685
rect 28460 2601 28494 2613
rect 28460 2480 28494 2541
rect 28556 3511 28590 3568
rect 28556 3439 28590 3451
rect 28556 3367 28590 3383
rect 28556 3295 28590 3315
rect 28556 3223 28590 3247
rect 28556 3151 28590 3179
rect 28556 3079 28590 3111
rect 28556 3009 28590 3043
rect 28556 2941 28590 2973
rect 28556 2873 28590 2901
rect 28556 2805 28590 2829
rect 28556 2737 28590 2757
rect 28556 2669 28590 2685
rect 28556 2601 28590 2613
rect 28556 2522 28590 2541
rect 28652 3511 28686 3530
rect 28652 3439 28686 3451
rect 28652 3367 28686 3383
rect 28652 3295 28686 3315
rect 28652 3223 28686 3247
rect 28652 3151 28686 3179
rect 28652 3079 28686 3111
rect 28652 3009 28686 3043
rect 28652 2941 28686 2973
rect 28652 2873 28686 2901
rect 28652 2805 28686 2829
rect 28652 2737 28686 2757
rect 28652 2669 28686 2685
rect 28652 2601 28686 2613
rect 28652 2480 28686 2541
rect 25064 2468 26454 2472
rect 26732 2468 28686 2480
rect 16686 2448 22198 2460
rect 14546 2394 14579 2428
rect 14613 2394 14646 2428
rect 14096 2339 14130 2371
rect 14426 2316 14692 2350
rect 16686 2342 22166 2448
rect 23172 2446 28686 2468
rect 14096 2269 14130 2303
rect 14096 2201 14130 2233
rect 14096 2133 14130 2161
rect 14096 2065 14130 2089
rect 14096 1997 14130 2017
rect 14096 1929 14130 1945
rect 14096 1861 14130 1873
rect 14096 1736 14130 1801
rect 13712 1702 14130 1736
rect 14500 2261 14534 2280
rect 14500 2193 14534 2195
rect 14500 2157 14534 2159
rect 10966 1656 11534 1690
rect 10966 1498 11000 1656
rect 13808 1652 13842 1702
rect 14500 1638 14534 2091
rect 14658 2261 14692 2316
rect 14658 2193 14692 2195
rect 14658 2157 14692 2159
rect 16650 2334 22268 2342
rect 23172 2340 28652 2446
rect 16650 2164 16688 2334
rect 22230 2164 22268 2334
rect 16650 2156 22268 2164
rect 23138 2332 28756 2340
rect 23138 2162 23176 2332
rect 28718 2162 28756 2332
rect 23138 2154 28756 2162
rect 14658 2070 14692 2091
rect 734 1346 768 1424
rect 252 1312 1248 1346
rect -1200 1264 -1095 1298
rect -1061 1264 -1045 1298
rect -915 1264 -899 1298
rect -865 1264 -849 1298
rect -1200 1178 -1166 1264
rect 158 1253 192 1272
rect 158 1181 192 1193
rect -1588 1144 -966 1178
rect -1686 1051 -1652 1072
rect -1686 979 -1652 991
rect -1686 907 -1652 923
rect -1686 835 -1652 855
rect -1686 763 -1652 787
rect -1686 691 -1652 719
rect -1686 619 -1652 651
rect -1686 549 -1652 583
rect -1686 481 -1652 513
rect -1686 413 -1652 441
rect -1686 345 -1652 369
rect -1686 277 -1652 297
rect -1686 209 -1652 225
rect -1686 141 -1652 153
rect -1686 -18 -1652 81
rect -1588 1051 -1554 1144
rect -1588 979 -1554 991
rect -1588 907 -1554 923
rect -1588 835 -1554 855
rect -1588 763 -1554 787
rect -1588 691 -1554 719
rect -1588 619 -1554 651
rect -1588 549 -1554 583
rect -1588 481 -1554 513
rect -1588 413 -1554 441
rect -1588 345 -1554 369
rect -1588 277 -1554 297
rect -1588 209 -1554 225
rect -1588 141 -1554 153
rect -1588 60 -1554 81
rect -1490 1051 -1456 1068
rect -1490 979 -1456 991
rect -1490 907 -1456 923
rect -1490 835 -1456 855
rect -1490 763 -1456 787
rect -1490 691 -1456 719
rect -1490 619 -1456 651
rect -1490 549 -1456 583
rect -1490 481 -1456 513
rect -1490 413 -1456 441
rect -1490 345 -1456 369
rect -1490 277 -1456 297
rect -1490 209 -1456 225
rect -1490 141 -1456 153
rect -1490 -18 -1456 81
rect -1392 1051 -1358 1144
rect -1392 979 -1358 991
rect -1392 907 -1358 923
rect -1392 835 -1358 855
rect -1392 763 -1358 787
rect -1392 691 -1358 719
rect -1392 619 -1358 651
rect -1392 549 -1358 583
rect -1392 481 -1358 513
rect -1392 413 -1358 441
rect -1392 345 -1358 369
rect -1392 277 -1358 297
rect -1392 209 -1358 225
rect -1392 141 -1358 153
rect -1392 60 -1358 81
rect -1294 1051 -1260 1068
rect -1294 979 -1260 991
rect -1294 907 -1260 923
rect -1294 835 -1260 855
rect -1294 763 -1260 787
rect -1294 691 -1260 719
rect -1294 619 -1260 651
rect -1294 549 -1260 583
rect -1294 481 -1260 513
rect -1294 413 -1260 441
rect -1294 345 -1260 369
rect -1294 277 -1260 297
rect -1294 209 -1260 225
rect -1294 141 -1260 153
rect -1294 -18 -1260 81
rect -1196 1051 -1162 1144
rect -1196 979 -1162 991
rect -1196 907 -1162 923
rect -1196 835 -1162 855
rect -1196 763 -1162 787
rect -1196 691 -1162 719
rect -1196 619 -1162 651
rect -1196 549 -1162 583
rect -1196 481 -1162 513
rect -1196 413 -1162 441
rect -1196 345 -1162 369
rect -1196 277 -1162 297
rect -1196 209 -1162 225
rect -1196 141 -1162 153
rect -1196 60 -1162 81
rect -1098 1051 -1064 1068
rect -1098 979 -1064 991
rect -1098 907 -1064 923
rect -1098 835 -1064 855
rect -1098 763 -1064 787
rect -1098 691 -1064 719
rect -1098 619 -1064 651
rect -1098 549 -1064 583
rect -1098 481 -1064 513
rect -1098 413 -1064 441
rect -1098 345 -1064 369
rect -1098 277 -1064 297
rect -1098 209 -1064 225
rect -1098 141 -1064 153
rect -1098 -18 -1064 81
rect -1000 1051 -966 1144
rect 158 1109 192 1125
rect -1000 979 -966 991
rect -1000 907 -966 923
rect -1000 835 -966 855
rect -1000 763 -966 787
rect -1000 691 -966 719
rect -1000 619 -966 651
rect -1000 549 -966 583
rect -1000 481 -966 513
rect -1000 413 -966 441
rect -1000 345 -966 369
rect -1000 277 -966 297
rect -1000 209 -966 225
rect -1000 141 -966 153
rect -1000 60 -966 81
rect -902 1051 -868 1070
rect -902 979 -868 991
rect -902 907 -868 923
rect -902 835 -868 855
rect -902 763 -868 787
rect -902 691 -868 719
rect -902 619 -868 651
rect -902 549 -868 583
rect -902 481 -868 513
rect -902 413 -868 441
rect -902 345 -868 369
rect -902 277 -868 297
rect -902 209 -868 225
rect 158 1037 192 1057
rect 158 965 192 989
rect 158 893 192 921
rect 158 821 192 853
rect 158 751 192 785
rect 158 683 192 715
rect 158 615 192 643
rect 158 547 192 571
rect 158 479 192 499
rect 158 411 192 427
rect 158 343 192 355
rect 158 214 192 283
rect 254 1253 288 1312
rect 254 1181 288 1193
rect 254 1109 288 1125
rect 254 1037 288 1057
rect 254 965 288 989
rect 254 893 288 921
rect 254 821 288 853
rect 254 751 288 785
rect 254 683 288 715
rect 254 615 288 643
rect 254 547 288 571
rect 254 479 288 499
rect 254 411 288 427
rect 254 343 288 355
rect 254 264 288 283
rect 350 1253 384 1270
rect 350 1181 384 1193
rect 350 1109 384 1125
rect 350 1037 384 1057
rect 350 965 384 989
rect 350 893 384 921
rect 350 821 384 853
rect 350 751 384 785
rect 350 683 384 715
rect 350 615 384 643
rect 350 547 384 571
rect 350 479 384 499
rect 350 411 384 427
rect 350 343 384 355
rect 350 214 384 283
rect 446 1253 480 1312
rect 446 1181 480 1193
rect 446 1109 480 1125
rect 446 1037 480 1057
rect 446 965 480 989
rect 446 893 480 921
rect 446 821 480 853
rect 446 751 480 785
rect 446 683 480 715
rect 446 615 480 643
rect 446 547 480 571
rect 446 479 480 499
rect 446 411 480 427
rect 446 343 480 355
rect 446 264 480 283
rect 542 1253 576 1270
rect 542 1181 576 1193
rect 542 1109 576 1125
rect 542 1037 576 1057
rect 542 965 576 989
rect 542 893 576 921
rect 542 821 576 853
rect 542 751 576 785
rect 542 683 576 715
rect 542 615 576 643
rect 542 547 576 571
rect 542 479 576 499
rect 542 411 576 427
rect 542 343 576 355
rect 542 214 576 283
rect 638 1253 672 1312
rect 638 1181 672 1193
rect 638 1109 672 1125
rect 638 1037 672 1057
rect 638 965 672 989
rect 638 893 672 921
rect 638 821 672 853
rect 638 751 672 785
rect 638 683 672 715
rect 638 615 672 643
rect 638 547 672 571
rect 638 479 672 499
rect 638 411 672 427
rect 638 343 672 355
rect 638 264 672 283
rect 734 1253 768 1270
rect 734 1181 768 1193
rect 734 1109 768 1125
rect 734 1037 768 1057
rect 734 965 768 989
rect 734 893 768 921
rect 734 821 768 853
rect 734 751 768 785
rect 734 683 768 715
rect 734 615 768 643
rect 734 547 768 571
rect 734 479 768 499
rect 734 411 768 427
rect 734 343 768 355
rect 734 214 768 283
rect 830 1253 864 1312
rect 830 1181 864 1193
rect 830 1109 864 1125
rect 830 1037 864 1057
rect 830 965 864 989
rect 830 893 864 921
rect 830 821 864 853
rect 830 751 864 785
rect 830 683 864 715
rect 830 615 864 643
rect 830 547 864 571
rect 830 479 864 499
rect 830 411 864 427
rect 830 343 864 355
rect 830 264 864 283
rect 926 1253 960 1270
rect 926 1181 960 1193
rect 926 1109 960 1125
rect 926 1037 960 1057
rect 926 965 960 989
rect 926 893 960 921
rect 926 821 960 853
rect 926 751 960 785
rect 926 683 960 715
rect 926 615 960 643
rect 926 547 960 571
rect 926 479 960 499
rect 926 411 960 427
rect 926 343 960 355
rect 926 214 960 283
rect 1022 1253 1056 1312
rect 1022 1181 1056 1193
rect 1022 1109 1056 1125
rect 1022 1037 1056 1057
rect 1022 965 1056 989
rect 1022 893 1056 921
rect 1022 821 1056 853
rect 1022 751 1056 785
rect 1022 683 1056 715
rect 1022 615 1056 643
rect 1022 547 1056 571
rect 1022 479 1056 499
rect 1022 411 1056 427
rect 1022 343 1056 355
rect 1022 264 1056 283
rect 1118 1253 1152 1270
rect 1118 1181 1152 1193
rect 1118 1109 1152 1125
rect 1118 1037 1152 1057
rect 1118 965 1152 989
rect 1118 893 1152 921
rect 1118 821 1152 853
rect 1118 751 1152 785
rect 1118 683 1152 715
rect 1118 615 1152 643
rect 1118 547 1152 571
rect 1118 479 1152 499
rect 1118 411 1152 427
rect 1118 343 1152 355
rect 1118 214 1152 283
rect 1214 1253 1248 1312
rect 1214 1181 1248 1193
rect 1214 1109 1248 1125
rect 1214 1037 1248 1057
rect 1214 965 1248 989
rect 1214 893 1248 921
rect 1214 821 1248 853
rect 1214 751 1248 785
rect 1214 683 1248 715
rect 1214 615 1248 643
rect 1214 547 1248 571
rect 1214 479 1248 499
rect 1214 411 1248 427
rect 1214 343 1248 355
rect 1214 266 1248 283
rect 1310 1253 1344 1270
rect 1310 1181 1344 1193
rect 1310 1109 1344 1125
rect 1310 1037 1344 1057
rect 1310 965 1344 989
rect 1310 893 1344 921
rect 1310 821 1344 853
rect 1310 751 1344 785
rect 1310 683 1344 715
rect 1310 615 1344 643
rect 1310 547 1344 571
rect 1310 479 1344 499
rect 1310 411 1344 427
rect 1310 343 1344 355
rect 1310 214 1344 283
rect 158 180 1344 214
rect -902 141 -868 153
rect 140 96 156 130
rect 190 96 206 130
rect -902 -18 -868 81
rect 626 -18 722 180
rect 830 120 864 180
rect -1700 -106 722 -18
rect 626 -338 722 -106
rect 1484 30 1734 1488
rect 4574 1456 5008 1490
rect 7618 1462 8036 1496
rect 10552 1464 11000 1498
rect 14152 1604 14534 1638
rect 2400 1368 2434 1418
rect 2022 1334 3016 1368
rect 1926 1253 1960 1272
rect 1926 1181 1960 1193
rect 1926 1109 1960 1125
rect 1926 1037 1960 1057
rect 1926 965 1960 989
rect 1926 893 1960 921
rect 1926 821 1960 853
rect 1926 751 1960 785
rect 1926 683 1960 715
rect 1926 615 1960 643
rect 1926 547 1960 571
rect 1926 479 1960 499
rect 1926 411 1960 427
rect 1926 343 1960 355
rect 1926 216 1960 283
rect 2022 1253 2056 1334
rect 2022 1181 2056 1193
rect 2022 1109 2056 1125
rect 2022 1037 2056 1057
rect 2022 965 2056 989
rect 2022 893 2056 921
rect 2022 821 2056 853
rect 2022 751 2056 785
rect 2022 683 2056 715
rect 2022 615 2056 643
rect 2022 547 2056 571
rect 2022 479 2056 499
rect 2022 411 2056 427
rect 2022 343 2056 355
rect 2022 264 2056 283
rect 2118 1253 2152 1272
rect 2118 1181 2152 1193
rect 2118 1109 2152 1125
rect 2118 1037 2152 1057
rect 2118 965 2152 989
rect 2118 893 2152 921
rect 2118 821 2152 853
rect 2118 751 2152 785
rect 2118 683 2152 715
rect 2118 615 2152 643
rect 2118 547 2152 571
rect 2118 479 2152 499
rect 2118 411 2152 427
rect 2118 343 2152 355
rect 2118 216 2152 283
rect 2214 1253 2248 1334
rect 2214 1181 2248 1193
rect 2214 1109 2248 1125
rect 2214 1037 2248 1057
rect 2214 965 2248 989
rect 2214 893 2248 921
rect 2214 821 2248 853
rect 2214 751 2248 785
rect 2214 683 2248 715
rect 2214 615 2248 643
rect 2214 547 2248 571
rect 2214 479 2248 499
rect 2214 411 2248 427
rect 2214 343 2248 355
rect 2214 264 2248 283
rect 2310 1253 2344 1272
rect 2310 1181 2344 1193
rect 2310 1109 2344 1125
rect 2310 1037 2344 1057
rect 2310 965 2344 989
rect 2310 893 2344 921
rect 2310 821 2344 853
rect 2310 751 2344 785
rect 2310 683 2344 715
rect 2310 615 2344 643
rect 2310 547 2344 571
rect 2310 479 2344 499
rect 2310 411 2344 427
rect 2310 343 2344 355
rect 2310 216 2344 283
rect 2406 1253 2440 1334
rect 2406 1181 2440 1193
rect 2406 1109 2440 1125
rect 2406 1037 2440 1057
rect 2406 965 2440 989
rect 2406 893 2440 921
rect 2406 821 2440 853
rect 2406 751 2440 785
rect 2406 683 2440 715
rect 2406 615 2440 643
rect 2406 547 2440 571
rect 2406 479 2440 499
rect 2406 411 2440 427
rect 2406 343 2440 355
rect 2406 264 2440 283
rect 2502 1253 2536 1272
rect 2502 1181 2536 1193
rect 2502 1109 2536 1125
rect 2502 1037 2536 1057
rect 2502 965 2536 989
rect 2502 893 2536 921
rect 2502 821 2536 853
rect 2502 751 2536 785
rect 2502 683 2536 715
rect 2502 615 2536 643
rect 2502 547 2536 571
rect 2502 479 2536 499
rect 2502 411 2536 427
rect 2502 343 2536 355
rect 2502 216 2536 283
rect 2598 1253 2632 1334
rect 2598 1181 2632 1193
rect 2598 1109 2632 1125
rect 2598 1037 2632 1057
rect 2598 965 2632 989
rect 2598 893 2632 921
rect 2598 821 2632 853
rect 2598 751 2632 785
rect 2598 683 2632 715
rect 2598 615 2632 643
rect 2598 547 2632 571
rect 2598 479 2632 499
rect 2598 411 2632 427
rect 2598 343 2632 355
rect 2598 266 2632 283
rect 2694 1253 2728 1272
rect 2694 1181 2728 1193
rect 2694 1109 2728 1125
rect 2694 1037 2728 1057
rect 2694 965 2728 989
rect 2694 893 2728 921
rect 2694 821 2728 853
rect 2694 751 2728 785
rect 2694 683 2728 715
rect 2694 615 2728 643
rect 2694 547 2728 571
rect 2694 479 2728 499
rect 2694 411 2728 427
rect 2694 343 2728 355
rect 2694 216 2728 283
rect 2790 1253 2824 1334
rect 2790 1181 2824 1193
rect 2790 1109 2824 1125
rect 2790 1037 2824 1057
rect 2790 965 2824 989
rect 2790 893 2824 921
rect 2790 821 2824 853
rect 2790 751 2824 785
rect 2790 683 2824 715
rect 2790 615 2824 643
rect 2790 547 2824 571
rect 2790 479 2824 499
rect 2790 411 2824 427
rect 2790 343 2824 355
rect 2790 266 2824 283
rect 2886 1253 2920 1272
rect 2886 1181 2920 1193
rect 2886 1109 2920 1125
rect 2886 1037 2920 1057
rect 2886 965 2920 989
rect 2886 893 2920 921
rect 2886 821 2920 853
rect 2886 751 2920 785
rect 2886 683 2920 715
rect 2886 615 2920 643
rect 2886 547 2920 571
rect 2886 479 2920 499
rect 2886 411 2920 427
rect 2886 343 2920 355
rect 2886 216 2920 283
rect 2982 1253 3016 1334
rect 3690 1330 3724 1408
rect 3208 1296 4204 1330
rect 2982 1181 3016 1193
rect 2982 1109 3016 1125
rect 2982 1037 3016 1057
rect 2982 965 3016 989
rect 2982 893 3016 921
rect 2982 821 3016 853
rect 2982 751 3016 785
rect 2982 683 3016 715
rect 2982 615 3016 643
rect 2982 547 3016 571
rect 2982 479 3016 499
rect 2982 411 3016 427
rect 2982 343 3016 355
rect 2982 266 3016 283
rect 3114 1237 3148 1256
rect 3114 1165 3148 1177
rect 3114 1093 3148 1109
rect 3114 1021 3148 1041
rect 3114 949 3148 973
rect 3114 877 3148 905
rect 3114 805 3148 837
rect 3114 735 3148 769
rect 3114 667 3148 699
rect 3114 599 3148 627
rect 3114 531 3148 555
rect 3114 463 3148 483
rect 3114 395 3148 411
rect 3114 327 3148 339
rect 1926 182 2920 216
rect 3114 198 3148 267
rect 3210 1237 3244 1296
rect 3210 1165 3244 1177
rect 3210 1093 3244 1109
rect 3210 1021 3244 1041
rect 3210 949 3244 973
rect 3210 877 3244 905
rect 3210 805 3244 837
rect 3210 735 3244 769
rect 3210 667 3244 699
rect 3210 599 3244 627
rect 3210 531 3244 555
rect 3210 463 3244 483
rect 3210 395 3244 411
rect 3210 327 3244 339
rect 3210 248 3244 267
rect 3306 1237 3340 1254
rect 3306 1165 3340 1177
rect 3306 1093 3340 1109
rect 3306 1021 3340 1041
rect 3306 949 3340 973
rect 3306 877 3340 905
rect 3306 805 3340 837
rect 3306 735 3340 769
rect 3306 667 3340 699
rect 3306 599 3340 627
rect 3306 531 3340 555
rect 3306 463 3340 483
rect 3306 395 3340 411
rect 3306 327 3340 339
rect 3306 198 3340 267
rect 3402 1237 3436 1296
rect 3402 1165 3436 1177
rect 3402 1093 3436 1109
rect 3402 1021 3436 1041
rect 3402 949 3436 973
rect 3402 877 3436 905
rect 3402 805 3436 837
rect 3402 735 3436 769
rect 3402 667 3436 699
rect 3402 599 3436 627
rect 3402 531 3436 555
rect 3402 463 3436 483
rect 3402 395 3436 411
rect 3402 327 3436 339
rect 3402 248 3436 267
rect 3498 1237 3532 1254
rect 3498 1165 3532 1177
rect 3498 1093 3532 1109
rect 3498 1021 3532 1041
rect 3498 949 3532 973
rect 3498 877 3532 905
rect 3498 805 3532 837
rect 3498 735 3532 769
rect 3498 667 3532 699
rect 3498 599 3532 627
rect 3498 531 3532 555
rect 3498 463 3532 483
rect 3498 395 3532 411
rect 3498 327 3532 339
rect 3498 198 3532 267
rect 3594 1237 3628 1296
rect 3594 1165 3628 1177
rect 3594 1093 3628 1109
rect 3594 1021 3628 1041
rect 3594 949 3628 973
rect 3594 877 3628 905
rect 3594 805 3628 837
rect 3594 735 3628 769
rect 3594 667 3628 699
rect 3594 599 3628 627
rect 3594 531 3628 555
rect 3594 463 3628 483
rect 3594 395 3628 411
rect 3594 327 3628 339
rect 3594 248 3628 267
rect 3690 1237 3724 1254
rect 3690 1165 3724 1177
rect 3690 1093 3724 1109
rect 3690 1021 3724 1041
rect 3690 949 3724 973
rect 3690 877 3724 905
rect 3690 805 3724 837
rect 3690 735 3724 769
rect 3690 667 3724 699
rect 3690 599 3724 627
rect 3690 531 3724 555
rect 3690 463 3724 483
rect 3690 395 3724 411
rect 3690 327 3724 339
rect 3690 198 3724 267
rect 3786 1237 3820 1296
rect 3786 1165 3820 1177
rect 3786 1093 3820 1109
rect 3786 1021 3820 1041
rect 3786 949 3820 973
rect 3786 877 3820 905
rect 3786 805 3820 837
rect 3786 735 3820 769
rect 3786 667 3820 699
rect 3786 599 3820 627
rect 3786 531 3820 555
rect 3786 463 3820 483
rect 3786 395 3820 411
rect 3786 327 3820 339
rect 3786 248 3820 267
rect 3882 1237 3916 1254
rect 3882 1165 3916 1177
rect 3882 1093 3916 1109
rect 3882 1021 3916 1041
rect 3882 949 3916 973
rect 3882 877 3916 905
rect 3882 805 3916 837
rect 3882 735 3916 769
rect 3882 667 3916 699
rect 3882 599 3916 627
rect 3882 531 3916 555
rect 3882 463 3916 483
rect 3882 395 3916 411
rect 3882 327 3916 339
rect 3882 198 3916 267
rect 3978 1237 4012 1296
rect 3978 1165 4012 1177
rect 3978 1093 4012 1109
rect 3978 1021 4012 1041
rect 3978 949 4012 973
rect 3978 877 4012 905
rect 3978 805 4012 837
rect 3978 735 4012 769
rect 3978 667 4012 699
rect 3978 599 4012 627
rect 3978 531 4012 555
rect 3978 463 4012 483
rect 3978 395 4012 411
rect 3978 327 4012 339
rect 3978 248 4012 267
rect 4074 1237 4108 1254
rect 4074 1165 4108 1177
rect 4074 1093 4108 1109
rect 4074 1021 4108 1041
rect 4074 949 4108 973
rect 4074 877 4108 905
rect 4074 805 4108 837
rect 4074 735 4108 769
rect 4074 667 4108 699
rect 4074 599 4108 627
rect 4074 531 4108 555
rect 4074 463 4108 483
rect 4074 395 4108 411
rect 4074 327 4108 339
rect 4074 198 4108 267
rect 4170 1237 4204 1296
rect 4170 1165 4204 1177
rect 4170 1093 4204 1109
rect 4170 1021 4204 1041
rect 4170 949 4204 973
rect 4170 877 4204 905
rect 4170 805 4204 837
rect 4170 735 4204 769
rect 4170 667 4204 699
rect 4170 599 4204 627
rect 4170 531 4204 555
rect 4170 463 4204 483
rect 4170 395 4204 411
rect 4170 327 4204 339
rect 4170 250 4204 267
rect 4266 1237 4300 1254
rect 4266 1165 4300 1177
rect 4266 1093 4300 1109
rect 4266 1021 4300 1041
rect 4266 949 4300 973
rect 4266 877 4300 905
rect 4266 805 4300 837
rect 4266 735 4300 769
rect 4266 667 4300 699
rect 4266 599 4300 627
rect 4266 531 4300 555
rect 4266 463 4300 483
rect 4266 395 4300 411
rect 4266 327 4300 339
rect 4266 198 4300 267
rect 2494 146 2528 182
rect 3114 164 4300 198
rect 2772 96 2788 130
rect 2822 96 2838 130
rect 3096 80 3112 114
rect 3146 80 3162 114
rect 3786 104 3820 164
rect 1484 -6 1498 30
rect 1720 -6 1734 30
rect 626 -946 720 -338
rect 592 -948 720 -946
rect 1484 -948 1734 -6
rect 4574 12 4824 1456
rect 5356 1352 5390 1402
rect 4978 1318 5972 1352
rect 6720 1330 6754 1408
rect 4882 1237 4916 1256
rect 4882 1165 4916 1177
rect 4882 1093 4916 1109
rect 4882 1021 4916 1041
rect 4882 949 4916 973
rect 4882 877 4916 905
rect 4882 805 4916 837
rect 4882 735 4916 769
rect 4882 667 4916 699
rect 4882 599 4916 627
rect 4882 531 4916 555
rect 4882 463 4916 483
rect 4882 395 4916 411
rect 4882 327 4916 339
rect 4882 200 4916 267
rect 4978 1237 5012 1318
rect 4978 1165 5012 1177
rect 4978 1093 5012 1109
rect 4978 1021 5012 1041
rect 4978 949 5012 973
rect 4978 877 5012 905
rect 4978 805 5012 837
rect 4978 735 5012 769
rect 4978 667 5012 699
rect 4978 599 5012 627
rect 4978 531 5012 555
rect 4978 463 5012 483
rect 4978 395 5012 411
rect 4978 327 5012 339
rect 4978 248 5012 267
rect 5074 1237 5108 1256
rect 5074 1165 5108 1177
rect 5074 1093 5108 1109
rect 5074 1021 5108 1041
rect 5074 949 5108 973
rect 5074 877 5108 905
rect 5074 805 5108 837
rect 5074 735 5108 769
rect 5074 667 5108 699
rect 5074 599 5108 627
rect 5074 531 5108 555
rect 5074 463 5108 483
rect 5074 395 5108 411
rect 5074 327 5108 339
rect 5074 200 5108 267
rect 5170 1237 5204 1318
rect 5170 1165 5204 1177
rect 5170 1093 5204 1109
rect 5170 1021 5204 1041
rect 5170 949 5204 973
rect 5170 877 5204 905
rect 5170 805 5204 837
rect 5170 735 5204 769
rect 5170 667 5204 699
rect 5170 599 5204 627
rect 5170 531 5204 555
rect 5170 463 5204 483
rect 5170 395 5204 411
rect 5170 327 5204 339
rect 5170 248 5204 267
rect 5266 1237 5300 1256
rect 5266 1165 5300 1177
rect 5266 1093 5300 1109
rect 5266 1021 5300 1041
rect 5266 949 5300 973
rect 5266 877 5300 905
rect 5266 805 5300 837
rect 5266 735 5300 769
rect 5266 667 5300 699
rect 5266 599 5300 627
rect 5266 531 5300 555
rect 5266 463 5300 483
rect 5266 395 5300 411
rect 5266 327 5300 339
rect 5266 200 5300 267
rect 5362 1237 5396 1318
rect 5362 1165 5396 1177
rect 5362 1093 5396 1109
rect 5362 1021 5396 1041
rect 5362 949 5396 973
rect 5362 877 5396 905
rect 5362 805 5396 837
rect 5362 735 5396 769
rect 5362 667 5396 699
rect 5362 599 5396 627
rect 5362 531 5396 555
rect 5362 463 5396 483
rect 5362 395 5396 411
rect 5362 327 5396 339
rect 5362 248 5396 267
rect 5458 1237 5492 1256
rect 5458 1165 5492 1177
rect 5458 1093 5492 1109
rect 5458 1021 5492 1041
rect 5458 949 5492 973
rect 5458 877 5492 905
rect 5458 805 5492 837
rect 5458 735 5492 769
rect 5458 667 5492 699
rect 5458 599 5492 627
rect 5458 531 5492 555
rect 5458 463 5492 483
rect 5458 395 5492 411
rect 5458 327 5492 339
rect 5458 200 5492 267
rect 5554 1237 5588 1318
rect 5554 1165 5588 1177
rect 5554 1093 5588 1109
rect 5554 1021 5588 1041
rect 5554 949 5588 973
rect 5554 877 5588 905
rect 5554 805 5588 837
rect 5554 735 5588 769
rect 5554 667 5588 699
rect 5554 599 5588 627
rect 5554 531 5588 555
rect 5554 463 5588 483
rect 5554 395 5588 411
rect 5554 327 5588 339
rect 5554 250 5588 267
rect 5650 1237 5684 1256
rect 5650 1165 5684 1177
rect 5650 1093 5684 1109
rect 5650 1021 5684 1041
rect 5650 949 5684 973
rect 5650 877 5684 905
rect 5650 805 5684 837
rect 5650 735 5684 769
rect 5650 667 5684 699
rect 5650 599 5684 627
rect 5650 531 5684 555
rect 5650 463 5684 483
rect 5650 395 5684 411
rect 5650 327 5684 339
rect 5650 200 5684 267
rect 5746 1237 5780 1318
rect 5746 1165 5780 1177
rect 5746 1093 5780 1109
rect 5746 1021 5780 1041
rect 5746 949 5780 973
rect 5746 877 5780 905
rect 5746 805 5780 837
rect 5746 735 5780 769
rect 5746 667 5780 699
rect 5746 599 5780 627
rect 5746 531 5780 555
rect 5746 463 5780 483
rect 5746 395 5780 411
rect 5746 327 5780 339
rect 5746 250 5780 267
rect 5842 1237 5876 1256
rect 5842 1165 5876 1177
rect 5842 1093 5876 1109
rect 5842 1021 5876 1041
rect 5842 949 5876 973
rect 5842 877 5876 905
rect 5842 805 5876 837
rect 5842 735 5876 769
rect 5842 667 5876 699
rect 5842 599 5876 627
rect 5842 531 5876 555
rect 5842 463 5876 483
rect 5842 395 5876 411
rect 5842 327 5876 339
rect 5842 200 5876 267
rect 5938 1237 5972 1318
rect 6238 1296 7234 1330
rect 5938 1165 5972 1177
rect 5938 1093 5972 1109
rect 5938 1021 5972 1041
rect 5938 949 5972 973
rect 5938 877 5972 905
rect 5938 805 5972 837
rect 5938 735 5972 769
rect 5938 667 5972 699
rect 5938 599 5972 627
rect 5938 531 5972 555
rect 5938 463 5972 483
rect 5938 395 5972 411
rect 5938 327 5972 339
rect 5938 250 5972 267
rect 6144 1237 6178 1256
rect 6144 1165 6178 1177
rect 6144 1093 6178 1109
rect 6144 1021 6178 1041
rect 6144 949 6178 973
rect 6144 877 6178 905
rect 6144 805 6178 837
rect 6144 735 6178 769
rect 6144 667 6178 699
rect 6144 599 6178 627
rect 6144 531 6178 555
rect 6144 463 6178 483
rect 6144 395 6178 411
rect 6144 327 6178 339
rect 4882 166 5876 200
rect 6144 198 6178 267
rect 6240 1237 6274 1296
rect 6240 1165 6274 1177
rect 6240 1093 6274 1109
rect 6240 1021 6274 1041
rect 6240 949 6274 973
rect 6240 877 6274 905
rect 6240 805 6274 837
rect 6240 735 6274 769
rect 6240 667 6274 699
rect 6240 599 6274 627
rect 6240 531 6274 555
rect 6240 463 6274 483
rect 6240 395 6274 411
rect 6240 327 6274 339
rect 6240 248 6274 267
rect 6336 1237 6370 1254
rect 6336 1165 6370 1177
rect 6336 1093 6370 1109
rect 6336 1021 6370 1041
rect 6336 949 6370 973
rect 6336 877 6370 905
rect 6336 805 6370 837
rect 6336 735 6370 769
rect 6336 667 6370 699
rect 6336 599 6370 627
rect 6336 531 6370 555
rect 6336 463 6370 483
rect 6336 395 6370 411
rect 6336 327 6370 339
rect 6336 198 6370 267
rect 6432 1237 6466 1296
rect 6432 1165 6466 1177
rect 6432 1093 6466 1109
rect 6432 1021 6466 1041
rect 6432 949 6466 973
rect 6432 877 6466 905
rect 6432 805 6466 837
rect 6432 735 6466 769
rect 6432 667 6466 699
rect 6432 599 6466 627
rect 6432 531 6466 555
rect 6432 463 6466 483
rect 6432 395 6466 411
rect 6432 327 6466 339
rect 6432 248 6466 267
rect 6528 1237 6562 1254
rect 6528 1165 6562 1177
rect 6528 1093 6562 1109
rect 6528 1021 6562 1041
rect 6528 949 6562 973
rect 6528 877 6562 905
rect 6528 805 6562 837
rect 6528 735 6562 769
rect 6528 667 6562 699
rect 6528 599 6562 627
rect 6528 531 6562 555
rect 6528 463 6562 483
rect 6528 395 6562 411
rect 6528 327 6562 339
rect 6528 198 6562 267
rect 6624 1237 6658 1296
rect 6624 1165 6658 1177
rect 6624 1093 6658 1109
rect 6624 1021 6658 1041
rect 6624 949 6658 973
rect 6624 877 6658 905
rect 6624 805 6658 837
rect 6624 735 6658 769
rect 6624 667 6658 699
rect 6624 599 6658 627
rect 6624 531 6658 555
rect 6624 463 6658 483
rect 6624 395 6658 411
rect 6624 327 6658 339
rect 6624 248 6658 267
rect 6720 1237 6754 1254
rect 6720 1165 6754 1177
rect 6720 1093 6754 1109
rect 6720 1021 6754 1041
rect 6720 949 6754 973
rect 6720 877 6754 905
rect 6720 805 6754 837
rect 6720 735 6754 769
rect 6720 667 6754 699
rect 6720 599 6754 627
rect 6720 531 6754 555
rect 6720 463 6754 483
rect 6720 395 6754 411
rect 6720 327 6754 339
rect 6720 198 6754 267
rect 6816 1237 6850 1296
rect 6816 1165 6850 1177
rect 6816 1093 6850 1109
rect 6816 1021 6850 1041
rect 6816 949 6850 973
rect 6816 877 6850 905
rect 6816 805 6850 837
rect 6816 735 6850 769
rect 6816 667 6850 699
rect 6816 599 6850 627
rect 6816 531 6850 555
rect 6816 463 6850 483
rect 6816 395 6850 411
rect 6816 327 6850 339
rect 6816 248 6850 267
rect 6912 1237 6946 1254
rect 6912 1165 6946 1177
rect 6912 1093 6946 1109
rect 6912 1021 6946 1041
rect 6912 949 6946 973
rect 6912 877 6946 905
rect 6912 805 6946 837
rect 6912 735 6946 769
rect 6912 667 6946 699
rect 6912 599 6946 627
rect 6912 531 6946 555
rect 6912 463 6946 483
rect 6912 395 6946 411
rect 6912 327 6946 339
rect 6912 198 6946 267
rect 7008 1237 7042 1296
rect 7008 1165 7042 1177
rect 7008 1093 7042 1109
rect 7008 1021 7042 1041
rect 7008 949 7042 973
rect 7008 877 7042 905
rect 7008 805 7042 837
rect 7008 735 7042 769
rect 7008 667 7042 699
rect 7008 599 7042 627
rect 7008 531 7042 555
rect 7008 463 7042 483
rect 7008 395 7042 411
rect 7008 327 7042 339
rect 7008 248 7042 267
rect 7104 1237 7138 1254
rect 7104 1165 7138 1177
rect 7104 1093 7138 1109
rect 7104 1021 7138 1041
rect 7104 949 7138 973
rect 7104 877 7138 905
rect 7104 805 7138 837
rect 7104 735 7138 769
rect 7104 667 7138 699
rect 7104 599 7138 627
rect 7104 531 7138 555
rect 7104 463 7138 483
rect 7104 395 7138 411
rect 7104 327 7138 339
rect 7104 198 7138 267
rect 7200 1237 7234 1296
rect 7200 1165 7234 1177
rect 7200 1093 7234 1109
rect 7200 1021 7234 1041
rect 7200 949 7234 973
rect 7200 877 7234 905
rect 7200 805 7234 837
rect 7200 735 7234 769
rect 7200 667 7234 699
rect 7200 599 7234 627
rect 7200 531 7234 555
rect 7200 463 7234 483
rect 7200 395 7234 411
rect 7200 327 7234 339
rect 7200 250 7234 267
rect 7296 1237 7330 1254
rect 7296 1165 7330 1177
rect 7296 1093 7330 1109
rect 7296 1021 7330 1041
rect 7296 949 7330 973
rect 7296 877 7330 905
rect 7296 805 7330 837
rect 7296 735 7330 769
rect 7296 667 7330 699
rect 7296 599 7330 627
rect 7296 531 7330 555
rect 7296 463 7330 483
rect 7296 395 7330 411
rect 7296 327 7330 339
rect 7296 198 7330 267
rect 5450 130 5484 166
rect 6144 164 7330 198
rect 5728 80 5744 114
rect 5778 80 5794 114
rect 6126 80 6142 114
rect 6176 80 6192 114
rect 6816 104 6850 164
rect 4574 -24 4584 12
rect 4806 -24 4824 12
rect 4574 -948 4824 -24
rect 7618 18 7868 1462
rect 8386 1352 8420 1402
rect 8008 1318 9002 1352
rect 9808 1328 9842 1406
rect 7912 1237 7946 1256
rect 7912 1165 7946 1177
rect 7912 1093 7946 1109
rect 7912 1021 7946 1041
rect 7912 949 7946 973
rect 7912 877 7946 905
rect 7912 805 7946 837
rect 7912 735 7946 769
rect 7912 667 7946 699
rect 7912 599 7946 627
rect 7912 531 7946 555
rect 7912 463 7946 483
rect 7912 395 7946 411
rect 7912 327 7946 339
rect 7912 200 7946 267
rect 8008 1237 8042 1318
rect 8008 1165 8042 1177
rect 8008 1093 8042 1109
rect 8008 1021 8042 1041
rect 8008 949 8042 973
rect 8008 877 8042 905
rect 8008 805 8042 837
rect 8008 735 8042 769
rect 8008 667 8042 699
rect 8008 599 8042 627
rect 8008 531 8042 555
rect 8008 463 8042 483
rect 8008 395 8042 411
rect 8008 327 8042 339
rect 8008 248 8042 267
rect 8104 1237 8138 1256
rect 8104 1165 8138 1177
rect 8104 1093 8138 1109
rect 8104 1021 8138 1041
rect 8104 949 8138 973
rect 8104 877 8138 905
rect 8104 805 8138 837
rect 8104 735 8138 769
rect 8104 667 8138 699
rect 8104 599 8138 627
rect 8104 531 8138 555
rect 8104 463 8138 483
rect 8104 395 8138 411
rect 8104 327 8138 339
rect 8104 200 8138 267
rect 8200 1237 8234 1318
rect 8200 1165 8234 1177
rect 8200 1093 8234 1109
rect 8200 1021 8234 1041
rect 8200 949 8234 973
rect 8200 877 8234 905
rect 8200 805 8234 837
rect 8200 735 8234 769
rect 8200 667 8234 699
rect 8200 599 8234 627
rect 8200 531 8234 555
rect 8200 463 8234 483
rect 8200 395 8234 411
rect 8200 327 8234 339
rect 8200 248 8234 267
rect 8296 1237 8330 1256
rect 8296 1165 8330 1177
rect 8296 1093 8330 1109
rect 8296 1021 8330 1041
rect 8296 949 8330 973
rect 8296 877 8330 905
rect 8296 805 8330 837
rect 8296 735 8330 769
rect 8296 667 8330 699
rect 8296 599 8330 627
rect 8296 531 8330 555
rect 8296 463 8330 483
rect 8296 395 8330 411
rect 8296 327 8330 339
rect 8296 200 8330 267
rect 8392 1237 8426 1318
rect 8392 1165 8426 1177
rect 8392 1093 8426 1109
rect 8392 1021 8426 1041
rect 8392 949 8426 973
rect 8392 877 8426 905
rect 8392 805 8426 837
rect 8392 735 8426 769
rect 8392 667 8426 699
rect 8392 599 8426 627
rect 8392 531 8426 555
rect 8392 463 8426 483
rect 8392 395 8426 411
rect 8392 327 8426 339
rect 8392 248 8426 267
rect 8488 1237 8522 1256
rect 8488 1165 8522 1177
rect 8488 1093 8522 1109
rect 8488 1021 8522 1041
rect 8488 949 8522 973
rect 8488 877 8522 905
rect 8488 805 8522 837
rect 8488 735 8522 769
rect 8488 667 8522 699
rect 8488 599 8522 627
rect 8488 531 8522 555
rect 8488 463 8522 483
rect 8488 395 8522 411
rect 8488 327 8522 339
rect 8488 200 8522 267
rect 8584 1237 8618 1318
rect 8584 1165 8618 1177
rect 8584 1093 8618 1109
rect 8584 1021 8618 1041
rect 8584 949 8618 973
rect 8584 877 8618 905
rect 8584 805 8618 837
rect 8584 735 8618 769
rect 8584 667 8618 699
rect 8584 599 8618 627
rect 8584 531 8618 555
rect 8584 463 8618 483
rect 8584 395 8618 411
rect 8584 327 8618 339
rect 8584 250 8618 267
rect 8680 1237 8714 1256
rect 8680 1165 8714 1177
rect 8680 1093 8714 1109
rect 8680 1021 8714 1041
rect 8680 949 8714 973
rect 8680 877 8714 905
rect 8680 805 8714 837
rect 8680 735 8714 769
rect 8680 667 8714 699
rect 8680 599 8714 627
rect 8680 531 8714 555
rect 8680 463 8714 483
rect 8680 395 8714 411
rect 8680 327 8714 339
rect 8680 200 8714 267
rect 8776 1237 8810 1318
rect 8776 1165 8810 1177
rect 8776 1093 8810 1109
rect 8776 1021 8810 1041
rect 8776 949 8810 973
rect 8776 877 8810 905
rect 8776 805 8810 837
rect 8776 735 8810 769
rect 8776 667 8810 699
rect 8776 599 8810 627
rect 8776 531 8810 555
rect 8776 463 8810 483
rect 8776 395 8810 411
rect 8776 327 8810 339
rect 8776 250 8810 267
rect 8872 1237 8906 1256
rect 8872 1165 8906 1177
rect 8872 1093 8906 1109
rect 8872 1021 8906 1041
rect 8872 949 8906 973
rect 8872 877 8906 905
rect 8872 805 8906 837
rect 8872 735 8906 769
rect 8872 667 8906 699
rect 8872 599 8906 627
rect 8872 531 8906 555
rect 8872 463 8906 483
rect 8872 395 8906 411
rect 8872 327 8906 339
rect 8872 200 8906 267
rect 8968 1237 9002 1318
rect 9326 1294 10322 1328
rect 8968 1165 9002 1177
rect 8968 1093 9002 1109
rect 8968 1021 9002 1041
rect 8968 949 9002 973
rect 8968 877 9002 905
rect 8968 805 9002 837
rect 8968 735 9002 769
rect 8968 667 9002 699
rect 8968 599 9002 627
rect 8968 531 9002 555
rect 8968 463 9002 483
rect 8968 395 9002 411
rect 8968 327 9002 339
rect 8968 250 9002 267
rect 9232 1235 9266 1254
rect 9232 1163 9266 1175
rect 9232 1091 9266 1107
rect 9232 1019 9266 1039
rect 9232 947 9266 971
rect 9232 875 9266 903
rect 9232 803 9266 835
rect 9232 733 9266 767
rect 9232 665 9266 697
rect 9232 597 9266 625
rect 9232 529 9266 553
rect 9232 461 9266 481
rect 9232 393 9266 409
rect 9232 325 9266 337
rect 7912 166 8906 200
rect 9232 196 9266 265
rect 9328 1235 9362 1294
rect 9328 1163 9362 1175
rect 9328 1091 9362 1107
rect 9328 1019 9362 1039
rect 9328 947 9362 971
rect 9328 875 9362 903
rect 9328 803 9362 835
rect 9328 733 9362 767
rect 9328 665 9362 697
rect 9328 597 9362 625
rect 9328 529 9362 553
rect 9328 461 9362 481
rect 9328 393 9362 409
rect 9328 325 9362 337
rect 9328 246 9362 265
rect 9424 1235 9458 1252
rect 9424 1163 9458 1175
rect 9424 1091 9458 1107
rect 9424 1019 9458 1039
rect 9424 947 9458 971
rect 9424 875 9458 903
rect 9424 803 9458 835
rect 9424 733 9458 767
rect 9424 665 9458 697
rect 9424 597 9458 625
rect 9424 529 9458 553
rect 9424 461 9458 481
rect 9424 393 9458 409
rect 9424 325 9458 337
rect 9424 196 9458 265
rect 9520 1235 9554 1294
rect 9520 1163 9554 1175
rect 9520 1091 9554 1107
rect 9520 1019 9554 1039
rect 9520 947 9554 971
rect 9520 875 9554 903
rect 9520 803 9554 835
rect 9520 733 9554 767
rect 9520 665 9554 697
rect 9520 597 9554 625
rect 9520 529 9554 553
rect 9520 461 9554 481
rect 9520 393 9554 409
rect 9520 325 9554 337
rect 9520 246 9554 265
rect 9616 1235 9650 1252
rect 9616 1163 9650 1175
rect 9616 1091 9650 1107
rect 9616 1019 9650 1039
rect 9616 947 9650 971
rect 9616 875 9650 903
rect 9616 803 9650 835
rect 9616 733 9650 767
rect 9616 665 9650 697
rect 9616 597 9650 625
rect 9616 529 9650 553
rect 9616 461 9650 481
rect 9616 393 9650 409
rect 9616 325 9650 337
rect 9616 196 9650 265
rect 9712 1235 9746 1294
rect 9712 1163 9746 1175
rect 9712 1091 9746 1107
rect 9712 1019 9746 1039
rect 9712 947 9746 971
rect 9712 875 9746 903
rect 9712 803 9746 835
rect 9712 733 9746 767
rect 9712 665 9746 697
rect 9712 597 9746 625
rect 9712 529 9746 553
rect 9712 461 9746 481
rect 9712 393 9746 409
rect 9712 325 9746 337
rect 9712 246 9746 265
rect 9808 1235 9842 1252
rect 9808 1163 9842 1175
rect 9808 1091 9842 1107
rect 9808 1019 9842 1039
rect 9808 947 9842 971
rect 9808 875 9842 903
rect 9808 803 9842 835
rect 9808 733 9842 767
rect 9808 665 9842 697
rect 9808 597 9842 625
rect 9808 529 9842 553
rect 9808 461 9842 481
rect 9808 393 9842 409
rect 9808 325 9842 337
rect 9808 196 9842 265
rect 9904 1235 9938 1294
rect 9904 1163 9938 1175
rect 9904 1091 9938 1107
rect 9904 1019 9938 1039
rect 9904 947 9938 971
rect 9904 875 9938 903
rect 9904 803 9938 835
rect 9904 733 9938 767
rect 9904 665 9938 697
rect 9904 597 9938 625
rect 9904 529 9938 553
rect 9904 461 9938 481
rect 9904 393 9938 409
rect 9904 325 9938 337
rect 9904 246 9938 265
rect 10000 1235 10034 1252
rect 10000 1163 10034 1175
rect 10000 1091 10034 1107
rect 10000 1019 10034 1039
rect 10000 947 10034 971
rect 10000 875 10034 903
rect 10000 803 10034 835
rect 10000 733 10034 767
rect 10000 665 10034 697
rect 10000 597 10034 625
rect 10000 529 10034 553
rect 10000 461 10034 481
rect 10000 393 10034 409
rect 10000 325 10034 337
rect 10000 196 10034 265
rect 10096 1235 10130 1294
rect 10096 1163 10130 1175
rect 10096 1091 10130 1107
rect 10096 1019 10130 1039
rect 10096 947 10130 971
rect 10096 875 10130 903
rect 10096 803 10130 835
rect 10096 733 10130 767
rect 10096 665 10130 697
rect 10096 597 10130 625
rect 10096 529 10130 553
rect 10096 461 10130 481
rect 10096 393 10130 409
rect 10096 325 10130 337
rect 10096 246 10130 265
rect 10192 1235 10226 1252
rect 10192 1163 10226 1175
rect 10192 1091 10226 1107
rect 10192 1019 10226 1039
rect 10192 947 10226 971
rect 10192 875 10226 903
rect 10192 803 10226 835
rect 10192 733 10226 767
rect 10192 665 10226 697
rect 10192 597 10226 625
rect 10192 529 10226 553
rect 10192 461 10226 481
rect 10192 393 10226 409
rect 10192 325 10226 337
rect 10192 196 10226 265
rect 10288 1235 10322 1294
rect 10288 1163 10322 1175
rect 10288 1091 10322 1107
rect 10288 1019 10322 1039
rect 10288 947 10322 971
rect 10288 875 10322 903
rect 10288 803 10322 835
rect 10288 733 10322 767
rect 10288 665 10322 697
rect 10288 597 10322 625
rect 10288 529 10322 553
rect 10288 461 10322 481
rect 10288 393 10322 409
rect 10288 325 10322 337
rect 10288 248 10322 265
rect 10384 1235 10418 1252
rect 10384 1163 10418 1175
rect 10384 1091 10418 1107
rect 10384 1019 10418 1039
rect 10384 947 10418 971
rect 10384 875 10418 903
rect 10384 803 10418 835
rect 10384 733 10418 767
rect 10384 665 10418 697
rect 10384 597 10418 625
rect 10384 529 10418 553
rect 10384 461 10418 481
rect 10384 393 10418 409
rect 10384 325 10418 337
rect 10384 196 10418 265
rect 8480 130 8514 166
rect 9232 162 10418 196
rect 8758 80 8774 114
rect 8808 80 8824 114
rect 9214 78 9230 112
rect 9264 78 9280 112
rect 9904 102 9938 162
rect 7618 -16 7632 18
rect 7854 -16 7868 18
rect 7618 -948 7868 -16
rect 10552 12 10802 1464
rect 14152 1448 14186 1604
rect 15450 1458 15466 1492
rect 15500 1458 15516 1492
rect 13848 1414 14186 1448
rect 11474 1350 11508 1400
rect 11096 1316 12090 1350
rect 11000 1235 11034 1254
rect 11000 1163 11034 1175
rect 11000 1091 11034 1107
rect 11000 1019 11034 1039
rect 11000 947 11034 971
rect 11000 875 11034 903
rect 11000 803 11034 835
rect 11000 733 11034 767
rect 11000 665 11034 697
rect 11000 597 11034 625
rect 11000 529 11034 553
rect 11000 461 11034 481
rect 11000 393 11034 409
rect 11000 325 11034 337
rect 11000 198 11034 265
rect 11096 1235 11130 1316
rect 11096 1163 11130 1175
rect 11096 1091 11130 1107
rect 11096 1019 11130 1039
rect 11096 947 11130 971
rect 11096 875 11130 903
rect 11096 803 11130 835
rect 11096 733 11130 767
rect 11096 665 11130 697
rect 11096 597 11130 625
rect 11096 529 11130 553
rect 11096 461 11130 481
rect 11096 393 11130 409
rect 11096 325 11130 337
rect 11096 246 11130 265
rect 11192 1235 11226 1254
rect 11192 1163 11226 1175
rect 11192 1091 11226 1107
rect 11192 1019 11226 1039
rect 11192 947 11226 971
rect 11192 875 11226 903
rect 11192 803 11226 835
rect 11192 733 11226 767
rect 11192 665 11226 697
rect 11192 597 11226 625
rect 11192 529 11226 553
rect 11192 461 11226 481
rect 11192 393 11226 409
rect 11192 325 11226 337
rect 11192 198 11226 265
rect 11288 1235 11322 1316
rect 11288 1163 11322 1175
rect 11288 1091 11322 1107
rect 11288 1019 11322 1039
rect 11288 947 11322 971
rect 11288 875 11322 903
rect 11288 803 11322 835
rect 11288 733 11322 767
rect 11288 665 11322 697
rect 11288 597 11322 625
rect 11288 529 11322 553
rect 11288 461 11322 481
rect 11288 393 11322 409
rect 11288 325 11322 337
rect 11288 246 11322 265
rect 11384 1235 11418 1254
rect 11384 1163 11418 1175
rect 11384 1091 11418 1107
rect 11384 1019 11418 1039
rect 11384 947 11418 971
rect 11384 875 11418 903
rect 11384 803 11418 835
rect 11384 733 11418 767
rect 11384 665 11418 697
rect 11384 597 11418 625
rect 11384 529 11418 553
rect 11384 461 11418 481
rect 11384 393 11418 409
rect 11384 325 11418 337
rect 11384 198 11418 265
rect 11480 1235 11514 1316
rect 11480 1163 11514 1175
rect 11480 1091 11514 1107
rect 11480 1019 11514 1039
rect 11480 947 11514 971
rect 11480 875 11514 903
rect 11480 803 11514 835
rect 11480 733 11514 767
rect 11480 665 11514 697
rect 11480 597 11514 625
rect 11480 529 11514 553
rect 11480 461 11514 481
rect 11480 393 11514 409
rect 11480 325 11514 337
rect 11480 246 11514 265
rect 11576 1235 11610 1254
rect 11576 1163 11610 1175
rect 11576 1091 11610 1107
rect 11576 1019 11610 1039
rect 11576 947 11610 971
rect 11576 875 11610 903
rect 11576 803 11610 835
rect 11576 733 11610 767
rect 11576 665 11610 697
rect 11576 597 11610 625
rect 11576 529 11610 553
rect 11576 461 11610 481
rect 11576 393 11610 409
rect 11576 325 11610 337
rect 11576 198 11610 265
rect 11672 1235 11706 1316
rect 11672 1163 11706 1175
rect 11672 1091 11706 1107
rect 11672 1019 11706 1039
rect 11672 947 11706 971
rect 11672 875 11706 903
rect 11672 803 11706 835
rect 11672 733 11706 767
rect 11672 665 11706 697
rect 11672 597 11706 625
rect 11672 529 11706 553
rect 11672 461 11706 481
rect 11672 393 11706 409
rect 11672 325 11706 337
rect 11672 248 11706 265
rect 11768 1235 11802 1254
rect 11768 1163 11802 1175
rect 11768 1091 11802 1107
rect 11768 1019 11802 1039
rect 11768 947 11802 971
rect 11768 875 11802 903
rect 11768 803 11802 835
rect 11768 733 11802 767
rect 11768 665 11802 697
rect 11768 597 11802 625
rect 11768 529 11802 553
rect 11768 461 11802 481
rect 11768 393 11802 409
rect 11768 325 11802 337
rect 11768 198 11802 265
rect 11864 1235 11898 1316
rect 11864 1163 11898 1175
rect 11864 1091 11898 1107
rect 11864 1019 11898 1039
rect 11864 947 11898 971
rect 11864 875 11898 903
rect 11864 803 11898 835
rect 11864 733 11898 767
rect 11864 665 11898 697
rect 11864 597 11898 625
rect 11864 529 11898 553
rect 11864 461 11898 481
rect 11864 393 11898 409
rect 11864 325 11898 337
rect 11864 248 11898 265
rect 11960 1235 11994 1254
rect 11960 1163 11994 1175
rect 11960 1091 11994 1107
rect 11960 1019 11994 1039
rect 11960 947 11994 971
rect 11960 875 11994 903
rect 11960 803 11994 835
rect 11960 733 11994 767
rect 11960 665 11994 697
rect 11960 597 11994 625
rect 11960 529 11994 553
rect 11960 461 11994 481
rect 11960 393 11994 409
rect 11960 325 11994 337
rect 11960 198 11994 265
rect 12056 1235 12090 1316
rect 12964 1302 12998 1380
rect 12482 1268 13478 1302
rect 12056 1163 12090 1175
rect 12056 1091 12090 1107
rect 12056 1019 12090 1039
rect 12056 947 12090 971
rect 12056 875 12090 903
rect 12056 803 12090 835
rect 12056 733 12090 767
rect 12056 665 12090 697
rect 12056 597 12090 625
rect 12056 529 12090 553
rect 12056 461 12090 481
rect 12056 393 12090 409
rect 12056 325 12090 337
rect 12056 248 12090 265
rect 12388 1209 12422 1228
rect 12388 1137 12422 1149
rect 12388 1065 12422 1081
rect 12388 993 12422 1013
rect 12388 921 12422 945
rect 12388 849 12422 877
rect 12388 777 12422 809
rect 12388 707 12422 741
rect 12388 639 12422 671
rect 12388 571 12422 599
rect 12388 503 12422 527
rect 12388 435 12422 455
rect 12388 367 12422 383
rect 12388 299 12422 311
rect 11000 164 11994 198
rect 12388 170 12422 239
rect 12484 1209 12518 1268
rect 12484 1137 12518 1149
rect 12484 1065 12518 1081
rect 12484 993 12518 1013
rect 12484 921 12518 945
rect 12484 849 12518 877
rect 12484 777 12518 809
rect 12484 707 12518 741
rect 12484 639 12518 671
rect 12484 571 12518 599
rect 12484 503 12518 527
rect 12484 435 12518 455
rect 12484 367 12518 383
rect 12484 299 12518 311
rect 12484 220 12518 239
rect 12580 1209 12614 1226
rect 12580 1137 12614 1149
rect 12580 1065 12614 1081
rect 12580 993 12614 1013
rect 12580 921 12614 945
rect 12580 849 12614 877
rect 12580 777 12614 809
rect 12580 707 12614 741
rect 12580 639 12614 671
rect 12580 571 12614 599
rect 12580 503 12614 527
rect 12580 435 12614 455
rect 12580 367 12614 383
rect 12580 299 12614 311
rect 12580 170 12614 239
rect 12676 1209 12710 1268
rect 12676 1137 12710 1149
rect 12676 1065 12710 1081
rect 12676 993 12710 1013
rect 12676 921 12710 945
rect 12676 849 12710 877
rect 12676 777 12710 809
rect 12676 707 12710 741
rect 12676 639 12710 671
rect 12676 571 12710 599
rect 12676 503 12710 527
rect 12676 435 12710 455
rect 12676 367 12710 383
rect 12676 299 12710 311
rect 12676 220 12710 239
rect 12772 1209 12806 1226
rect 12772 1137 12806 1149
rect 12772 1065 12806 1081
rect 12772 993 12806 1013
rect 12772 921 12806 945
rect 12772 849 12806 877
rect 12772 777 12806 809
rect 12772 707 12806 741
rect 12772 639 12806 671
rect 12772 571 12806 599
rect 12772 503 12806 527
rect 12772 435 12806 455
rect 12772 367 12806 383
rect 12772 299 12806 311
rect 12772 170 12806 239
rect 12868 1209 12902 1268
rect 12868 1137 12902 1149
rect 12868 1065 12902 1081
rect 12868 993 12902 1013
rect 12868 921 12902 945
rect 12868 849 12902 877
rect 12868 777 12902 809
rect 12868 707 12902 741
rect 12868 639 12902 671
rect 12868 571 12902 599
rect 12868 503 12902 527
rect 12868 435 12902 455
rect 12868 367 12902 383
rect 12868 299 12902 311
rect 12868 220 12902 239
rect 12964 1209 12998 1226
rect 12964 1137 12998 1149
rect 12964 1065 12998 1081
rect 12964 993 12998 1013
rect 12964 921 12998 945
rect 12964 849 12998 877
rect 12964 777 12998 809
rect 12964 707 12998 741
rect 12964 639 12998 671
rect 12964 571 12998 599
rect 12964 503 12998 527
rect 12964 435 12998 455
rect 12964 367 12998 383
rect 12964 299 12998 311
rect 12964 170 12998 239
rect 13060 1209 13094 1268
rect 13060 1137 13094 1149
rect 13060 1065 13094 1081
rect 13060 993 13094 1013
rect 13060 921 13094 945
rect 13060 849 13094 877
rect 13060 777 13094 809
rect 13060 707 13094 741
rect 13060 639 13094 671
rect 13060 571 13094 599
rect 13060 503 13094 527
rect 13060 435 13094 455
rect 13060 367 13094 383
rect 13060 299 13094 311
rect 13060 220 13094 239
rect 13156 1209 13190 1226
rect 13156 1137 13190 1149
rect 13156 1065 13190 1081
rect 13156 993 13190 1013
rect 13156 921 13190 945
rect 13156 849 13190 877
rect 13156 777 13190 809
rect 13156 707 13190 741
rect 13156 639 13190 671
rect 13156 571 13190 599
rect 13156 503 13190 527
rect 13156 435 13190 455
rect 13156 367 13190 383
rect 13156 299 13190 311
rect 13156 170 13190 239
rect 13252 1209 13286 1268
rect 13252 1137 13286 1149
rect 13252 1065 13286 1081
rect 13252 993 13286 1013
rect 13252 921 13286 945
rect 13252 849 13286 877
rect 13252 777 13286 809
rect 13252 707 13286 741
rect 13252 639 13286 671
rect 13252 571 13286 599
rect 13252 503 13286 527
rect 13252 435 13286 455
rect 13252 367 13286 383
rect 13252 299 13286 311
rect 13252 220 13286 239
rect 13348 1209 13382 1226
rect 13348 1137 13382 1149
rect 13348 1065 13382 1081
rect 13348 993 13382 1013
rect 13348 921 13382 945
rect 13348 849 13382 877
rect 13348 777 13382 809
rect 13348 707 13382 741
rect 13348 639 13382 671
rect 13348 571 13382 599
rect 13348 503 13382 527
rect 13348 435 13382 455
rect 13348 367 13382 383
rect 13348 299 13382 311
rect 13348 170 13382 239
rect 13444 1209 13478 1268
rect 13444 1137 13478 1149
rect 13444 1065 13478 1081
rect 13444 993 13478 1013
rect 13444 921 13478 945
rect 13444 849 13478 877
rect 13444 777 13478 809
rect 13444 707 13478 741
rect 13444 639 13478 671
rect 13444 571 13478 599
rect 13444 503 13478 527
rect 13444 435 13478 455
rect 13444 367 13478 383
rect 13444 299 13478 311
rect 13444 222 13478 239
rect 13540 1209 13574 1226
rect 13540 1137 13574 1149
rect 13540 1065 13574 1081
rect 13540 993 13574 1013
rect 13540 921 13574 945
rect 13540 849 13574 877
rect 13540 777 13574 809
rect 13540 707 13574 741
rect 13540 639 13574 671
rect 13540 571 13574 599
rect 13540 503 13574 527
rect 13540 435 13574 455
rect 13540 367 13574 383
rect 13540 299 13574 311
rect 13540 170 13574 239
rect 11568 128 11602 164
rect 12388 136 13574 170
rect 11846 78 11862 112
rect 11896 78 11912 112
rect 12370 52 12386 86
rect 12420 52 12436 86
rect 13060 76 13094 136
rect 10552 -24 10562 12
rect 10796 -24 10802 12
rect 10552 -948 10802 -24
rect 13848 -14 14098 1414
rect 14630 1324 14664 1374
rect 14252 1290 15246 1324
rect 14156 1209 14190 1228
rect 14156 1137 14190 1149
rect 14156 1065 14190 1081
rect 14156 993 14190 1013
rect 14156 921 14190 945
rect 14156 849 14190 877
rect 14156 777 14190 809
rect 14156 707 14190 741
rect 14156 639 14190 671
rect 14156 571 14190 599
rect 14156 503 14190 527
rect 14156 435 14190 455
rect 14156 367 14190 383
rect 14156 299 14190 311
rect 14156 172 14190 239
rect 14252 1209 14286 1290
rect 14252 1137 14286 1149
rect 14252 1065 14286 1081
rect 14252 993 14286 1013
rect 14252 921 14286 945
rect 14252 849 14286 877
rect 14252 777 14286 809
rect 14252 707 14286 741
rect 14252 639 14286 671
rect 14252 571 14286 599
rect 14252 503 14286 527
rect 14252 435 14286 455
rect 14252 367 14286 383
rect 14252 299 14286 311
rect 14252 220 14286 239
rect 14348 1209 14382 1228
rect 14348 1137 14382 1149
rect 14348 1065 14382 1081
rect 14348 993 14382 1013
rect 14348 921 14382 945
rect 14348 849 14382 877
rect 14348 777 14382 809
rect 14348 707 14382 741
rect 14348 639 14382 671
rect 14348 571 14382 599
rect 14348 503 14382 527
rect 14348 435 14382 455
rect 14348 367 14382 383
rect 14348 299 14382 311
rect 14348 172 14382 239
rect 14444 1209 14478 1290
rect 14444 1137 14478 1149
rect 14444 1065 14478 1081
rect 14444 993 14478 1013
rect 14444 921 14478 945
rect 14444 849 14478 877
rect 14444 777 14478 809
rect 14444 707 14478 741
rect 14444 639 14478 671
rect 14444 571 14478 599
rect 14444 503 14478 527
rect 14444 435 14478 455
rect 14444 367 14478 383
rect 14444 299 14478 311
rect 14444 220 14478 239
rect 14540 1209 14574 1228
rect 14540 1137 14574 1149
rect 14540 1065 14574 1081
rect 14540 993 14574 1013
rect 14540 921 14574 945
rect 14540 849 14574 877
rect 14540 777 14574 809
rect 14540 707 14574 741
rect 14540 639 14574 671
rect 14540 571 14574 599
rect 14540 503 14574 527
rect 14540 435 14574 455
rect 14540 367 14574 383
rect 14540 299 14574 311
rect 14540 172 14574 239
rect 14636 1209 14670 1290
rect 14636 1137 14670 1149
rect 14636 1065 14670 1081
rect 14636 993 14670 1013
rect 14636 921 14670 945
rect 14636 849 14670 877
rect 14636 777 14670 809
rect 14636 707 14670 741
rect 14636 639 14670 671
rect 14636 571 14670 599
rect 14636 503 14670 527
rect 14636 435 14670 455
rect 14636 367 14670 383
rect 14636 299 14670 311
rect 14636 220 14670 239
rect 14732 1209 14766 1228
rect 14732 1137 14766 1149
rect 14732 1065 14766 1081
rect 14732 993 14766 1013
rect 14732 921 14766 945
rect 14732 849 14766 877
rect 14732 777 14766 809
rect 14732 707 14766 741
rect 14732 639 14766 671
rect 14732 571 14766 599
rect 14732 503 14766 527
rect 14732 435 14766 455
rect 14732 367 14766 383
rect 14732 299 14766 311
rect 14732 172 14766 239
rect 14828 1209 14862 1290
rect 14828 1137 14862 1149
rect 14828 1065 14862 1081
rect 14828 993 14862 1013
rect 14828 921 14862 945
rect 14828 849 14862 877
rect 14828 777 14862 809
rect 14828 707 14862 741
rect 14828 639 14862 671
rect 14828 571 14862 599
rect 14828 503 14862 527
rect 14828 435 14862 455
rect 14828 367 14862 383
rect 14828 299 14862 311
rect 14828 222 14862 239
rect 14924 1209 14958 1228
rect 14924 1137 14958 1149
rect 14924 1065 14958 1081
rect 14924 993 14958 1013
rect 14924 921 14958 945
rect 14924 849 14958 877
rect 14924 777 14958 809
rect 14924 707 14958 741
rect 14924 639 14958 671
rect 14924 571 14958 599
rect 14924 503 14958 527
rect 14924 435 14958 455
rect 14924 367 14958 383
rect 14924 299 14958 311
rect 14924 172 14958 239
rect 15020 1209 15054 1290
rect 15020 1137 15054 1149
rect 15020 1065 15054 1081
rect 15020 993 15054 1013
rect 15020 921 15054 945
rect 15020 849 15054 877
rect 15020 777 15054 809
rect 15020 707 15054 741
rect 15020 639 15054 671
rect 15020 571 15054 599
rect 15020 503 15054 527
rect 15020 435 15054 455
rect 15020 367 15054 383
rect 15020 299 15054 311
rect 15020 222 15054 239
rect 15116 1209 15150 1228
rect 15116 1137 15150 1149
rect 15116 1065 15150 1081
rect 15116 993 15150 1013
rect 15116 921 15150 945
rect 15116 849 15150 877
rect 15116 777 15150 809
rect 15116 707 15150 741
rect 15116 639 15150 671
rect 15116 571 15150 599
rect 15116 503 15150 527
rect 15116 435 15150 455
rect 15116 367 15150 383
rect 15116 299 15150 311
rect 15116 172 15150 239
rect 15212 1209 15246 1290
rect 15212 1137 15246 1149
rect 15212 1065 15246 1081
rect 15212 993 15246 1013
rect 15212 921 15246 945
rect 15212 849 15246 877
rect 15212 777 15246 809
rect 15212 707 15246 741
rect 15212 639 15246 671
rect 15212 571 15246 599
rect 15212 503 15246 527
rect 15212 435 15246 455
rect 15212 367 15246 383
rect 15212 299 15246 311
rect 15212 222 15246 239
rect 15422 1261 15456 1336
rect 15422 1193 15456 1223
rect 15422 1125 15456 1151
rect 15422 1057 15456 1079
rect 15422 989 15456 1007
rect 15422 921 15456 935
rect 15422 853 15456 863
rect 15422 785 15456 791
rect 15422 717 15456 719
rect 15422 681 15456 683
rect 15422 609 15456 615
rect 15422 537 15456 547
rect 15422 465 15456 479
rect 15422 393 15456 411
rect 15422 321 15456 343
rect 15422 249 15456 275
rect 14156 138 15150 172
rect 15422 177 15456 207
rect 14724 102 14758 138
rect 15422 96 15456 139
rect 15510 1261 15544 1304
rect 15510 1193 15544 1223
rect 15510 1125 15544 1151
rect 15510 1057 15544 1079
rect 15510 989 15544 1007
rect 15510 921 15544 935
rect 15510 853 15544 863
rect 15510 785 15544 791
rect 15510 717 15544 719
rect 15510 681 15544 683
rect 15510 609 15544 615
rect 15510 537 15544 547
rect 15510 465 15544 479
rect 15510 393 15544 411
rect 15510 321 15544 343
rect 15510 249 15544 275
rect 15510 177 15544 207
rect 15002 52 15018 86
rect 15052 52 15068 86
rect 15510 52 15544 139
rect 15510 16 15544 18
rect 13848 -50 13856 -14
rect 14090 -50 14098 -14
rect 13848 -948 14098 -50
rect 258 -963 15772 -948
rect 258 -1269 280 -963
rect 15750 -1269 15772 -963
rect 258 -1284 15772 -1269
rect 2238 -1465 2478 -1284
rect 2238 -1643 2269 -1465
rect 2447 -1643 2478 -1465
rect 2238 -1648 2478 -1643
rect 4238 -1465 4478 -1284
rect 4238 -1643 4269 -1465
rect 4447 -1643 4478 -1465
rect 4238 -1648 4478 -1643
rect 6238 -1465 6478 -1284
rect 6238 -1643 6269 -1465
rect 6447 -1643 6478 -1465
rect 6238 -1648 6478 -1643
rect 8462 -1482 8702 -1284
rect 8462 -1660 8493 -1482
rect 8671 -1660 8702 -1482
rect 10238 -1465 10478 -1284
rect 10238 -1643 10269 -1465
rect 10447 -1643 10478 -1465
rect 10238 -1648 10478 -1643
rect 12238 -1465 12478 -1284
rect 12238 -1643 12269 -1465
rect 12447 -1643 12478 -1465
rect 12238 -1648 12478 -1643
rect 14238 -1465 14478 -1284
rect 14238 -1643 14269 -1465
rect 14447 -1643 14478 -1465
rect 14238 -1648 14478 -1643
rect 8462 -1664 8702 -1660
<< viali >>
rect -344 8844 -166 9022
rect 1656 8844 1834 9022
rect 3656 8844 3834 9022
rect 5656 8844 5834 9022
rect 7656 8844 7834 9022
rect 9656 8844 9834 9022
rect 11656 8844 11834 9022
rect 13656 8844 13834 9022
rect 15454 8879 15632 9057
rect -1251 7921 -857 8099
rect 15491 7928 15741 8106
rect 764 6858 798 6892
rect 288 6773 322 6807
rect 1694 6792 1888 6896
rect 3720 6842 3754 6876
rect 2440 6754 2474 6788
rect 2728 6769 2762 6803
rect 3244 6757 3278 6791
rect 4552 6776 4746 6880
rect 6750 6842 6784 6876
rect 5396 6738 5430 6772
rect 5684 6753 5718 6787
rect 6274 6757 6308 6791
rect 194 6565 228 6591
rect 194 6557 228 6565
rect 194 6497 228 6519
rect 194 6485 228 6497
rect 194 6429 228 6447
rect 194 6413 228 6429
rect 194 6361 228 6375
rect 194 6341 228 6361
rect 194 6293 228 6303
rect 194 6269 228 6293
rect 194 6225 228 6231
rect 194 6197 228 6225
rect 194 6157 228 6159
rect 194 6125 228 6157
rect 194 6055 228 6087
rect 194 6053 228 6055
rect -1652 5895 -1618 5921
rect -1652 5887 -1618 5895
rect -1652 5827 -1618 5849
rect -1652 5815 -1618 5827
rect -1652 5759 -1618 5777
rect -1652 5743 -1618 5759
rect -1652 5691 -1618 5705
rect -1652 5671 -1618 5691
rect -1652 5623 -1618 5633
rect -1652 5599 -1618 5623
rect -1652 5555 -1618 5561
rect -1652 5527 -1618 5555
rect -1652 5487 -1618 5489
rect -1652 5455 -1618 5487
rect -1652 5385 -1618 5417
rect -1652 5383 -1618 5385
rect -1652 5317 -1618 5345
rect -1652 5311 -1618 5317
rect -1652 5249 -1618 5273
rect -1652 5239 -1618 5249
rect -1652 5181 -1618 5201
rect -1652 5167 -1618 5181
rect -1652 5113 -1618 5129
rect -1652 5095 -1618 5113
rect -1652 5045 -1618 5057
rect -1652 5023 -1618 5045
rect -1652 4977 -1618 4985
rect -1652 4951 -1618 4977
rect -1554 5895 -1520 5921
rect -1554 5887 -1520 5895
rect -1554 5827 -1520 5849
rect -1554 5815 -1520 5827
rect -1554 5759 -1520 5777
rect -1554 5743 -1520 5759
rect -1554 5691 -1520 5705
rect -1554 5671 -1520 5691
rect -1554 5623 -1520 5633
rect -1554 5599 -1520 5623
rect -1554 5555 -1520 5561
rect -1554 5527 -1520 5555
rect -1554 5487 -1520 5489
rect -1554 5455 -1520 5487
rect -1554 5385 -1520 5417
rect -1554 5383 -1520 5385
rect -1554 5317 -1520 5345
rect -1554 5311 -1520 5317
rect -1554 5249 -1520 5273
rect -1554 5239 -1520 5249
rect -1554 5181 -1520 5201
rect -1554 5167 -1520 5181
rect -1554 5113 -1520 5129
rect -1554 5095 -1520 5113
rect -1554 5045 -1520 5057
rect -1554 5023 -1520 5045
rect -1554 4977 -1520 4985
rect -1554 4951 -1520 4977
rect -1456 5895 -1422 5921
rect -1456 5887 -1422 5895
rect -1456 5827 -1422 5849
rect -1456 5815 -1422 5827
rect -1456 5759 -1422 5777
rect -1456 5743 -1422 5759
rect -1456 5691 -1422 5705
rect -1456 5671 -1422 5691
rect -1456 5623 -1422 5633
rect -1456 5599 -1422 5623
rect -1456 5555 -1422 5561
rect -1456 5527 -1422 5555
rect -1456 5487 -1422 5489
rect -1456 5455 -1422 5487
rect -1456 5385 -1422 5417
rect -1456 5383 -1422 5385
rect -1456 5317 -1422 5345
rect -1456 5311 -1422 5317
rect -1456 5249 -1422 5273
rect -1456 5239 -1422 5249
rect -1456 5181 -1422 5201
rect -1456 5167 -1422 5181
rect -1456 5113 -1422 5129
rect -1456 5095 -1422 5113
rect -1456 5045 -1422 5057
rect -1456 5023 -1422 5045
rect -1456 4977 -1422 4985
rect -1456 4951 -1422 4977
rect -1358 5895 -1324 5921
rect -1358 5887 -1324 5895
rect -1358 5827 -1324 5849
rect -1358 5815 -1324 5827
rect -1358 5759 -1324 5777
rect -1358 5743 -1324 5759
rect -1358 5691 -1324 5705
rect -1358 5671 -1324 5691
rect -1358 5623 -1324 5633
rect -1358 5599 -1324 5623
rect -1358 5555 -1324 5561
rect -1358 5527 -1324 5555
rect -1358 5487 -1324 5489
rect -1358 5455 -1324 5487
rect -1358 5385 -1324 5417
rect -1358 5383 -1324 5385
rect -1358 5317 -1324 5345
rect -1358 5311 -1324 5317
rect -1358 5249 -1324 5273
rect -1358 5239 -1324 5249
rect -1358 5181 -1324 5201
rect -1358 5167 -1324 5181
rect -1358 5113 -1324 5129
rect -1358 5095 -1324 5113
rect -1358 5045 -1324 5057
rect -1358 5023 -1324 5045
rect -1358 4977 -1324 4985
rect -1358 4951 -1324 4977
rect -1260 5895 -1226 5921
rect -1260 5887 -1226 5895
rect -1260 5827 -1226 5849
rect -1260 5815 -1226 5827
rect -1260 5759 -1226 5777
rect -1260 5743 -1226 5759
rect -1260 5691 -1226 5705
rect -1260 5671 -1226 5691
rect -1260 5623 -1226 5633
rect -1260 5599 -1226 5623
rect -1260 5555 -1226 5561
rect -1260 5527 -1226 5555
rect -1260 5487 -1226 5489
rect -1260 5455 -1226 5487
rect -1260 5385 -1226 5417
rect -1260 5383 -1226 5385
rect -1260 5317 -1226 5345
rect -1260 5311 -1226 5317
rect -1260 5249 -1226 5273
rect -1260 5239 -1226 5249
rect -1260 5181 -1226 5201
rect -1260 5167 -1226 5181
rect -1260 5113 -1226 5129
rect -1260 5095 -1226 5113
rect -1260 5045 -1226 5057
rect -1260 5023 -1226 5045
rect -1260 4977 -1226 4985
rect -1260 4951 -1226 4977
rect -1162 5895 -1128 5921
rect -1162 5887 -1128 5895
rect -1162 5827 -1128 5849
rect -1162 5815 -1128 5827
rect -1162 5759 -1128 5777
rect -1162 5743 -1128 5759
rect -1162 5691 -1128 5705
rect -1162 5671 -1128 5691
rect -1162 5623 -1128 5633
rect -1162 5599 -1128 5623
rect -1162 5555 -1128 5561
rect -1162 5527 -1128 5555
rect -1162 5487 -1128 5489
rect -1162 5455 -1128 5487
rect -1162 5385 -1128 5417
rect -1162 5383 -1128 5385
rect -1162 5317 -1128 5345
rect -1162 5311 -1128 5317
rect -1162 5249 -1128 5273
rect -1162 5239 -1128 5249
rect -1162 5181 -1128 5201
rect -1162 5167 -1128 5181
rect -1162 5113 -1128 5129
rect -1162 5095 -1128 5113
rect -1162 5045 -1128 5057
rect -1162 5023 -1128 5045
rect -1162 4977 -1128 4985
rect -1162 4951 -1128 4977
rect -1064 5895 -1030 5921
rect -1064 5887 -1030 5895
rect -1064 5827 -1030 5849
rect -1064 5815 -1030 5827
rect -1064 5759 -1030 5777
rect -1064 5743 -1030 5759
rect -1064 5691 -1030 5705
rect -1064 5671 -1030 5691
rect -1064 5623 -1030 5633
rect -1064 5599 -1030 5623
rect -1064 5555 -1030 5561
rect -1064 5527 -1030 5555
rect -1064 5487 -1030 5489
rect -1064 5455 -1030 5487
rect -1064 5385 -1030 5417
rect -1064 5383 -1030 5385
rect -1064 5317 -1030 5345
rect -1064 5311 -1030 5317
rect -1064 5249 -1030 5273
rect -1064 5239 -1030 5249
rect -1064 5181 -1030 5201
rect -1064 5167 -1030 5181
rect -1064 5113 -1030 5129
rect -1064 5095 -1030 5113
rect -1064 5045 -1030 5057
rect -1064 5023 -1030 5045
rect -1064 4977 -1030 4985
rect -1064 4951 -1030 4977
rect -966 5895 -932 5921
rect -966 5887 -932 5895
rect -966 5827 -932 5849
rect -966 5815 -932 5827
rect -966 5759 -932 5777
rect -966 5743 -932 5759
rect -966 5691 -932 5705
rect -966 5671 -932 5691
rect -966 5623 -932 5633
rect -966 5599 -932 5623
rect -966 5555 -932 5561
rect -966 5527 -932 5555
rect -966 5487 -932 5489
rect -966 5455 -932 5487
rect -966 5385 -932 5417
rect -966 5383 -932 5385
rect -966 5317 -932 5345
rect -966 5311 -932 5317
rect -966 5249 -932 5273
rect -966 5239 -932 5249
rect -966 5181 -932 5201
rect -966 5167 -932 5181
rect -966 5113 -932 5129
rect -966 5095 -932 5113
rect -966 5045 -932 5057
rect -966 5023 -932 5045
rect -966 4977 -932 4985
rect -966 4951 -932 4977
rect -868 5895 -834 5921
rect -868 5887 -834 5895
rect -868 5827 -834 5849
rect -868 5815 -834 5827
rect -868 5759 -834 5777
rect -868 5743 -834 5759
rect -868 5691 -834 5705
rect -868 5671 -834 5691
rect -868 5623 -834 5633
rect -868 5599 -834 5623
rect 194 5987 228 6015
rect 194 5981 228 5987
rect 194 5919 228 5943
rect 194 5909 228 5919
rect 194 5851 228 5871
rect 194 5837 228 5851
rect 194 5783 228 5799
rect 194 5765 228 5783
rect 194 5715 228 5727
rect 194 5693 228 5715
rect 194 5647 228 5655
rect 194 5621 228 5647
rect 290 6565 324 6591
rect 290 6557 324 6565
rect 290 6497 324 6519
rect 290 6485 324 6497
rect 290 6429 324 6447
rect 290 6413 324 6429
rect 290 6361 324 6375
rect 290 6341 324 6361
rect 290 6293 324 6303
rect 290 6269 324 6293
rect 290 6225 324 6231
rect 290 6197 324 6225
rect 290 6157 324 6159
rect 290 6125 324 6157
rect 290 6055 324 6087
rect 290 6053 324 6055
rect 290 5987 324 6015
rect 290 5981 324 5987
rect 290 5919 324 5943
rect 290 5909 324 5919
rect 290 5851 324 5871
rect 290 5837 324 5851
rect 290 5783 324 5799
rect 290 5765 324 5783
rect 290 5715 324 5727
rect 290 5693 324 5715
rect 290 5647 324 5655
rect 290 5621 324 5647
rect -868 5555 -834 5561
rect -868 5527 -834 5555
rect 386 6565 420 6591
rect 386 6557 420 6565
rect 386 6497 420 6519
rect 386 6485 420 6497
rect 386 6429 420 6447
rect 386 6413 420 6429
rect 386 6361 420 6375
rect 386 6341 420 6361
rect 386 6293 420 6303
rect 386 6269 420 6293
rect 386 6225 420 6231
rect 386 6197 420 6225
rect 386 6157 420 6159
rect 386 6125 420 6157
rect 386 6055 420 6087
rect 386 6053 420 6055
rect 386 5987 420 6015
rect 386 5981 420 5987
rect 386 5919 420 5943
rect 386 5909 420 5919
rect 386 5851 420 5871
rect 386 5837 420 5851
rect 386 5783 420 5799
rect 386 5765 420 5783
rect 386 5715 420 5727
rect 386 5693 420 5715
rect 386 5647 420 5655
rect 386 5621 420 5647
rect 482 6565 516 6591
rect 482 6557 516 6565
rect 482 6497 516 6519
rect 482 6485 516 6497
rect 482 6429 516 6447
rect 482 6413 516 6429
rect 482 6361 516 6375
rect 482 6341 516 6361
rect 482 6293 516 6303
rect 482 6269 516 6293
rect 482 6225 516 6231
rect 482 6197 516 6225
rect 482 6157 516 6159
rect 482 6125 516 6157
rect 482 6055 516 6087
rect 482 6053 516 6055
rect 482 5987 516 6015
rect 482 5981 516 5987
rect 482 5919 516 5943
rect 482 5909 516 5919
rect 482 5851 516 5871
rect 482 5837 516 5851
rect 482 5783 516 5799
rect 482 5765 516 5783
rect 482 5715 516 5727
rect 482 5693 516 5715
rect 482 5647 516 5655
rect 482 5621 516 5647
rect 578 6565 612 6591
rect 578 6557 612 6565
rect 578 6497 612 6519
rect 578 6485 612 6497
rect 578 6429 612 6447
rect 578 6413 612 6429
rect 578 6361 612 6375
rect 578 6341 612 6361
rect 578 6293 612 6303
rect 578 6269 612 6293
rect 578 6225 612 6231
rect 578 6197 612 6225
rect 578 6157 612 6159
rect 578 6125 612 6157
rect 578 6055 612 6087
rect 578 6053 612 6055
rect 578 5987 612 6015
rect 578 5981 612 5987
rect 578 5919 612 5943
rect 578 5909 612 5919
rect 578 5851 612 5871
rect 578 5837 612 5851
rect 578 5783 612 5799
rect 578 5765 612 5783
rect 578 5715 612 5727
rect 578 5693 612 5715
rect 578 5647 612 5655
rect 578 5621 612 5647
rect 674 6565 708 6591
rect 674 6557 708 6565
rect 674 6497 708 6519
rect 674 6485 708 6497
rect 674 6429 708 6447
rect 674 6413 708 6429
rect 674 6361 708 6375
rect 674 6341 708 6361
rect 674 6293 708 6303
rect 674 6269 708 6293
rect 674 6225 708 6231
rect 674 6197 708 6225
rect 674 6157 708 6159
rect 674 6125 708 6157
rect 674 6055 708 6087
rect 674 6053 708 6055
rect 674 5987 708 6015
rect 674 5981 708 5987
rect 674 5919 708 5943
rect 674 5909 708 5919
rect 674 5851 708 5871
rect 674 5837 708 5851
rect 674 5783 708 5799
rect 674 5765 708 5783
rect 674 5715 708 5727
rect 674 5693 708 5715
rect 674 5647 708 5655
rect 674 5621 708 5647
rect 770 6565 804 6591
rect 770 6557 804 6565
rect 770 6497 804 6519
rect 770 6485 804 6497
rect 770 6429 804 6447
rect 770 6413 804 6429
rect 770 6361 804 6375
rect 770 6341 804 6361
rect 770 6293 804 6303
rect 770 6269 804 6293
rect 770 6225 804 6231
rect 770 6197 804 6225
rect 770 6157 804 6159
rect 770 6125 804 6157
rect 770 6055 804 6087
rect 770 6053 804 6055
rect 770 5987 804 6015
rect 770 5981 804 5987
rect 770 5919 804 5943
rect 770 5909 804 5919
rect 770 5851 804 5871
rect 770 5837 804 5851
rect 770 5783 804 5799
rect 770 5765 804 5783
rect 770 5715 804 5727
rect 770 5693 804 5715
rect 770 5647 804 5655
rect 770 5621 804 5647
rect 866 6565 900 6591
rect 866 6557 900 6565
rect 866 6497 900 6519
rect 866 6485 900 6497
rect 866 6429 900 6447
rect 866 6413 900 6429
rect 866 6361 900 6375
rect 866 6341 900 6361
rect 866 6293 900 6303
rect 866 6269 900 6293
rect 866 6225 900 6231
rect 866 6197 900 6225
rect 866 6157 900 6159
rect 866 6125 900 6157
rect 866 6055 900 6087
rect 866 6053 900 6055
rect 866 5987 900 6015
rect 866 5981 900 5987
rect 866 5919 900 5943
rect 866 5909 900 5919
rect 866 5851 900 5871
rect 866 5837 900 5851
rect 866 5783 900 5799
rect 866 5765 900 5783
rect 866 5715 900 5727
rect 866 5693 900 5715
rect 866 5647 900 5655
rect 866 5621 900 5647
rect 962 6565 996 6591
rect 962 6557 996 6565
rect 962 6497 996 6519
rect 962 6485 996 6497
rect 962 6429 996 6447
rect 962 6413 996 6429
rect 962 6361 996 6375
rect 962 6341 996 6361
rect 962 6293 996 6303
rect 962 6269 996 6293
rect 962 6225 996 6231
rect 962 6197 996 6225
rect 962 6157 996 6159
rect 962 6125 996 6157
rect 962 6055 996 6087
rect 962 6053 996 6055
rect 962 5987 996 6015
rect 962 5981 996 5987
rect 962 5919 996 5943
rect 962 5909 996 5919
rect 962 5851 996 5871
rect 962 5837 996 5851
rect 962 5783 996 5799
rect 962 5765 996 5783
rect 962 5715 996 5727
rect 962 5693 996 5715
rect 962 5647 996 5655
rect 962 5621 996 5647
rect 1058 6565 1092 6591
rect 1058 6557 1092 6565
rect 1058 6497 1092 6519
rect 1058 6485 1092 6497
rect 1058 6429 1092 6447
rect 1058 6413 1092 6429
rect 1058 6361 1092 6375
rect 1058 6341 1092 6361
rect 1058 6293 1092 6303
rect 1058 6269 1092 6293
rect 1058 6225 1092 6231
rect 1058 6197 1092 6225
rect 1058 6157 1092 6159
rect 1058 6125 1092 6157
rect 1058 6055 1092 6087
rect 1058 6053 1092 6055
rect 1058 5987 1092 6015
rect 1058 5981 1092 5987
rect 1058 5919 1092 5943
rect 1058 5909 1092 5919
rect 1058 5851 1092 5871
rect 1058 5837 1092 5851
rect 1058 5783 1092 5799
rect 1058 5765 1092 5783
rect 1058 5715 1092 5727
rect 1058 5693 1092 5715
rect 1058 5647 1092 5655
rect 1058 5621 1092 5647
rect 1154 6565 1188 6591
rect 1154 6557 1188 6565
rect 1154 6497 1188 6519
rect 1154 6485 1188 6497
rect 1154 6429 1188 6447
rect 1154 6413 1188 6429
rect 1154 6361 1188 6375
rect 1154 6341 1188 6361
rect 1154 6293 1188 6303
rect 1154 6269 1188 6293
rect 1154 6225 1188 6231
rect 1154 6197 1188 6225
rect 1154 6157 1188 6159
rect 1154 6125 1188 6157
rect 1154 6055 1188 6087
rect 1154 6053 1188 6055
rect 1154 5987 1188 6015
rect 1154 5981 1188 5987
rect 1154 5919 1188 5943
rect 1154 5909 1188 5919
rect 1154 5851 1188 5871
rect 1154 5837 1188 5851
rect 1154 5783 1188 5799
rect 1154 5765 1188 5783
rect 1154 5715 1188 5727
rect 1154 5693 1188 5715
rect 1154 5647 1188 5655
rect 1154 5621 1188 5647
rect 1250 6565 1284 6591
rect 1250 6557 1284 6565
rect 1250 6497 1284 6519
rect 1250 6485 1284 6497
rect 1250 6429 1284 6447
rect 1250 6413 1284 6429
rect 1250 6361 1284 6375
rect 1250 6341 1284 6361
rect 1250 6293 1284 6303
rect 1250 6269 1284 6293
rect 1250 6225 1284 6231
rect 1250 6197 1284 6225
rect 1250 6157 1284 6159
rect 1250 6125 1284 6157
rect 1250 6055 1284 6087
rect 1250 6053 1284 6055
rect 1250 5987 1284 6015
rect 1250 5981 1284 5987
rect 1250 5919 1284 5943
rect 1250 5909 1284 5919
rect 1250 5851 1284 5871
rect 1250 5837 1284 5851
rect 1250 5783 1284 5799
rect 1250 5765 1284 5783
rect 1250 5715 1284 5727
rect 1250 5693 1284 5715
rect 1250 5647 1284 5655
rect 1250 5621 1284 5647
rect 1346 6565 1380 6591
rect 1346 6557 1380 6565
rect 1346 6497 1380 6519
rect 1346 6485 1380 6497
rect 1346 6429 1380 6447
rect 1346 6413 1380 6429
rect 1346 6361 1380 6375
rect 1346 6341 1380 6361
rect 1346 6293 1380 6303
rect 1346 6269 1380 6293
rect 1346 6225 1380 6231
rect 1346 6197 1380 6225
rect 1346 6157 1380 6159
rect 1346 6125 1380 6157
rect 1346 6055 1380 6087
rect 1346 6053 1380 6055
rect 1346 5987 1380 6015
rect 1346 5981 1380 5987
rect 1346 5919 1380 5943
rect 1346 5909 1380 5919
rect 1346 5851 1380 5871
rect 1346 5837 1380 5851
rect 1346 5783 1380 5799
rect 1346 5765 1380 5783
rect 1346 5715 1380 5727
rect 1346 5693 1380 5715
rect 1346 5647 1380 5655
rect 1346 5621 1380 5647
rect 1960 6561 1994 6587
rect 1960 6553 1994 6561
rect 1960 6493 1994 6515
rect 1960 6481 1994 6493
rect 1960 6425 1994 6443
rect 1960 6409 1994 6425
rect 1960 6357 1994 6371
rect 1960 6337 1994 6357
rect 1960 6289 1994 6299
rect 1960 6265 1994 6289
rect 1960 6221 1994 6227
rect 1960 6193 1994 6221
rect 1960 6153 1994 6155
rect 1960 6121 1994 6153
rect 1960 6051 1994 6083
rect 1960 6049 1994 6051
rect 1960 5983 1994 6011
rect 1960 5977 1994 5983
rect 1960 5915 1994 5939
rect 1960 5905 1994 5915
rect 1960 5847 1994 5867
rect 1960 5833 1994 5847
rect 1960 5779 1994 5795
rect 1960 5761 1994 5779
rect 1960 5711 1994 5723
rect 1960 5689 1994 5711
rect 1960 5643 1994 5651
rect 1960 5617 1994 5643
rect 2056 6561 2090 6587
rect 2056 6553 2090 6561
rect 2056 6493 2090 6515
rect 2056 6481 2090 6493
rect 2056 6425 2090 6443
rect 2056 6409 2090 6425
rect 2056 6357 2090 6371
rect 2056 6337 2090 6357
rect 2056 6289 2090 6299
rect 2056 6265 2090 6289
rect 2056 6221 2090 6227
rect 2056 6193 2090 6221
rect 2056 6153 2090 6155
rect 2056 6121 2090 6153
rect 2056 6051 2090 6083
rect 2056 6049 2090 6051
rect 2056 5983 2090 6011
rect 2056 5977 2090 5983
rect 2056 5915 2090 5939
rect 2056 5905 2090 5915
rect 2056 5847 2090 5867
rect 2056 5833 2090 5847
rect 2056 5779 2090 5795
rect 2056 5761 2090 5779
rect 2056 5711 2090 5723
rect 2056 5689 2090 5711
rect 2056 5643 2090 5651
rect 2056 5617 2090 5643
rect 2152 6561 2186 6587
rect 2152 6553 2186 6561
rect 2152 6493 2186 6515
rect 2152 6481 2186 6493
rect 2152 6425 2186 6443
rect 2152 6409 2186 6425
rect 2152 6357 2186 6371
rect 2152 6337 2186 6357
rect 2152 6289 2186 6299
rect 2152 6265 2186 6289
rect 2152 6221 2186 6227
rect 2152 6193 2186 6221
rect 2152 6153 2186 6155
rect 2152 6121 2186 6153
rect 2152 6051 2186 6083
rect 2152 6049 2186 6051
rect 2152 5983 2186 6011
rect 2152 5977 2186 5983
rect 2152 5915 2186 5939
rect 2152 5905 2186 5915
rect 2152 5847 2186 5867
rect 2152 5833 2186 5847
rect 2152 5779 2186 5795
rect 2152 5761 2186 5779
rect 2152 5711 2186 5723
rect 2152 5689 2186 5711
rect 2152 5643 2186 5651
rect 2152 5617 2186 5643
rect 2248 6561 2282 6587
rect 2248 6553 2282 6561
rect 2248 6493 2282 6515
rect 2248 6481 2282 6493
rect 2248 6425 2282 6443
rect 2248 6409 2282 6425
rect 2248 6357 2282 6371
rect 2248 6337 2282 6357
rect 2248 6289 2282 6299
rect 2248 6265 2282 6289
rect 2248 6221 2282 6227
rect 2248 6193 2282 6221
rect 2248 6153 2282 6155
rect 2248 6121 2282 6153
rect 2248 6051 2282 6083
rect 2248 6049 2282 6051
rect 2248 5983 2282 6011
rect 2248 5977 2282 5983
rect 2248 5915 2282 5939
rect 2248 5905 2282 5915
rect 2248 5847 2282 5867
rect 2248 5833 2282 5847
rect 2248 5779 2282 5795
rect 2248 5761 2282 5779
rect 2248 5711 2282 5723
rect 2248 5689 2282 5711
rect 2248 5643 2282 5651
rect 2248 5617 2282 5643
rect 2344 6561 2378 6587
rect 2344 6553 2378 6561
rect 2344 6493 2378 6515
rect 2344 6481 2378 6493
rect 2344 6425 2378 6443
rect 2344 6409 2378 6425
rect 2344 6357 2378 6371
rect 2344 6337 2378 6357
rect 2344 6289 2378 6299
rect 2344 6265 2378 6289
rect 2344 6221 2378 6227
rect 2344 6193 2378 6221
rect 2344 6153 2378 6155
rect 2344 6121 2378 6153
rect 2344 6051 2378 6083
rect 2344 6049 2378 6051
rect 2344 5983 2378 6011
rect 2344 5977 2378 5983
rect 2344 5915 2378 5939
rect 2344 5905 2378 5915
rect 2344 5847 2378 5867
rect 2344 5833 2378 5847
rect 2344 5779 2378 5795
rect 2344 5761 2378 5779
rect 2344 5711 2378 5723
rect 2344 5689 2378 5711
rect 2344 5643 2378 5651
rect 2344 5617 2378 5643
rect 2440 6561 2474 6587
rect 2440 6553 2474 6561
rect 2440 6493 2474 6515
rect 2440 6481 2474 6493
rect 2440 6425 2474 6443
rect 2440 6409 2474 6425
rect 2440 6357 2474 6371
rect 2440 6337 2474 6357
rect 2440 6289 2474 6299
rect 2440 6265 2474 6289
rect 2440 6221 2474 6227
rect 2440 6193 2474 6221
rect 2440 6153 2474 6155
rect 2440 6121 2474 6153
rect 2440 6051 2474 6083
rect 2440 6049 2474 6051
rect 2440 5983 2474 6011
rect 2440 5977 2474 5983
rect 2440 5915 2474 5939
rect 2440 5905 2474 5915
rect 2440 5847 2474 5867
rect 2440 5833 2474 5847
rect 2440 5779 2474 5795
rect 2440 5761 2474 5779
rect 2440 5711 2474 5723
rect 2440 5689 2474 5711
rect 2440 5643 2474 5651
rect 2440 5617 2474 5643
rect 2536 6561 2570 6587
rect 2536 6553 2570 6561
rect 2536 6493 2570 6515
rect 2536 6481 2570 6493
rect 2536 6425 2570 6443
rect 2536 6409 2570 6425
rect 2536 6357 2570 6371
rect 2536 6337 2570 6357
rect 2536 6289 2570 6299
rect 2536 6265 2570 6289
rect 2536 6221 2570 6227
rect 2536 6193 2570 6221
rect 2536 6153 2570 6155
rect 2536 6121 2570 6153
rect 2536 6051 2570 6083
rect 2536 6049 2570 6051
rect 2536 5983 2570 6011
rect 2536 5977 2570 5983
rect 2536 5915 2570 5939
rect 2536 5905 2570 5915
rect 2536 5847 2570 5867
rect 2536 5833 2570 5847
rect 2536 5779 2570 5795
rect 2536 5761 2570 5779
rect 2536 5711 2570 5723
rect 2536 5689 2570 5711
rect 2536 5643 2570 5651
rect 2536 5617 2570 5643
rect 2632 6561 2666 6587
rect 2632 6553 2666 6561
rect 2632 6493 2666 6515
rect 2632 6481 2666 6493
rect 2632 6425 2666 6443
rect 2632 6409 2666 6425
rect 2632 6357 2666 6371
rect 2632 6337 2666 6357
rect 2632 6289 2666 6299
rect 2632 6265 2666 6289
rect 2632 6221 2666 6227
rect 2632 6193 2666 6221
rect 2632 6153 2666 6155
rect 2632 6121 2666 6153
rect 2632 6051 2666 6083
rect 2632 6049 2666 6051
rect 2632 5983 2666 6011
rect 2632 5977 2666 5983
rect 2632 5915 2666 5939
rect 2632 5905 2666 5915
rect 2632 5847 2666 5867
rect 2632 5833 2666 5847
rect 2632 5779 2666 5795
rect 2632 5761 2666 5779
rect 2632 5711 2666 5723
rect 2632 5689 2666 5711
rect 2632 5643 2666 5651
rect 2632 5617 2666 5643
rect 2728 6561 2762 6587
rect 2728 6553 2762 6561
rect 2728 6493 2762 6515
rect 2728 6481 2762 6493
rect 2728 6425 2762 6443
rect 2728 6409 2762 6425
rect 2728 6357 2762 6371
rect 2728 6337 2762 6357
rect 2728 6289 2762 6299
rect 2728 6265 2762 6289
rect 2728 6221 2762 6227
rect 2728 6193 2762 6221
rect 2728 6153 2762 6155
rect 2728 6121 2762 6153
rect 2728 6051 2762 6083
rect 2728 6049 2762 6051
rect 2728 5983 2762 6011
rect 2728 5977 2762 5983
rect 2728 5915 2762 5939
rect 2728 5905 2762 5915
rect 2728 5847 2762 5867
rect 2728 5833 2762 5847
rect 2728 5779 2762 5795
rect 2728 5761 2762 5779
rect 2728 5711 2762 5723
rect 2728 5689 2762 5711
rect 2728 5643 2762 5651
rect 2728 5617 2762 5643
rect 7486 6774 7680 6878
rect 9838 6840 9872 6874
rect 8426 6738 8460 6772
rect 8714 6753 8748 6787
rect 9362 6755 9396 6789
rect 3150 6549 3184 6575
rect 3150 6541 3184 6549
rect 3150 6481 3184 6503
rect 3150 6469 3184 6481
rect 3150 6413 3184 6431
rect 3150 6397 3184 6413
rect 3150 6345 3184 6359
rect 3150 6325 3184 6345
rect 3150 6277 3184 6287
rect 3150 6253 3184 6277
rect 3150 6209 3184 6215
rect 3150 6181 3184 6209
rect 3150 6141 3184 6143
rect 3150 6109 3184 6141
rect 3150 6039 3184 6071
rect 3150 6037 3184 6039
rect 3150 5971 3184 5999
rect 3150 5965 3184 5971
rect 3150 5903 3184 5927
rect 3150 5893 3184 5903
rect 3150 5835 3184 5855
rect 3150 5821 3184 5835
rect 3150 5767 3184 5783
rect 3150 5749 3184 5767
rect 3150 5699 3184 5711
rect 3150 5677 3184 5699
rect 3150 5631 3184 5639
rect 3150 5605 3184 5631
rect 3246 6549 3280 6575
rect 3246 6541 3280 6549
rect 3246 6481 3280 6503
rect 3246 6469 3280 6481
rect 3246 6413 3280 6431
rect 3246 6397 3280 6413
rect 3246 6345 3280 6359
rect 3246 6325 3280 6345
rect 3246 6277 3280 6287
rect 3246 6253 3280 6277
rect 3246 6209 3280 6215
rect 3246 6181 3280 6209
rect 3246 6141 3280 6143
rect 3246 6109 3280 6141
rect 3246 6039 3280 6071
rect 3246 6037 3280 6039
rect 3246 5971 3280 5999
rect 3246 5965 3280 5971
rect 3246 5903 3280 5927
rect 3246 5893 3280 5903
rect 3246 5835 3280 5855
rect 3246 5821 3280 5835
rect 3246 5767 3280 5783
rect 3246 5749 3280 5767
rect 3246 5699 3280 5711
rect 3246 5677 3280 5699
rect 3246 5631 3280 5639
rect 3246 5605 3280 5631
rect -868 5487 -834 5489
rect -868 5455 -834 5487
rect -868 5385 -834 5417
rect -868 5383 -834 5385
rect 3342 6549 3376 6575
rect 3342 6541 3376 6549
rect 3342 6481 3376 6503
rect 3342 6469 3376 6481
rect 3342 6413 3376 6431
rect 3342 6397 3376 6413
rect 3342 6345 3376 6359
rect 3342 6325 3376 6345
rect 3342 6277 3376 6287
rect 3342 6253 3376 6277
rect 3342 6209 3376 6215
rect 3342 6181 3376 6209
rect 3342 6141 3376 6143
rect 3342 6109 3376 6141
rect 3342 6039 3376 6071
rect 3342 6037 3376 6039
rect 3342 5971 3376 5999
rect 3342 5965 3376 5971
rect 3342 5903 3376 5927
rect 3342 5893 3376 5903
rect 3342 5835 3376 5855
rect 3342 5821 3376 5835
rect 3342 5767 3376 5783
rect 3342 5749 3376 5767
rect 3342 5699 3376 5711
rect 3342 5677 3376 5699
rect 3342 5631 3376 5639
rect 3342 5605 3376 5631
rect 3438 6549 3472 6575
rect 3438 6541 3472 6549
rect 3438 6481 3472 6503
rect 3438 6469 3472 6481
rect 3438 6413 3472 6431
rect 3438 6397 3472 6413
rect 3438 6345 3472 6359
rect 3438 6325 3472 6345
rect 3438 6277 3472 6287
rect 3438 6253 3472 6277
rect 3438 6209 3472 6215
rect 3438 6181 3472 6209
rect 3438 6141 3472 6143
rect 3438 6109 3472 6141
rect 3438 6039 3472 6071
rect 3438 6037 3472 6039
rect 3438 5971 3472 5999
rect 3438 5965 3472 5971
rect 3438 5903 3472 5927
rect 3438 5893 3472 5903
rect 3438 5835 3472 5855
rect 3438 5821 3472 5835
rect 3438 5767 3472 5783
rect 3438 5749 3472 5767
rect 3438 5699 3472 5711
rect 3438 5677 3472 5699
rect 3438 5631 3472 5639
rect 3438 5605 3472 5631
rect 3534 6549 3568 6575
rect 3534 6541 3568 6549
rect 3534 6481 3568 6503
rect 3534 6469 3568 6481
rect 3534 6413 3568 6431
rect 3534 6397 3568 6413
rect 3534 6345 3568 6359
rect 3534 6325 3568 6345
rect 3534 6277 3568 6287
rect 3534 6253 3568 6277
rect 3534 6209 3568 6215
rect 3534 6181 3568 6209
rect 3534 6141 3568 6143
rect 3534 6109 3568 6141
rect 3534 6039 3568 6071
rect 3534 6037 3568 6039
rect 3534 5971 3568 5999
rect 3534 5965 3568 5971
rect 3534 5903 3568 5927
rect 3534 5893 3568 5903
rect 3534 5835 3568 5855
rect 3534 5821 3568 5835
rect 3534 5767 3568 5783
rect 3534 5749 3568 5767
rect 3534 5699 3568 5711
rect 3534 5677 3568 5699
rect 3534 5631 3568 5639
rect 3534 5605 3568 5631
rect 3630 6549 3664 6575
rect 3630 6541 3664 6549
rect 3630 6481 3664 6503
rect 3630 6469 3664 6481
rect 3630 6413 3664 6431
rect 3630 6397 3664 6413
rect 3630 6345 3664 6359
rect 3630 6325 3664 6345
rect 3630 6277 3664 6287
rect 3630 6253 3664 6277
rect 3630 6209 3664 6215
rect 3630 6181 3664 6209
rect 3630 6141 3664 6143
rect 3630 6109 3664 6141
rect 3630 6039 3664 6071
rect 3630 6037 3664 6039
rect 3630 5971 3664 5999
rect 3630 5965 3664 5971
rect 3630 5903 3664 5927
rect 3630 5893 3664 5903
rect 3630 5835 3664 5855
rect 3630 5821 3664 5835
rect 3630 5767 3664 5783
rect 3630 5749 3664 5767
rect 3630 5699 3664 5711
rect 3630 5677 3664 5699
rect 3630 5631 3664 5639
rect 3630 5605 3664 5631
rect 3726 6549 3760 6575
rect 3726 6541 3760 6549
rect 3726 6481 3760 6503
rect 3726 6469 3760 6481
rect 3726 6413 3760 6431
rect 3726 6397 3760 6413
rect 3726 6345 3760 6359
rect 3726 6325 3760 6345
rect 3726 6277 3760 6287
rect 3726 6253 3760 6277
rect 3726 6209 3760 6215
rect 3726 6181 3760 6209
rect 3726 6141 3760 6143
rect 3726 6109 3760 6141
rect 3726 6039 3760 6071
rect 3726 6037 3760 6039
rect 3726 5971 3760 5999
rect 3726 5965 3760 5971
rect 3726 5903 3760 5927
rect 3726 5893 3760 5903
rect 3726 5835 3760 5855
rect 3726 5821 3760 5835
rect 3726 5767 3760 5783
rect 3726 5749 3760 5767
rect 3726 5699 3760 5711
rect 3726 5677 3760 5699
rect 3726 5631 3760 5639
rect 3726 5605 3760 5631
rect 3822 6549 3856 6575
rect 3822 6541 3856 6549
rect 3822 6481 3856 6503
rect 3822 6469 3856 6481
rect 3822 6413 3856 6431
rect 3822 6397 3856 6413
rect 3822 6345 3856 6359
rect 3822 6325 3856 6345
rect 3822 6277 3856 6287
rect 3822 6253 3856 6277
rect 3822 6209 3856 6215
rect 3822 6181 3856 6209
rect 3822 6141 3856 6143
rect 3822 6109 3856 6141
rect 3822 6039 3856 6071
rect 3822 6037 3856 6039
rect 3822 5971 3856 5999
rect 3822 5965 3856 5971
rect 3822 5903 3856 5927
rect 3822 5893 3856 5903
rect 3822 5835 3856 5855
rect 3822 5821 3856 5835
rect 3822 5767 3856 5783
rect 3822 5749 3856 5767
rect 3822 5699 3856 5711
rect 3822 5677 3856 5699
rect 3822 5631 3856 5639
rect 3822 5605 3856 5631
rect 3918 6549 3952 6575
rect 3918 6541 3952 6549
rect 3918 6481 3952 6503
rect 3918 6469 3952 6481
rect 3918 6413 3952 6431
rect 3918 6397 3952 6413
rect 3918 6345 3952 6359
rect 3918 6325 3952 6345
rect 3918 6277 3952 6287
rect 3918 6253 3952 6277
rect 3918 6209 3952 6215
rect 3918 6181 3952 6209
rect 3918 6141 3952 6143
rect 3918 6109 3952 6141
rect 3918 6039 3952 6071
rect 3918 6037 3952 6039
rect 3918 5971 3952 5999
rect 3918 5965 3952 5971
rect 3918 5903 3952 5927
rect 3918 5893 3952 5903
rect 3918 5835 3952 5855
rect 3918 5821 3952 5835
rect 3918 5767 3952 5783
rect 3918 5749 3952 5767
rect 3918 5699 3952 5711
rect 3918 5677 3952 5699
rect 3918 5631 3952 5639
rect 3918 5605 3952 5631
rect 4014 6549 4048 6575
rect 4014 6541 4048 6549
rect 4014 6481 4048 6503
rect 4014 6469 4048 6481
rect 4014 6413 4048 6431
rect 4014 6397 4048 6413
rect 4014 6345 4048 6359
rect 4014 6325 4048 6345
rect 4014 6277 4048 6287
rect 4014 6253 4048 6277
rect 4014 6209 4048 6215
rect 4014 6181 4048 6209
rect 4014 6141 4048 6143
rect 4014 6109 4048 6141
rect 4014 6039 4048 6071
rect 4014 6037 4048 6039
rect 4014 5971 4048 5999
rect 4014 5965 4048 5971
rect 4014 5903 4048 5927
rect 4014 5893 4048 5903
rect 4014 5835 4048 5855
rect 4014 5821 4048 5835
rect 4014 5767 4048 5783
rect 4014 5749 4048 5767
rect 4014 5699 4048 5711
rect 4014 5677 4048 5699
rect 4014 5631 4048 5639
rect 4014 5605 4048 5631
rect 4110 6549 4144 6575
rect 4110 6541 4144 6549
rect 4110 6481 4144 6503
rect 4110 6469 4144 6481
rect 4110 6413 4144 6431
rect 4110 6397 4144 6413
rect 4110 6345 4144 6359
rect 4110 6325 4144 6345
rect 4110 6277 4144 6287
rect 4110 6253 4144 6277
rect 4110 6209 4144 6215
rect 4110 6181 4144 6209
rect 4110 6141 4144 6143
rect 4110 6109 4144 6141
rect 4110 6039 4144 6071
rect 4110 6037 4144 6039
rect 4110 5971 4144 5999
rect 4110 5965 4144 5971
rect 4110 5903 4144 5927
rect 4110 5893 4144 5903
rect 4110 5835 4144 5855
rect 4110 5821 4144 5835
rect 4110 5767 4144 5783
rect 4110 5749 4144 5767
rect 4110 5699 4144 5711
rect 4110 5677 4144 5699
rect 4110 5631 4144 5639
rect 4110 5605 4144 5631
rect 4206 6549 4240 6575
rect 4206 6541 4240 6549
rect 4206 6481 4240 6503
rect 4206 6469 4240 6481
rect 4206 6413 4240 6431
rect 4206 6397 4240 6413
rect 4206 6345 4240 6359
rect 4206 6325 4240 6345
rect 4206 6277 4240 6287
rect 4206 6253 4240 6277
rect 4206 6209 4240 6215
rect 4206 6181 4240 6209
rect 4206 6141 4240 6143
rect 4206 6109 4240 6141
rect 4206 6039 4240 6071
rect 4206 6037 4240 6039
rect 4206 5971 4240 5999
rect 4206 5965 4240 5971
rect 4206 5903 4240 5927
rect 4206 5893 4240 5903
rect 4206 5835 4240 5855
rect 4206 5821 4240 5835
rect 4206 5767 4240 5783
rect 4206 5749 4240 5767
rect 4206 5699 4240 5711
rect 4206 5677 4240 5699
rect 4206 5631 4240 5639
rect 4206 5605 4240 5631
rect 4302 6549 4336 6575
rect 4302 6541 4336 6549
rect 4302 6481 4336 6503
rect 4302 6469 4336 6481
rect 4302 6413 4336 6431
rect 4302 6397 4336 6413
rect 4302 6345 4336 6359
rect 4302 6325 4336 6345
rect 4302 6277 4336 6287
rect 4302 6253 4336 6277
rect 4302 6209 4336 6215
rect 4302 6181 4336 6209
rect 4302 6141 4336 6143
rect 4302 6109 4336 6141
rect 4302 6039 4336 6071
rect 4302 6037 4336 6039
rect 4302 5971 4336 5999
rect 4302 5965 4336 5971
rect 4302 5903 4336 5927
rect 4302 5893 4336 5903
rect 4302 5835 4336 5855
rect 4302 5821 4336 5835
rect 4302 5767 4336 5783
rect 4302 5749 4336 5767
rect 4302 5699 4336 5711
rect 4302 5677 4336 5699
rect 4302 5631 4336 5639
rect 4302 5605 4336 5631
rect 4916 6545 4950 6571
rect 4916 6537 4950 6545
rect 4916 6477 4950 6499
rect 4916 6465 4950 6477
rect 4916 6409 4950 6427
rect 4916 6393 4950 6409
rect 4916 6341 4950 6355
rect 4916 6321 4950 6341
rect 4916 6273 4950 6283
rect 4916 6249 4950 6273
rect 4916 6205 4950 6211
rect 4916 6177 4950 6205
rect 4916 6137 4950 6139
rect 4916 6105 4950 6137
rect 4916 6035 4950 6067
rect 4916 6033 4950 6035
rect 4916 5967 4950 5995
rect 4916 5961 4950 5967
rect 4916 5899 4950 5923
rect 4916 5889 4950 5899
rect 4916 5831 4950 5851
rect 4916 5817 4950 5831
rect 4916 5763 4950 5779
rect 4916 5745 4950 5763
rect 4916 5695 4950 5707
rect 4916 5673 4950 5695
rect 4916 5627 4950 5635
rect 4916 5601 4950 5627
rect 5012 6545 5046 6571
rect 5012 6537 5046 6545
rect 5012 6477 5046 6499
rect 5012 6465 5046 6477
rect 5012 6409 5046 6427
rect 5012 6393 5046 6409
rect 5012 6341 5046 6355
rect 5012 6321 5046 6341
rect 5012 6273 5046 6283
rect 5012 6249 5046 6273
rect 5012 6205 5046 6211
rect 5012 6177 5046 6205
rect 5012 6137 5046 6139
rect 5012 6105 5046 6137
rect 5012 6035 5046 6067
rect 5012 6033 5046 6035
rect 5012 5967 5046 5995
rect 5012 5961 5046 5967
rect 5012 5899 5046 5923
rect 5012 5889 5046 5899
rect 5012 5831 5046 5851
rect 5012 5817 5046 5831
rect 5012 5763 5046 5779
rect 5012 5745 5046 5763
rect 5012 5695 5046 5707
rect 5012 5673 5046 5695
rect 5012 5627 5046 5635
rect 5012 5601 5046 5627
rect 880 5372 982 5418
rect 5108 6545 5142 6571
rect 5108 6537 5142 6545
rect 5108 6477 5142 6499
rect 5108 6465 5142 6477
rect 5108 6409 5142 6427
rect 5108 6393 5142 6409
rect 5108 6341 5142 6355
rect 5108 6321 5142 6341
rect 5108 6273 5142 6283
rect 5108 6249 5142 6273
rect 5108 6205 5142 6211
rect 5108 6177 5142 6205
rect 5108 6137 5142 6139
rect 5108 6105 5142 6137
rect 5108 6035 5142 6067
rect 5108 6033 5142 6035
rect 5108 5967 5142 5995
rect 5108 5961 5142 5967
rect 5108 5899 5142 5923
rect 5108 5889 5142 5899
rect 5108 5831 5142 5851
rect 5108 5817 5142 5831
rect 5108 5763 5142 5779
rect 5108 5745 5142 5763
rect 5108 5695 5142 5707
rect 5108 5673 5142 5695
rect 5108 5627 5142 5635
rect 5108 5601 5142 5627
rect 5204 6545 5238 6571
rect 5204 6537 5238 6545
rect 5204 6477 5238 6499
rect 5204 6465 5238 6477
rect 5204 6409 5238 6427
rect 5204 6393 5238 6409
rect 5204 6341 5238 6355
rect 5204 6321 5238 6341
rect 5204 6273 5238 6283
rect 5204 6249 5238 6273
rect 5204 6205 5238 6211
rect 5204 6177 5238 6205
rect 5204 6137 5238 6139
rect 5204 6105 5238 6137
rect 5204 6035 5238 6067
rect 5204 6033 5238 6035
rect 5204 5967 5238 5995
rect 5204 5961 5238 5967
rect 5204 5899 5238 5923
rect 5204 5889 5238 5899
rect 5204 5831 5238 5851
rect 5204 5817 5238 5831
rect 5204 5763 5238 5779
rect 5204 5745 5238 5763
rect 5204 5695 5238 5707
rect 5204 5673 5238 5695
rect 5204 5627 5238 5635
rect 5204 5601 5238 5627
rect 5300 6545 5334 6571
rect 5300 6537 5334 6545
rect 5300 6477 5334 6499
rect 5300 6465 5334 6477
rect 5300 6409 5334 6427
rect 5300 6393 5334 6409
rect 5300 6341 5334 6355
rect 5300 6321 5334 6341
rect 5300 6273 5334 6283
rect 5300 6249 5334 6273
rect 5300 6205 5334 6211
rect 5300 6177 5334 6205
rect 5300 6137 5334 6139
rect 5300 6105 5334 6137
rect 5300 6035 5334 6067
rect 5300 6033 5334 6035
rect 5300 5967 5334 5995
rect 5300 5961 5334 5967
rect 5300 5899 5334 5923
rect 5300 5889 5334 5899
rect 5300 5831 5334 5851
rect 5300 5817 5334 5831
rect 5300 5763 5334 5779
rect 5300 5745 5334 5763
rect 5300 5695 5334 5707
rect 5300 5673 5334 5695
rect 5300 5627 5334 5635
rect 5300 5601 5334 5627
rect 5396 6545 5430 6571
rect 5396 6537 5430 6545
rect 5396 6477 5430 6499
rect 5396 6465 5430 6477
rect 5396 6409 5430 6427
rect 5396 6393 5430 6409
rect 5396 6341 5430 6355
rect 5396 6321 5430 6341
rect 5396 6273 5430 6283
rect 5396 6249 5430 6273
rect 5396 6205 5430 6211
rect 5396 6177 5430 6205
rect 5396 6137 5430 6139
rect 5396 6105 5430 6137
rect 5396 6035 5430 6067
rect 5396 6033 5430 6035
rect 5396 5967 5430 5995
rect 5396 5961 5430 5967
rect 5396 5899 5430 5923
rect 5396 5889 5430 5899
rect 5396 5831 5430 5851
rect 5396 5817 5430 5831
rect 5396 5763 5430 5779
rect 5396 5745 5430 5763
rect 5396 5695 5430 5707
rect 5396 5673 5430 5695
rect 5396 5627 5430 5635
rect 5396 5601 5430 5627
rect 5492 6545 5526 6571
rect 5492 6537 5526 6545
rect 5492 6477 5526 6499
rect 5492 6465 5526 6477
rect 5492 6409 5526 6427
rect 5492 6393 5526 6409
rect 5492 6341 5526 6355
rect 5492 6321 5526 6341
rect 5492 6273 5526 6283
rect 5492 6249 5526 6273
rect 5492 6205 5526 6211
rect 5492 6177 5526 6205
rect 5492 6137 5526 6139
rect 5492 6105 5526 6137
rect 5492 6035 5526 6067
rect 5492 6033 5526 6035
rect 5492 5967 5526 5995
rect 5492 5961 5526 5967
rect 5492 5899 5526 5923
rect 5492 5889 5526 5899
rect 5492 5831 5526 5851
rect 5492 5817 5526 5831
rect 5492 5763 5526 5779
rect 5492 5745 5526 5763
rect 5492 5695 5526 5707
rect 5492 5673 5526 5695
rect 5492 5627 5526 5635
rect 5492 5601 5526 5627
rect 5588 6545 5622 6571
rect 5588 6537 5622 6545
rect 5588 6477 5622 6499
rect 5588 6465 5622 6477
rect 5588 6409 5622 6427
rect 5588 6393 5622 6409
rect 5588 6341 5622 6355
rect 5588 6321 5622 6341
rect 5588 6273 5622 6283
rect 5588 6249 5622 6273
rect 5588 6205 5622 6211
rect 5588 6177 5622 6205
rect 5588 6137 5622 6139
rect 5588 6105 5622 6137
rect 5588 6035 5622 6067
rect 5588 6033 5622 6035
rect 5588 5967 5622 5995
rect 5588 5961 5622 5967
rect 5588 5899 5622 5923
rect 5588 5889 5622 5899
rect 5588 5831 5622 5851
rect 5588 5817 5622 5831
rect 5588 5763 5622 5779
rect 5588 5745 5622 5763
rect 5588 5695 5622 5707
rect 5588 5673 5622 5695
rect 5588 5627 5622 5635
rect 5588 5601 5622 5627
rect 5684 6545 5718 6571
rect 5684 6537 5718 6545
rect 5684 6477 5718 6499
rect 5684 6465 5718 6477
rect 5684 6409 5718 6427
rect 5684 6393 5718 6409
rect 5684 6341 5718 6355
rect 5684 6321 5718 6341
rect 5684 6273 5718 6283
rect 5684 6249 5718 6273
rect 5684 6205 5718 6211
rect 5684 6177 5718 6205
rect 5684 6137 5718 6139
rect 5684 6105 5718 6137
rect 5684 6035 5718 6067
rect 5684 6033 5718 6035
rect 5684 5967 5718 5995
rect 5684 5961 5718 5967
rect 5684 5899 5718 5923
rect 5684 5889 5718 5899
rect 5684 5831 5718 5851
rect 5684 5817 5718 5831
rect 5684 5763 5718 5779
rect 5684 5745 5718 5763
rect 5684 5695 5718 5707
rect 5684 5673 5718 5695
rect 5684 5627 5718 5635
rect 5684 5601 5718 5627
rect 10568 6774 10762 6878
rect 12994 6814 13028 6848
rect 11514 6736 11548 6770
rect 11802 6751 11836 6785
rect 12518 6729 12552 6763
rect 6180 6549 6214 6575
rect 6180 6541 6214 6549
rect 6180 6481 6214 6503
rect 6180 6469 6214 6481
rect 6180 6413 6214 6431
rect 6180 6397 6214 6413
rect 6180 6345 6214 6359
rect 6180 6325 6214 6345
rect 6180 6277 6214 6287
rect 6180 6253 6214 6277
rect 6180 6209 6214 6215
rect 6180 6181 6214 6209
rect 6180 6141 6214 6143
rect 6180 6109 6214 6141
rect 6180 6039 6214 6071
rect 6180 6037 6214 6039
rect 6180 5971 6214 5999
rect 6180 5965 6214 5971
rect 6180 5903 6214 5927
rect 6180 5893 6214 5903
rect 6180 5835 6214 5855
rect 6180 5821 6214 5835
rect 6180 5767 6214 5783
rect 6180 5749 6214 5767
rect 6180 5699 6214 5711
rect 6180 5677 6214 5699
rect 6180 5631 6214 5639
rect 6180 5605 6214 5631
rect 6276 6549 6310 6575
rect 6276 6541 6310 6549
rect 6276 6481 6310 6503
rect 6276 6469 6310 6481
rect 6276 6413 6310 6431
rect 6276 6397 6310 6413
rect 6276 6345 6310 6359
rect 6276 6325 6310 6345
rect 6276 6277 6310 6287
rect 6276 6253 6310 6277
rect 6276 6209 6310 6215
rect 6276 6181 6310 6209
rect 6276 6141 6310 6143
rect 6276 6109 6310 6141
rect 6276 6039 6310 6071
rect 6276 6037 6310 6039
rect 6276 5971 6310 5999
rect 6276 5965 6310 5971
rect 6276 5903 6310 5927
rect 6276 5893 6310 5903
rect 6276 5835 6310 5855
rect 6276 5821 6310 5835
rect 6276 5767 6310 5783
rect 6276 5749 6310 5767
rect 6276 5699 6310 5711
rect 6276 5677 6310 5699
rect 6276 5631 6310 5639
rect 6276 5605 6310 5631
rect 2278 5372 2380 5418
rect 6372 6549 6406 6575
rect 6372 6541 6406 6549
rect 6372 6481 6406 6503
rect 6372 6469 6406 6481
rect 6372 6413 6406 6431
rect 6372 6397 6406 6413
rect 6372 6345 6406 6359
rect 6372 6325 6406 6345
rect 6372 6277 6406 6287
rect 6372 6253 6406 6277
rect 6372 6209 6406 6215
rect 6372 6181 6406 6209
rect 6372 6141 6406 6143
rect 6372 6109 6406 6141
rect 6372 6039 6406 6071
rect 6372 6037 6406 6039
rect 6372 5971 6406 5999
rect 6372 5965 6406 5971
rect 6372 5903 6406 5927
rect 6372 5893 6406 5903
rect 6372 5835 6406 5855
rect 6372 5821 6406 5835
rect 6372 5767 6406 5783
rect 6372 5749 6406 5767
rect 6372 5699 6406 5711
rect 6372 5677 6406 5699
rect 6372 5631 6406 5639
rect 6372 5605 6406 5631
rect 6468 6549 6502 6575
rect 6468 6541 6502 6549
rect 6468 6481 6502 6503
rect 6468 6469 6502 6481
rect 6468 6413 6502 6431
rect 6468 6397 6502 6413
rect 6468 6345 6502 6359
rect 6468 6325 6502 6345
rect 6468 6277 6502 6287
rect 6468 6253 6502 6277
rect 6468 6209 6502 6215
rect 6468 6181 6502 6209
rect 6468 6141 6502 6143
rect 6468 6109 6502 6141
rect 6468 6039 6502 6071
rect 6468 6037 6502 6039
rect 6468 5971 6502 5999
rect 6468 5965 6502 5971
rect 6468 5903 6502 5927
rect 6468 5893 6502 5903
rect 6468 5835 6502 5855
rect 6468 5821 6502 5835
rect 6468 5767 6502 5783
rect 6468 5749 6502 5767
rect 6468 5699 6502 5711
rect 6468 5677 6502 5699
rect 6468 5631 6502 5639
rect 6468 5605 6502 5631
rect 6564 6549 6598 6575
rect 6564 6541 6598 6549
rect 6564 6481 6598 6503
rect 6564 6469 6598 6481
rect 6564 6413 6598 6431
rect 6564 6397 6598 6413
rect 6564 6345 6598 6359
rect 6564 6325 6598 6345
rect 6564 6277 6598 6287
rect 6564 6253 6598 6277
rect 6564 6209 6598 6215
rect 6564 6181 6598 6209
rect 6564 6141 6598 6143
rect 6564 6109 6598 6141
rect 6564 6039 6598 6071
rect 6564 6037 6598 6039
rect 6564 5971 6598 5999
rect 6564 5965 6598 5971
rect 6564 5903 6598 5927
rect 6564 5893 6598 5903
rect 6564 5835 6598 5855
rect 6564 5821 6598 5835
rect 6564 5767 6598 5783
rect 6564 5749 6598 5767
rect 6564 5699 6598 5711
rect 6564 5677 6598 5699
rect 6564 5631 6598 5639
rect 6564 5605 6598 5631
rect 6660 6549 6694 6575
rect 6660 6541 6694 6549
rect 6660 6481 6694 6503
rect 6660 6469 6694 6481
rect 6660 6413 6694 6431
rect 6660 6397 6694 6413
rect 6660 6345 6694 6359
rect 6660 6325 6694 6345
rect 6660 6277 6694 6287
rect 6660 6253 6694 6277
rect 6660 6209 6694 6215
rect 6660 6181 6694 6209
rect 6660 6141 6694 6143
rect 6660 6109 6694 6141
rect 6660 6039 6694 6071
rect 6660 6037 6694 6039
rect 6660 5971 6694 5999
rect 6660 5965 6694 5971
rect 6660 5903 6694 5927
rect 6660 5893 6694 5903
rect 6660 5835 6694 5855
rect 6660 5821 6694 5835
rect 6660 5767 6694 5783
rect 6660 5749 6694 5767
rect 6660 5699 6694 5711
rect 6660 5677 6694 5699
rect 6660 5631 6694 5639
rect 6660 5605 6694 5631
rect 6756 6549 6790 6575
rect 6756 6541 6790 6549
rect 6756 6481 6790 6503
rect 6756 6469 6790 6481
rect 6756 6413 6790 6431
rect 6756 6397 6790 6413
rect 6756 6345 6790 6359
rect 6756 6325 6790 6345
rect 6756 6277 6790 6287
rect 6756 6253 6790 6277
rect 6756 6209 6790 6215
rect 6756 6181 6790 6209
rect 6756 6141 6790 6143
rect 6756 6109 6790 6141
rect 6756 6039 6790 6071
rect 6756 6037 6790 6039
rect 6756 5971 6790 5999
rect 6756 5965 6790 5971
rect 6756 5903 6790 5927
rect 6756 5893 6790 5903
rect 6756 5835 6790 5855
rect 6756 5821 6790 5835
rect 6756 5767 6790 5783
rect 6756 5749 6790 5767
rect 6756 5699 6790 5711
rect 6756 5677 6790 5699
rect 6756 5631 6790 5639
rect 6756 5605 6790 5631
rect 6852 6549 6886 6575
rect 6852 6541 6886 6549
rect 6852 6481 6886 6503
rect 6852 6469 6886 6481
rect 6852 6413 6886 6431
rect 6852 6397 6886 6413
rect 6852 6345 6886 6359
rect 6852 6325 6886 6345
rect 6852 6277 6886 6287
rect 6852 6253 6886 6277
rect 6852 6209 6886 6215
rect 6852 6181 6886 6209
rect 6852 6141 6886 6143
rect 6852 6109 6886 6141
rect 6852 6039 6886 6071
rect 6852 6037 6886 6039
rect 6852 5971 6886 5999
rect 6852 5965 6886 5971
rect 6852 5903 6886 5927
rect 6852 5893 6886 5903
rect 6852 5835 6886 5855
rect 6852 5821 6886 5835
rect 6852 5767 6886 5783
rect 6852 5749 6886 5767
rect 6852 5699 6886 5711
rect 6852 5677 6886 5699
rect 6852 5631 6886 5639
rect 6852 5605 6886 5631
rect 6948 6549 6982 6575
rect 6948 6541 6982 6549
rect 6948 6481 6982 6503
rect 6948 6469 6982 6481
rect 6948 6413 6982 6431
rect 6948 6397 6982 6413
rect 6948 6345 6982 6359
rect 6948 6325 6982 6345
rect 6948 6277 6982 6287
rect 6948 6253 6982 6277
rect 6948 6209 6982 6215
rect 6948 6181 6982 6209
rect 6948 6141 6982 6143
rect 6948 6109 6982 6141
rect 6948 6039 6982 6071
rect 6948 6037 6982 6039
rect 6948 5971 6982 5999
rect 6948 5965 6982 5971
rect 6948 5903 6982 5927
rect 6948 5893 6982 5903
rect 6948 5835 6982 5855
rect 6948 5821 6982 5835
rect 6948 5767 6982 5783
rect 6948 5749 6982 5767
rect 6948 5699 6982 5711
rect 6948 5677 6982 5699
rect 6948 5631 6982 5639
rect 6948 5605 6982 5631
rect 7044 6549 7078 6575
rect 7044 6541 7078 6549
rect 7044 6481 7078 6503
rect 7044 6469 7078 6481
rect 7044 6413 7078 6431
rect 7044 6397 7078 6413
rect 7044 6345 7078 6359
rect 7044 6325 7078 6345
rect 7044 6277 7078 6287
rect 7044 6253 7078 6277
rect 7044 6209 7078 6215
rect 7044 6181 7078 6209
rect 7044 6141 7078 6143
rect 7044 6109 7078 6141
rect 7044 6039 7078 6071
rect 7044 6037 7078 6039
rect 7044 5971 7078 5999
rect 7044 5965 7078 5971
rect 7044 5903 7078 5927
rect 7044 5893 7078 5903
rect 7044 5835 7078 5855
rect 7044 5821 7078 5835
rect 7044 5767 7078 5783
rect 7044 5749 7078 5767
rect 7044 5699 7078 5711
rect 7044 5677 7078 5699
rect 7044 5631 7078 5639
rect 7044 5605 7078 5631
rect 7140 6549 7174 6575
rect 7140 6541 7174 6549
rect 7140 6481 7174 6503
rect 7140 6469 7174 6481
rect 7140 6413 7174 6431
rect 7140 6397 7174 6413
rect 7140 6345 7174 6359
rect 7140 6325 7174 6345
rect 7140 6277 7174 6287
rect 7140 6253 7174 6277
rect 7140 6209 7174 6215
rect 7140 6181 7174 6209
rect 7140 6141 7174 6143
rect 7140 6109 7174 6141
rect 7140 6039 7174 6071
rect 7140 6037 7174 6039
rect 7140 5971 7174 5999
rect 7140 5965 7174 5971
rect 7140 5903 7174 5927
rect 7140 5893 7174 5903
rect 7140 5835 7174 5855
rect 7140 5821 7174 5835
rect 7140 5767 7174 5783
rect 7140 5749 7174 5767
rect 7140 5699 7174 5711
rect 7140 5677 7174 5699
rect 7140 5631 7174 5639
rect 7140 5605 7174 5631
rect 7236 6549 7270 6575
rect 7236 6541 7270 6549
rect 7236 6481 7270 6503
rect 7236 6469 7270 6481
rect 7236 6413 7270 6431
rect 7236 6397 7270 6413
rect 7236 6345 7270 6359
rect 7236 6325 7270 6345
rect 7236 6277 7270 6287
rect 7236 6253 7270 6277
rect 7236 6209 7270 6215
rect 7236 6181 7270 6209
rect 7236 6141 7270 6143
rect 7236 6109 7270 6141
rect 7236 6039 7270 6071
rect 7236 6037 7270 6039
rect 7236 5971 7270 5999
rect 7236 5965 7270 5971
rect 7236 5903 7270 5927
rect 7236 5893 7270 5903
rect 7236 5835 7270 5855
rect 7236 5821 7270 5835
rect 7236 5767 7270 5783
rect 7236 5749 7270 5767
rect 7236 5699 7270 5711
rect 7236 5677 7270 5699
rect 7236 5631 7270 5639
rect 7236 5605 7270 5631
rect 7332 6549 7366 6575
rect 7332 6541 7366 6549
rect 7332 6481 7366 6503
rect 7332 6469 7366 6481
rect 7332 6413 7366 6431
rect 7332 6397 7366 6413
rect 7332 6345 7366 6359
rect 7332 6325 7366 6345
rect 7332 6277 7366 6287
rect 7332 6253 7366 6277
rect 7332 6209 7366 6215
rect 7332 6181 7366 6209
rect 7332 6141 7366 6143
rect 7332 6109 7366 6141
rect 7332 6039 7366 6071
rect 7332 6037 7366 6039
rect 7332 5971 7366 5999
rect 7332 5965 7366 5971
rect 7332 5903 7366 5927
rect 7332 5893 7366 5903
rect 7332 5835 7366 5855
rect 7332 5821 7366 5835
rect 7332 5767 7366 5783
rect 7332 5749 7366 5767
rect 7332 5699 7366 5711
rect 7332 5677 7366 5699
rect 7332 5631 7366 5639
rect 7332 5605 7366 5631
rect 7946 6545 7980 6571
rect 7946 6537 7980 6545
rect 7946 6477 7980 6499
rect 7946 6465 7980 6477
rect 7946 6409 7980 6427
rect 7946 6393 7980 6409
rect 7946 6341 7980 6355
rect 7946 6321 7980 6341
rect 7946 6273 7980 6283
rect 7946 6249 7980 6273
rect 7946 6205 7980 6211
rect 7946 6177 7980 6205
rect 7946 6137 7980 6139
rect 7946 6105 7980 6137
rect 7946 6035 7980 6067
rect 7946 6033 7980 6035
rect 7946 5967 7980 5995
rect 7946 5961 7980 5967
rect 7946 5899 7980 5923
rect 7946 5889 7980 5899
rect 7946 5831 7980 5851
rect 7946 5817 7980 5831
rect 7946 5763 7980 5779
rect 7946 5745 7980 5763
rect 7946 5695 7980 5707
rect 7946 5673 7980 5695
rect 7946 5627 7980 5635
rect 7946 5601 7980 5627
rect 8042 6545 8076 6571
rect 8042 6537 8076 6545
rect 8042 6477 8076 6499
rect 8042 6465 8076 6477
rect 8042 6409 8076 6427
rect 8042 6393 8076 6409
rect 8042 6341 8076 6355
rect 8042 6321 8076 6341
rect 8042 6273 8076 6283
rect 8042 6249 8076 6273
rect 8042 6205 8076 6211
rect 8042 6177 8076 6205
rect 8042 6137 8076 6139
rect 8042 6105 8076 6137
rect 8042 6035 8076 6067
rect 8042 6033 8076 6035
rect 8042 5967 8076 5995
rect 8042 5961 8076 5967
rect 8042 5899 8076 5923
rect 8042 5889 8076 5899
rect 8042 5831 8076 5851
rect 8042 5817 8076 5831
rect 8042 5763 8076 5779
rect 8042 5745 8076 5763
rect 8042 5695 8076 5707
rect 8042 5673 8076 5695
rect 8042 5627 8076 5635
rect 8042 5601 8076 5627
rect 8138 6545 8172 6571
rect 8138 6537 8172 6545
rect 8138 6477 8172 6499
rect 8138 6465 8172 6477
rect 8138 6409 8172 6427
rect 8138 6393 8172 6409
rect 8138 6341 8172 6355
rect 8138 6321 8172 6341
rect 8138 6273 8172 6283
rect 8138 6249 8172 6273
rect 8138 6205 8172 6211
rect 8138 6177 8172 6205
rect 8138 6137 8172 6139
rect 8138 6105 8172 6137
rect 8138 6035 8172 6067
rect 8138 6033 8172 6035
rect 8138 5967 8172 5995
rect 8138 5961 8172 5967
rect 8138 5899 8172 5923
rect 8138 5889 8172 5899
rect 8138 5831 8172 5851
rect 8138 5817 8172 5831
rect 8138 5763 8172 5779
rect 8138 5745 8172 5763
rect 8138 5695 8172 5707
rect 8138 5673 8172 5695
rect 8138 5627 8172 5635
rect 8138 5601 8172 5627
rect 8234 6545 8268 6571
rect 8234 6537 8268 6545
rect 8234 6477 8268 6499
rect 8234 6465 8268 6477
rect 8234 6409 8268 6427
rect 8234 6393 8268 6409
rect 8234 6341 8268 6355
rect 8234 6321 8268 6341
rect 8234 6273 8268 6283
rect 8234 6249 8268 6273
rect 8234 6205 8268 6211
rect 8234 6177 8268 6205
rect 8234 6137 8268 6139
rect 8234 6105 8268 6137
rect 8234 6035 8268 6067
rect 8234 6033 8268 6035
rect 8234 5967 8268 5995
rect 8234 5961 8268 5967
rect 8234 5899 8268 5923
rect 8234 5889 8268 5899
rect 8234 5831 8268 5851
rect 8234 5817 8268 5831
rect 8234 5763 8268 5779
rect 8234 5745 8268 5763
rect 8234 5695 8268 5707
rect 8234 5673 8268 5695
rect 8234 5627 8268 5635
rect 8234 5601 8268 5627
rect 8330 6545 8364 6571
rect 8330 6537 8364 6545
rect 8330 6477 8364 6499
rect 8330 6465 8364 6477
rect 8330 6409 8364 6427
rect 8330 6393 8364 6409
rect 8330 6341 8364 6355
rect 8330 6321 8364 6341
rect 8330 6273 8364 6283
rect 8330 6249 8364 6273
rect 8330 6205 8364 6211
rect 8330 6177 8364 6205
rect 8330 6137 8364 6139
rect 8330 6105 8364 6137
rect 8330 6035 8364 6067
rect 8330 6033 8364 6035
rect 8330 5967 8364 5995
rect 8330 5961 8364 5967
rect 8330 5899 8364 5923
rect 8330 5889 8364 5899
rect 8330 5831 8364 5851
rect 8330 5817 8364 5831
rect 8330 5763 8364 5779
rect 8330 5745 8364 5763
rect 8330 5695 8364 5707
rect 8330 5673 8364 5695
rect 8330 5627 8364 5635
rect 8330 5601 8364 5627
rect 8426 6545 8460 6571
rect 8426 6537 8460 6545
rect 8426 6477 8460 6499
rect 8426 6465 8460 6477
rect 8426 6409 8460 6427
rect 8426 6393 8460 6409
rect 8426 6341 8460 6355
rect 8426 6321 8460 6341
rect 8426 6273 8460 6283
rect 8426 6249 8460 6273
rect 8426 6205 8460 6211
rect 8426 6177 8460 6205
rect 8426 6137 8460 6139
rect 8426 6105 8460 6137
rect 8426 6035 8460 6067
rect 8426 6033 8460 6035
rect 8426 5967 8460 5995
rect 8426 5961 8460 5967
rect 8426 5899 8460 5923
rect 8426 5889 8460 5899
rect 8426 5831 8460 5851
rect 8426 5817 8460 5831
rect 8426 5763 8460 5779
rect 8426 5745 8460 5763
rect 8426 5695 8460 5707
rect 8426 5673 8460 5695
rect 8426 5627 8460 5635
rect 8426 5601 8460 5627
rect 8522 6545 8556 6571
rect 8522 6537 8556 6545
rect 8522 6477 8556 6499
rect 8522 6465 8556 6477
rect 8522 6409 8556 6427
rect 8522 6393 8556 6409
rect 8522 6341 8556 6355
rect 8522 6321 8556 6341
rect 8522 6273 8556 6283
rect 8522 6249 8556 6273
rect 8522 6205 8556 6211
rect 8522 6177 8556 6205
rect 8522 6137 8556 6139
rect 8522 6105 8556 6137
rect 8522 6035 8556 6067
rect 8522 6033 8556 6035
rect 8522 5967 8556 5995
rect 8522 5961 8556 5967
rect 8522 5899 8556 5923
rect 8522 5889 8556 5899
rect 8522 5831 8556 5851
rect 8522 5817 8556 5831
rect 8522 5763 8556 5779
rect 8522 5745 8556 5763
rect 8522 5695 8556 5707
rect 8522 5673 8556 5695
rect 8522 5627 8556 5635
rect 8522 5601 8556 5627
rect 8618 6545 8652 6571
rect 8618 6537 8652 6545
rect 8618 6477 8652 6499
rect 8618 6465 8652 6477
rect 8618 6409 8652 6427
rect 8618 6393 8652 6409
rect 8618 6341 8652 6355
rect 8618 6321 8652 6341
rect 8618 6273 8652 6283
rect 8618 6249 8652 6273
rect 8618 6205 8652 6211
rect 8618 6177 8652 6205
rect 8618 6137 8652 6139
rect 8618 6105 8652 6137
rect 8618 6035 8652 6067
rect 8618 6033 8652 6035
rect 8618 5967 8652 5995
rect 8618 5961 8652 5967
rect 8618 5899 8652 5923
rect 8618 5889 8652 5899
rect 8618 5831 8652 5851
rect 8618 5817 8652 5831
rect 8618 5763 8652 5779
rect 8618 5745 8652 5763
rect 8618 5695 8652 5707
rect 8618 5673 8652 5695
rect 8618 5627 8652 5635
rect 8618 5601 8652 5627
rect 8714 6545 8748 6571
rect 8714 6537 8748 6545
rect 8714 6477 8748 6499
rect 8714 6465 8748 6477
rect 8714 6409 8748 6427
rect 8714 6393 8748 6409
rect 8714 6341 8748 6355
rect 8714 6321 8748 6341
rect 8714 6273 8748 6283
rect 8714 6249 8748 6273
rect 8714 6205 8748 6211
rect 8714 6177 8748 6205
rect 8714 6137 8748 6139
rect 8714 6105 8748 6137
rect 8714 6035 8748 6067
rect 8714 6033 8748 6035
rect 8714 5967 8748 5995
rect 8714 5961 8748 5967
rect 8714 5899 8748 5923
rect 8714 5889 8748 5899
rect 8714 5831 8748 5851
rect 8714 5817 8748 5831
rect 8714 5763 8748 5779
rect 8714 5745 8748 5763
rect 8714 5695 8748 5707
rect 8714 5673 8748 5695
rect 8714 5627 8748 5635
rect 8714 5601 8748 5627
rect 13724 6748 13918 6852
rect 14670 6710 14704 6744
rect 14958 6725 14992 6759
rect 9268 6547 9302 6573
rect 9268 6539 9302 6547
rect 9268 6479 9302 6501
rect 9268 6467 9302 6479
rect 9268 6411 9302 6429
rect 9268 6395 9302 6411
rect 9268 6343 9302 6357
rect 9268 6323 9302 6343
rect 9268 6275 9302 6285
rect 9268 6251 9302 6275
rect 9268 6207 9302 6213
rect 9268 6179 9302 6207
rect 9268 6139 9302 6141
rect 9268 6107 9302 6139
rect 9268 6037 9302 6069
rect 9268 6035 9302 6037
rect 9268 5969 9302 5997
rect 9268 5963 9302 5969
rect 9268 5901 9302 5925
rect 9268 5891 9302 5901
rect 9268 5833 9302 5853
rect 9268 5819 9302 5833
rect 9268 5765 9302 5781
rect 9268 5747 9302 5765
rect 9268 5697 9302 5709
rect 9268 5675 9302 5697
rect 9268 5629 9302 5637
rect 9268 5603 9302 5629
rect 9364 6547 9398 6573
rect 9364 6539 9398 6547
rect 9364 6479 9398 6501
rect 9364 6467 9398 6479
rect 9364 6411 9398 6429
rect 9364 6395 9398 6411
rect 9364 6343 9398 6357
rect 9364 6323 9398 6343
rect 9364 6275 9398 6285
rect 9364 6251 9398 6275
rect 9364 6207 9398 6213
rect 9364 6179 9398 6207
rect 9364 6139 9398 6141
rect 9364 6107 9398 6139
rect 9364 6037 9398 6069
rect 9364 6035 9398 6037
rect 9364 5969 9398 5997
rect 9364 5963 9398 5969
rect 9364 5901 9398 5925
rect 9364 5891 9398 5901
rect 9364 5833 9398 5853
rect 9364 5819 9398 5833
rect 9364 5765 9398 5781
rect 9364 5747 9398 5765
rect 9364 5697 9398 5709
rect 9364 5675 9398 5697
rect 9364 5629 9398 5637
rect 9364 5603 9398 5629
rect 3824 5354 3926 5400
rect -868 5317 -834 5345
rect 5234 5352 5336 5398
rect 9460 6547 9494 6573
rect 9460 6539 9494 6547
rect 9460 6479 9494 6501
rect 9460 6467 9494 6479
rect 9460 6411 9494 6429
rect 9460 6395 9494 6411
rect 9460 6343 9494 6357
rect 9460 6323 9494 6343
rect 9460 6275 9494 6285
rect 9460 6251 9494 6275
rect 9460 6207 9494 6213
rect 9460 6179 9494 6207
rect 9460 6139 9494 6141
rect 9460 6107 9494 6139
rect 9460 6037 9494 6069
rect 9460 6035 9494 6037
rect 9460 5969 9494 5997
rect 9460 5963 9494 5969
rect 9460 5901 9494 5925
rect 9460 5891 9494 5901
rect 9460 5833 9494 5853
rect 9460 5819 9494 5833
rect 9460 5765 9494 5781
rect 9460 5747 9494 5765
rect 9460 5697 9494 5709
rect 9460 5675 9494 5697
rect 9460 5629 9494 5637
rect 9460 5603 9494 5629
rect 9556 6547 9590 6573
rect 9556 6539 9590 6547
rect 9556 6479 9590 6501
rect 9556 6467 9590 6479
rect 9556 6411 9590 6429
rect 9556 6395 9590 6411
rect 9556 6343 9590 6357
rect 9556 6323 9590 6343
rect 9556 6275 9590 6285
rect 9556 6251 9590 6275
rect 9556 6207 9590 6213
rect 9556 6179 9590 6207
rect 9556 6139 9590 6141
rect 9556 6107 9590 6139
rect 9556 6037 9590 6069
rect 9556 6035 9590 6037
rect 9556 5969 9590 5997
rect 9556 5963 9590 5969
rect 9556 5901 9590 5925
rect 9556 5891 9590 5901
rect 9556 5833 9590 5853
rect 9556 5819 9590 5833
rect 9556 5765 9590 5781
rect 9556 5747 9590 5765
rect 9556 5697 9590 5709
rect 9556 5675 9590 5697
rect 9556 5629 9590 5637
rect 9556 5603 9590 5629
rect 9652 6547 9686 6573
rect 9652 6539 9686 6547
rect 9652 6479 9686 6501
rect 9652 6467 9686 6479
rect 9652 6411 9686 6429
rect 9652 6395 9686 6411
rect 9652 6343 9686 6357
rect 9652 6323 9686 6343
rect 9652 6275 9686 6285
rect 9652 6251 9686 6275
rect 9652 6207 9686 6213
rect 9652 6179 9686 6207
rect 9652 6139 9686 6141
rect 9652 6107 9686 6139
rect 9652 6037 9686 6069
rect 9652 6035 9686 6037
rect 9652 5969 9686 5997
rect 9652 5963 9686 5969
rect 9652 5901 9686 5925
rect 9652 5891 9686 5901
rect 9652 5833 9686 5853
rect 9652 5819 9686 5833
rect 9652 5765 9686 5781
rect 9652 5747 9686 5765
rect 9652 5697 9686 5709
rect 9652 5675 9686 5697
rect 9652 5629 9686 5637
rect 9652 5603 9686 5629
rect 9748 6547 9782 6573
rect 9748 6539 9782 6547
rect 9748 6479 9782 6501
rect 9748 6467 9782 6479
rect 9748 6411 9782 6429
rect 9748 6395 9782 6411
rect 9748 6343 9782 6357
rect 9748 6323 9782 6343
rect 9748 6275 9782 6285
rect 9748 6251 9782 6275
rect 9748 6207 9782 6213
rect 9748 6179 9782 6207
rect 9748 6139 9782 6141
rect 9748 6107 9782 6139
rect 9748 6037 9782 6069
rect 9748 6035 9782 6037
rect 9748 5969 9782 5997
rect 9748 5963 9782 5969
rect 9748 5901 9782 5925
rect 9748 5891 9782 5901
rect 9748 5833 9782 5853
rect 9748 5819 9782 5833
rect 9748 5765 9782 5781
rect 9748 5747 9782 5765
rect 9748 5697 9782 5709
rect 9748 5675 9782 5697
rect 9748 5629 9782 5637
rect 9748 5603 9782 5629
rect 9844 6547 9878 6573
rect 9844 6539 9878 6547
rect 9844 6479 9878 6501
rect 9844 6467 9878 6479
rect 9844 6411 9878 6429
rect 9844 6395 9878 6411
rect 9844 6343 9878 6357
rect 9844 6323 9878 6343
rect 9844 6275 9878 6285
rect 9844 6251 9878 6275
rect 9844 6207 9878 6213
rect 9844 6179 9878 6207
rect 9844 6139 9878 6141
rect 9844 6107 9878 6139
rect 9844 6037 9878 6069
rect 9844 6035 9878 6037
rect 9844 5969 9878 5997
rect 9844 5963 9878 5969
rect 9844 5901 9878 5925
rect 9844 5891 9878 5901
rect 9844 5833 9878 5853
rect 9844 5819 9878 5833
rect 9844 5765 9878 5781
rect 9844 5747 9878 5765
rect 9844 5697 9878 5709
rect 9844 5675 9878 5697
rect 9844 5629 9878 5637
rect 9844 5603 9878 5629
rect 9940 6547 9974 6573
rect 9940 6539 9974 6547
rect 9940 6479 9974 6501
rect 9940 6467 9974 6479
rect 9940 6411 9974 6429
rect 9940 6395 9974 6411
rect 9940 6343 9974 6357
rect 9940 6323 9974 6343
rect 9940 6275 9974 6285
rect 9940 6251 9974 6275
rect 9940 6207 9974 6213
rect 9940 6179 9974 6207
rect 9940 6139 9974 6141
rect 9940 6107 9974 6139
rect 9940 6037 9974 6069
rect 9940 6035 9974 6037
rect 9940 5969 9974 5997
rect 9940 5963 9974 5969
rect 9940 5901 9974 5925
rect 9940 5891 9974 5901
rect 9940 5833 9974 5853
rect 9940 5819 9974 5833
rect 9940 5765 9974 5781
rect 9940 5747 9974 5765
rect 9940 5697 9974 5709
rect 9940 5675 9974 5697
rect 9940 5629 9974 5637
rect 9940 5603 9974 5629
rect 10036 6547 10070 6573
rect 10036 6539 10070 6547
rect 10036 6479 10070 6501
rect 10036 6467 10070 6479
rect 10036 6411 10070 6429
rect 10036 6395 10070 6411
rect 10036 6343 10070 6357
rect 10036 6323 10070 6343
rect 10036 6275 10070 6285
rect 10036 6251 10070 6275
rect 10036 6207 10070 6213
rect 10036 6179 10070 6207
rect 10036 6139 10070 6141
rect 10036 6107 10070 6139
rect 10036 6037 10070 6069
rect 10036 6035 10070 6037
rect 10036 5969 10070 5997
rect 10036 5963 10070 5969
rect 10036 5901 10070 5925
rect 10036 5891 10070 5901
rect 10036 5833 10070 5853
rect 10036 5819 10070 5833
rect 10036 5765 10070 5781
rect 10036 5747 10070 5765
rect 10036 5697 10070 5709
rect 10036 5675 10070 5697
rect 10036 5629 10070 5637
rect 10036 5603 10070 5629
rect 10132 6547 10166 6573
rect 10132 6539 10166 6547
rect 10132 6479 10166 6501
rect 10132 6467 10166 6479
rect 10132 6411 10166 6429
rect 10132 6395 10166 6411
rect 10132 6343 10166 6357
rect 10132 6323 10166 6343
rect 10132 6275 10166 6285
rect 10132 6251 10166 6275
rect 10132 6207 10166 6213
rect 10132 6179 10166 6207
rect 10132 6139 10166 6141
rect 10132 6107 10166 6139
rect 10132 6037 10166 6069
rect 10132 6035 10166 6037
rect 10132 5969 10166 5997
rect 10132 5963 10166 5969
rect 10132 5901 10166 5925
rect 10132 5891 10166 5901
rect 10132 5833 10166 5853
rect 10132 5819 10166 5833
rect 10132 5765 10166 5781
rect 10132 5747 10166 5765
rect 10132 5697 10166 5709
rect 10132 5675 10166 5697
rect 10132 5629 10166 5637
rect 10132 5603 10166 5629
rect 10228 6547 10262 6573
rect 10228 6539 10262 6547
rect 10228 6479 10262 6501
rect 10228 6467 10262 6479
rect 10228 6411 10262 6429
rect 10228 6395 10262 6411
rect 10228 6343 10262 6357
rect 10228 6323 10262 6343
rect 10228 6275 10262 6285
rect 10228 6251 10262 6275
rect 10228 6207 10262 6213
rect 10228 6179 10262 6207
rect 10228 6139 10262 6141
rect 10228 6107 10262 6139
rect 10228 6037 10262 6069
rect 10228 6035 10262 6037
rect 10228 5969 10262 5997
rect 10228 5963 10262 5969
rect 10228 5901 10262 5925
rect 10228 5891 10262 5901
rect 10228 5833 10262 5853
rect 10228 5819 10262 5833
rect 10228 5765 10262 5781
rect 10228 5747 10262 5765
rect 10228 5697 10262 5709
rect 10228 5675 10262 5697
rect 10228 5629 10262 5637
rect 10228 5603 10262 5629
rect 10324 6547 10358 6573
rect 10324 6539 10358 6547
rect 10324 6479 10358 6501
rect 10324 6467 10358 6479
rect 10324 6411 10358 6429
rect 10324 6395 10358 6411
rect 10324 6343 10358 6357
rect 10324 6323 10358 6343
rect 10324 6275 10358 6285
rect 10324 6251 10358 6275
rect 10324 6207 10358 6213
rect 10324 6179 10358 6207
rect 10324 6139 10358 6141
rect 10324 6107 10358 6139
rect 10324 6037 10358 6069
rect 10324 6035 10358 6037
rect 10324 5969 10358 5997
rect 10324 5963 10358 5969
rect 10324 5901 10358 5925
rect 10324 5891 10358 5901
rect 10324 5833 10358 5853
rect 10324 5819 10358 5833
rect 10324 5765 10358 5781
rect 10324 5747 10358 5765
rect 10324 5697 10358 5709
rect 10324 5675 10358 5697
rect 10324 5629 10358 5637
rect 10324 5603 10358 5629
rect 10420 6547 10454 6573
rect 10420 6539 10454 6547
rect 10420 6479 10454 6501
rect 10420 6467 10454 6479
rect 10420 6411 10454 6429
rect 10420 6395 10454 6411
rect 10420 6343 10454 6357
rect 10420 6323 10454 6343
rect 10420 6275 10454 6285
rect 10420 6251 10454 6275
rect 10420 6207 10454 6213
rect 10420 6179 10454 6207
rect 10420 6139 10454 6141
rect 10420 6107 10454 6139
rect 10420 6037 10454 6069
rect 10420 6035 10454 6037
rect 10420 5969 10454 5997
rect 10420 5963 10454 5969
rect 10420 5901 10454 5925
rect 10420 5891 10454 5901
rect 10420 5833 10454 5853
rect 10420 5819 10454 5833
rect 10420 5765 10454 5781
rect 10420 5747 10454 5765
rect 10420 5697 10454 5709
rect 10420 5675 10454 5697
rect 10420 5629 10454 5637
rect 10420 5603 10454 5629
rect 11034 6543 11068 6569
rect 11034 6535 11068 6543
rect 11034 6475 11068 6497
rect 11034 6463 11068 6475
rect 11034 6407 11068 6425
rect 11034 6391 11068 6407
rect 11034 6339 11068 6353
rect 11034 6319 11068 6339
rect 11034 6271 11068 6281
rect 11034 6247 11068 6271
rect 11034 6203 11068 6209
rect 11034 6175 11068 6203
rect 11034 6135 11068 6137
rect 11034 6103 11068 6135
rect 11034 6033 11068 6065
rect 11034 6031 11068 6033
rect 11034 5965 11068 5993
rect 11034 5959 11068 5965
rect 11034 5897 11068 5921
rect 11034 5887 11068 5897
rect 11034 5829 11068 5849
rect 11034 5815 11068 5829
rect 11034 5761 11068 5777
rect 11034 5743 11068 5761
rect 11034 5693 11068 5705
rect 11034 5671 11068 5693
rect 11034 5625 11068 5633
rect 11034 5599 11068 5625
rect 11130 6543 11164 6569
rect 11130 6535 11164 6543
rect 11130 6475 11164 6497
rect 11130 6463 11164 6475
rect 11130 6407 11164 6425
rect 11130 6391 11164 6407
rect 11130 6339 11164 6353
rect 11130 6319 11164 6339
rect 11130 6271 11164 6281
rect 11130 6247 11164 6271
rect 11130 6203 11164 6209
rect 11130 6175 11164 6203
rect 11130 6135 11164 6137
rect 11130 6103 11164 6135
rect 11130 6033 11164 6065
rect 11130 6031 11164 6033
rect 11130 5965 11164 5993
rect 11130 5959 11164 5965
rect 11130 5897 11164 5921
rect 11130 5887 11164 5897
rect 11130 5829 11164 5849
rect 11130 5815 11164 5829
rect 11130 5761 11164 5777
rect 11130 5743 11164 5761
rect 11130 5693 11164 5705
rect 11130 5671 11164 5693
rect 11130 5625 11164 5633
rect 11130 5599 11164 5625
rect 11226 6543 11260 6569
rect 11226 6535 11260 6543
rect 11226 6475 11260 6497
rect 11226 6463 11260 6475
rect 11226 6407 11260 6425
rect 11226 6391 11260 6407
rect 11226 6339 11260 6353
rect 11226 6319 11260 6339
rect 11226 6271 11260 6281
rect 11226 6247 11260 6271
rect 11226 6203 11260 6209
rect 11226 6175 11260 6203
rect 11226 6135 11260 6137
rect 11226 6103 11260 6135
rect 11226 6033 11260 6065
rect 11226 6031 11260 6033
rect 11226 5965 11260 5993
rect 11226 5959 11260 5965
rect 11226 5897 11260 5921
rect 11226 5887 11260 5897
rect 11226 5829 11260 5849
rect 11226 5815 11260 5829
rect 11226 5761 11260 5777
rect 11226 5743 11260 5761
rect 11226 5693 11260 5705
rect 11226 5671 11260 5693
rect 11226 5625 11260 5633
rect 11226 5599 11260 5625
rect 11322 6543 11356 6569
rect 11322 6535 11356 6543
rect 11322 6475 11356 6497
rect 11322 6463 11356 6475
rect 11322 6407 11356 6425
rect 11322 6391 11356 6407
rect 11322 6339 11356 6353
rect 11322 6319 11356 6339
rect 11322 6271 11356 6281
rect 11322 6247 11356 6271
rect 11322 6203 11356 6209
rect 11322 6175 11356 6203
rect 11322 6135 11356 6137
rect 11322 6103 11356 6135
rect 11322 6033 11356 6065
rect 11322 6031 11356 6033
rect 11322 5965 11356 5993
rect 11322 5959 11356 5965
rect 11322 5897 11356 5921
rect 11322 5887 11356 5897
rect 11322 5829 11356 5849
rect 11322 5815 11356 5829
rect 11322 5761 11356 5777
rect 11322 5743 11356 5761
rect 11322 5693 11356 5705
rect 11322 5671 11356 5693
rect 11322 5625 11356 5633
rect 11322 5599 11356 5625
rect 11418 6543 11452 6569
rect 11418 6535 11452 6543
rect 11418 6475 11452 6497
rect 11418 6463 11452 6475
rect 11418 6407 11452 6425
rect 11418 6391 11452 6407
rect 11418 6339 11452 6353
rect 11418 6319 11452 6339
rect 11418 6271 11452 6281
rect 11418 6247 11452 6271
rect 11418 6203 11452 6209
rect 11418 6175 11452 6203
rect 11418 6135 11452 6137
rect 11418 6103 11452 6135
rect 11418 6033 11452 6065
rect 11418 6031 11452 6033
rect 11418 5965 11452 5993
rect 11418 5959 11452 5965
rect 11418 5897 11452 5921
rect 11418 5887 11452 5897
rect 11418 5829 11452 5849
rect 11418 5815 11452 5829
rect 11418 5761 11452 5777
rect 11418 5743 11452 5761
rect 11418 5693 11452 5705
rect 11418 5671 11452 5693
rect 11418 5625 11452 5633
rect 11418 5599 11452 5625
rect 11514 6543 11548 6569
rect 11514 6535 11548 6543
rect 11514 6475 11548 6497
rect 11514 6463 11548 6475
rect 11514 6407 11548 6425
rect 11514 6391 11548 6407
rect 11514 6339 11548 6353
rect 11514 6319 11548 6339
rect 11514 6271 11548 6281
rect 11514 6247 11548 6271
rect 11514 6203 11548 6209
rect 11514 6175 11548 6203
rect 11514 6135 11548 6137
rect 11514 6103 11548 6135
rect 11514 6033 11548 6065
rect 11514 6031 11548 6033
rect 11514 5965 11548 5993
rect 11514 5959 11548 5965
rect 11514 5897 11548 5921
rect 11514 5887 11548 5897
rect 11514 5829 11548 5849
rect 11514 5815 11548 5829
rect 11514 5761 11548 5777
rect 11514 5743 11548 5761
rect 11514 5693 11548 5705
rect 11514 5671 11548 5693
rect 11514 5625 11548 5633
rect 11514 5599 11548 5625
rect 11610 6543 11644 6569
rect 11610 6535 11644 6543
rect 11610 6475 11644 6497
rect 11610 6463 11644 6475
rect 11610 6407 11644 6425
rect 11610 6391 11644 6407
rect 11610 6339 11644 6353
rect 11610 6319 11644 6339
rect 11610 6271 11644 6281
rect 11610 6247 11644 6271
rect 11610 6203 11644 6209
rect 11610 6175 11644 6203
rect 11610 6135 11644 6137
rect 11610 6103 11644 6135
rect 11610 6033 11644 6065
rect 11610 6031 11644 6033
rect 11610 5965 11644 5993
rect 11610 5959 11644 5965
rect 11610 5897 11644 5921
rect 11610 5887 11644 5897
rect 11610 5829 11644 5849
rect 11610 5815 11644 5829
rect 11610 5761 11644 5777
rect 11610 5743 11644 5761
rect 11610 5693 11644 5705
rect 11610 5671 11644 5693
rect 11610 5625 11644 5633
rect 11610 5599 11644 5625
rect 11706 6543 11740 6569
rect 11706 6535 11740 6543
rect 11706 6475 11740 6497
rect 11706 6463 11740 6475
rect 11706 6407 11740 6425
rect 11706 6391 11740 6407
rect 11706 6339 11740 6353
rect 11706 6319 11740 6339
rect 11706 6271 11740 6281
rect 11706 6247 11740 6271
rect 11706 6203 11740 6209
rect 11706 6175 11740 6203
rect 11706 6135 11740 6137
rect 11706 6103 11740 6135
rect 11706 6033 11740 6065
rect 11706 6031 11740 6033
rect 11706 5965 11740 5993
rect 11706 5959 11740 5965
rect 11706 5897 11740 5921
rect 11706 5887 11740 5897
rect 11706 5829 11740 5849
rect 11706 5815 11740 5829
rect 11706 5761 11740 5777
rect 11706 5743 11740 5761
rect 11706 5693 11740 5705
rect 11706 5671 11740 5693
rect 11706 5625 11740 5633
rect 11706 5599 11740 5625
rect 11802 6543 11836 6569
rect 11802 6535 11836 6543
rect 11802 6475 11836 6497
rect 11802 6463 11836 6475
rect 11802 6407 11836 6425
rect 11802 6391 11836 6407
rect 11802 6339 11836 6353
rect 11802 6319 11836 6339
rect 11802 6271 11836 6281
rect 11802 6247 11836 6271
rect 11802 6203 11836 6209
rect 11802 6175 11836 6203
rect 11802 6135 11836 6137
rect 11802 6103 11836 6135
rect 11802 6033 11836 6065
rect 11802 6031 11836 6033
rect 11802 5965 11836 5993
rect 11802 5959 11836 5965
rect 11802 5897 11836 5921
rect 11802 5887 11836 5897
rect 11802 5829 11836 5849
rect 11802 5815 11836 5829
rect 11802 5761 11836 5777
rect 11802 5743 11836 5761
rect 11802 5693 11836 5705
rect 11802 5671 11836 5693
rect 11802 5625 11836 5633
rect 11802 5599 11836 5625
rect 12424 6521 12458 6547
rect 12424 6513 12458 6521
rect 12424 6453 12458 6475
rect 12424 6441 12458 6453
rect 12424 6385 12458 6403
rect 12424 6369 12458 6385
rect 12424 6317 12458 6331
rect 12424 6297 12458 6317
rect 12424 6249 12458 6259
rect 12424 6225 12458 6249
rect 12424 6181 12458 6187
rect 12424 6153 12458 6181
rect 12424 6113 12458 6115
rect 12424 6081 12458 6113
rect 12424 6011 12458 6043
rect 12424 6009 12458 6011
rect 12424 5943 12458 5971
rect 12424 5937 12458 5943
rect 12424 5875 12458 5899
rect 12424 5865 12458 5875
rect 12424 5807 12458 5827
rect 12424 5793 12458 5807
rect 12424 5739 12458 5755
rect 12424 5721 12458 5739
rect 12424 5671 12458 5683
rect 12424 5649 12458 5671
rect 12424 5603 12458 5611
rect 12424 5577 12458 5603
rect 12520 6521 12554 6547
rect 12520 6513 12554 6521
rect 12520 6453 12554 6475
rect 12520 6441 12554 6453
rect 12520 6385 12554 6403
rect 12520 6369 12554 6385
rect 12520 6317 12554 6331
rect 12520 6297 12554 6317
rect 12520 6249 12554 6259
rect 12520 6225 12554 6249
rect 12520 6181 12554 6187
rect 12520 6153 12554 6181
rect 12520 6113 12554 6115
rect 12520 6081 12554 6113
rect 12520 6011 12554 6043
rect 12520 6009 12554 6011
rect 12520 5943 12554 5971
rect 12520 5937 12554 5943
rect 12520 5875 12554 5899
rect 12520 5865 12554 5875
rect 12520 5807 12554 5827
rect 12520 5793 12554 5807
rect 12520 5739 12554 5755
rect 12520 5721 12554 5739
rect 12520 5671 12554 5683
rect 12520 5649 12554 5671
rect 12520 5603 12554 5611
rect 12520 5577 12554 5603
rect 6854 5352 6956 5398
rect 8268 5356 8370 5402
rect 12616 6521 12650 6547
rect 12616 6513 12650 6521
rect 12616 6453 12650 6475
rect 12616 6441 12650 6453
rect 12616 6385 12650 6403
rect 12616 6369 12650 6385
rect 12616 6317 12650 6331
rect 12616 6297 12650 6317
rect 12616 6249 12650 6259
rect 12616 6225 12650 6249
rect 12616 6181 12650 6187
rect 12616 6153 12650 6181
rect 12616 6113 12650 6115
rect 12616 6081 12650 6113
rect 12616 6011 12650 6043
rect 12616 6009 12650 6011
rect 12616 5943 12650 5971
rect 12616 5937 12650 5943
rect 12616 5875 12650 5899
rect 12616 5865 12650 5875
rect 12616 5807 12650 5827
rect 12616 5793 12650 5807
rect 12616 5739 12650 5755
rect 12616 5721 12650 5739
rect 12616 5671 12650 5683
rect 12616 5649 12650 5671
rect 12616 5603 12650 5611
rect 12616 5577 12650 5603
rect 12712 6521 12746 6547
rect 12712 6513 12746 6521
rect 12712 6453 12746 6475
rect 12712 6441 12746 6453
rect 12712 6385 12746 6403
rect 12712 6369 12746 6385
rect 12712 6317 12746 6331
rect 12712 6297 12746 6317
rect 12712 6249 12746 6259
rect 12712 6225 12746 6249
rect 12712 6181 12746 6187
rect 12712 6153 12746 6181
rect 12712 6113 12746 6115
rect 12712 6081 12746 6113
rect 12712 6011 12746 6043
rect 12712 6009 12746 6011
rect 12712 5943 12746 5971
rect 12712 5937 12746 5943
rect 12712 5875 12746 5899
rect 12712 5865 12746 5875
rect 12712 5807 12746 5827
rect 12712 5793 12746 5807
rect 12712 5739 12746 5755
rect 12712 5721 12746 5739
rect 12712 5671 12746 5683
rect 12712 5649 12746 5671
rect 12712 5603 12746 5611
rect 12712 5577 12746 5603
rect 12808 6521 12842 6547
rect 12808 6513 12842 6521
rect 12808 6453 12842 6475
rect 12808 6441 12842 6453
rect 12808 6385 12842 6403
rect 12808 6369 12842 6385
rect 12808 6317 12842 6331
rect 12808 6297 12842 6317
rect 12808 6249 12842 6259
rect 12808 6225 12842 6249
rect 12808 6181 12842 6187
rect 12808 6153 12842 6181
rect 12808 6113 12842 6115
rect 12808 6081 12842 6113
rect 12808 6011 12842 6043
rect 12808 6009 12842 6011
rect 12808 5943 12842 5971
rect 12808 5937 12842 5943
rect 12808 5875 12842 5899
rect 12808 5865 12842 5875
rect 12808 5807 12842 5827
rect 12808 5793 12842 5807
rect 12808 5739 12842 5755
rect 12808 5721 12842 5739
rect 12808 5671 12842 5683
rect 12808 5649 12842 5671
rect 12808 5603 12842 5611
rect 12808 5577 12842 5603
rect 12904 6521 12938 6547
rect 12904 6513 12938 6521
rect 12904 6453 12938 6475
rect 12904 6441 12938 6453
rect 12904 6385 12938 6403
rect 12904 6369 12938 6385
rect 12904 6317 12938 6331
rect 12904 6297 12938 6317
rect 12904 6249 12938 6259
rect 12904 6225 12938 6249
rect 12904 6181 12938 6187
rect 12904 6153 12938 6181
rect 12904 6113 12938 6115
rect 12904 6081 12938 6113
rect 12904 6011 12938 6043
rect 12904 6009 12938 6011
rect 12904 5943 12938 5971
rect 12904 5937 12938 5943
rect 12904 5875 12938 5899
rect 12904 5865 12938 5875
rect 12904 5807 12938 5827
rect 12904 5793 12938 5807
rect 12904 5739 12938 5755
rect 12904 5721 12938 5739
rect 12904 5671 12938 5683
rect 12904 5649 12938 5671
rect 12904 5603 12938 5611
rect 12904 5577 12938 5603
rect 13000 6521 13034 6547
rect 13000 6513 13034 6521
rect 13000 6453 13034 6475
rect 13000 6441 13034 6453
rect 13000 6385 13034 6403
rect 13000 6369 13034 6385
rect 13000 6317 13034 6331
rect 13000 6297 13034 6317
rect 13000 6249 13034 6259
rect 13000 6225 13034 6249
rect 13000 6181 13034 6187
rect 13000 6153 13034 6181
rect 13000 6113 13034 6115
rect 13000 6081 13034 6113
rect 13000 6011 13034 6043
rect 13000 6009 13034 6011
rect 13000 5943 13034 5971
rect 13000 5937 13034 5943
rect 13000 5875 13034 5899
rect 13000 5865 13034 5875
rect 13000 5807 13034 5827
rect 13000 5793 13034 5807
rect 13000 5739 13034 5755
rect 13000 5721 13034 5739
rect 13000 5671 13034 5683
rect 13000 5649 13034 5671
rect 13000 5603 13034 5611
rect 13000 5577 13034 5603
rect 13096 6521 13130 6547
rect 13096 6513 13130 6521
rect 13096 6453 13130 6475
rect 13096 6441 13130 6453
rect 13096 6385 13130 6403
rect 13096 6369 13130 6385
rect 13096 6317 13130 6331
rect 13096 6297 13130 6317
rect 13096 6249 13130 6259
rect 13096 6225 13130 6249
rect 13096 6181 13130 6187
rect 13096 6153 13130 6181
rect 13096 6113 13130 6115
rect 13096 6081 13130 6113
rect 13096 6011 13130 6043
rect 13096 6009 13130 6011
rect 13096 5943 13130 5971
rect 13096 5937 13130 5943
rect 13096 5875 13130 5899
rect 13096 5865 13130 5875
rect 13096 5807 13130 5827
rect 13096 5793 13130 5807
rect 13096 5739 13130 5755
rect 13096 5721 13130 5739
rect 13096 5671 13130 5683
rect 13096 5649 13130 5671
rect 13096 5603 13130 5611
rect 13096 5577 13130 5603
rect 13192 6521 13226 6547
rect 13192 6513 13226 6521
rect 13192 6453 13226 6475
rect 13192 6441 13226 6453
rect 13192 6385 13226 6403
rect 13192 6369 13226 6385
rect 13192 6317 13226 6331
rect 13192 6297 13226 6317
rect 13192 6249 13226 6259
rect 13192 6225 13226 6249
rect 13192 6181 13226 6187
rect 13192 6153 13226 6181
rect 13192 6113 13226 6115
rect 13192 6081 13226 6113
rect 13192 6011 13226 6043
rect 13192 6009 13226 6011
rect 13192 5943 13226 5971
rect 13192 5937 13226 5943
rect 13192 5875 13226 5899
rect 13192 5865 13226 5875
rect 13192 5807 13226 5827
rect 13192 5793 13226 5807
rect 13192 5739 13226 5755
rect 13192 5721 13226 5739
rect 13192 5671 13226 5683
rect 13192 5649 13226 5671
rect 13192 5603 13226 5611
rect 13192 5577 13226 5603
rect 13288 6521 13322 6547
rect 13288 6513 13322 6521
rect 13288 6453 13322 6475
rect 13288 6441 13322 6453
rect 13288 6385 13322 6403
rect 13288 6369 13322 6385
rect 13288 6317 13322 6331
rect 13288 6297 13322 6317
rect 13288 6249 13322 6259
rect 13288 6225 13322 6249
rect 13288 6181 13322 6187
rect 13288 6153 13322 6181
rect 13288 6113 13322 6115
rect 13288 6081 13322 6113
rect 13288 6011 13322 6043
rect 13288 6009 13322 6011
rect 13288 5943 13322 5971
rect 13288 5937 13322 5943
rect 13288 5875 13322 5899
rect 13288 5865 13322 5875
rect 13288 5807 13322 5827
rect 13288 5793 13322 5807
rect 13288 5739 13322 5755
rect 13288 5721 13322 5739
rect 13288 5671 13322 5683
rect 13288 5649 13322 5671
rect 13288 5603 13322 5611
rect 13288 5577 13322 5603
rect 13384 6521 13418 6547
rect 13384 6513 13418 6521
rect 13384 6453 13418 6475
rect 13384 6441 13418 6453
rect 13384 6385 13418 6403
rect 13384 6369 13418 6385
rect 13384 6317 13418 6331
rect 13384 6297 13418 6317
rect 13384 6249 13418 6259
rect 13384 6225 13418 6249
rect 13384 6181 13418 6187
rect 13384 6153 13418 6181
rect 13384 6113 13418 6115
rect 13384 6081 13418 6113
rect 13384 6011 13418 6043
rect 13384 6009 13418 6011
rect 13384 5943 13418 5971
rect 13384 5937 13418 5943
rect 13384 5875 13418 5899
rect 13384 5865 13418 5875
rect 13384 5807 13418 5827
rect 13384 5793 13418 5807
rect 13384 5739 13418 5755
rect 13384 5721 13418 5739
rect 13384 5671 13418 5683
rect 13384 5649 13418 5671
rect 13384 5603 13418 5611
rect 13384 5577 13418 5603
rect 13480 6521 13514 6547
rect 13480 6513 13514 6521
rect 13480 6453 13514 6475
rect 13480 6441 13514 6453
rect 13480 6385 13514 6403
rect 13480 6369 13514 6385
rect 13480 6317 13514 6331
rect 13480 6297 13514 6317
rect 13480 6249 13514 6259
rect 13480 6225 13514 6249
rect 13480 6181 13514 6187
rect 13480 6153 13514 6181
rect 13480 6113 13514 6115
rect 13480 6081 13514 6113
rect 13480 6011 13514 6043
rect 13480 6009 13514 6011
rect 13480 5943 13514 5971
rect 13480 5937 13514 5943
rect 13480 5875 13514 5899
rect 13480 5865 13514 5875
rect 13480 5807 13514 5827
rect 13480 5793 13514 5807
rect 13480 5739 13514 5755
rect 13480 5721 13514 5739
rect 13480 5671 13514 5683
rect 13480 5649 13514 5671
rect 13480 5603 13514 5611
rect 13480 5577 13514 5603
rect 13576 6521 13610 6547
rect 13576 6513 13610 6521
rect 13576 6453 13610 6475
rect 13576 6441 13610 6453
rect 13576 6385 13610 6403
rect 13576 6369 13610 6385
rect 13576 6317 13610 6331
rect 13576 6297 13610 6317
rect 13576 6249 13610 6259
rect 13576 6225 13610 6249
rect 13576 6181 13610 6187
rect 13576 6153 13610 6181
rect 13576 6113 13610 6115
rect 13576 6081 13610 6113
rect 13576 6011 13610 6043
rect 13576 6009 13610 6011
rect 13576 5943 13610 5971
rect 13576 5937 13610 5943
rect 13576 5875 13610 5899
rect 13576 5865 13610 5875
rect 13576 5807 13610 5827
rect 13576 5793 13610 5807
rect 13576 5739 13610 5755
rect 13576 5721 13610 5739
rect 13576 5671 13610 5683
rect 13576 5649 13610 5671
rect 13576 5603 13610 5611
rect 13576 5577 13610 5603
rect 14190 6517 14224 6543
rect 14190 6509 14224 6517
rect 14190 6449 14224 6471
rect 14190 6437 14224 6449
rect 14190 6381 14224 6399
rect 14190 6365 14224 6381
rect 14190 6313 14224 6327
rect 14190 6293 14224 6313
rect 14190 6245 14224 6255
rect 14190 6221 14224 6245
rect 14190 6177 14224 6183
rect 14190 6149 14224 6177
rect 14190 6109 14224 6111
rect 14190 6077 14224 6109
rect 14190 6007 14224 6039
rect 14190 6005 14224 6007
rect 14190 5939 14224 5967
rect 14190 5933 14224 5939
rect 14190 5871 14224 5895
rect 14190 5861 14224 5871
rect 14190 5803 14224 5823
rect 14190 5789 14224 5803
rect 14190 5735 14224 5751
rect 14190 5717 14224 5735
rect 14190 5667 14224 5679
rect 14190 5645 14224 5667
rect 14190 5599 14224 5607
rect 14190 5573 14224 5599
rect 14286 6517 14320 6543
rect 14286 6509 14320 6517
rect 14286 6449 14320 6471
rect 14286 6437 14320 6449
rect 14286 6381 14320 6399
rect 14286 6365 14320 6381
rect 14286 6313 14320 6327
rect 14286 6293 14320 6313
rect 14286 6245 14320 6255
rect 14286 6221 14320 6245
rect 14286 6177 14320 6183
rect 14286 6149 14320 6177
rect 14286 6109 14320 6111
rect 14286 6077 14320 6109
rect 14286 6007 14320 6039
rect 14286 6005 14320 6007
rect 14286 5939 14320 5967
rect 14286 5933 14320 5939
rect 14286 5871 14320 5895
rect 14286 5861 14320 5871
rect 14286 5803 14320 5823
rect 14286 5789 14320 5803
rect 14286 5735 14320 5751
rect 14286 5717 14320 5735
rect 14286 5667 14320 5679
rect 14286 5645 14320 5667
rect 14286 5599 14320 5607
rect 14286 5573 14320 5599
rect 9950 5346 10052 5392
rect 14382 6517 14416 6543
rect 14382 6509 14416 6517
rect 14382 6449 14416 6471
rect 14382 6437 14416 6449
rect 14382 6381 14416 6399
rect 14382 6365 14416 6381
rect 14382 6313 14416 6327
rect 14382 6293 14416 6313
rect 14382 6245 14416 6255
rect 14382 6221 14416 6245
rect 14382 6177 14416 6183
rect 14382 6149 14416 6177
rect 14382 6109 14416 6111
rect 14382 6077 14416 6109
rect 14382 6007 14416 6039
rect 14382 6005 14416 6007
rect 14382 5939 14416 5967
rect 14382 5933 14416 5939
rect 14382 5871 14416 5895
rect 14382 5861 14416 5871
rect 14382 5803 14416 5823
rect 14382 5789 14416 5803
rect 14382 5735 14416 5751
rect 14382 5717 14416 5735
rect 14382 5667 14416 5679
rect 14382 5645 14416 5667
rect 14382 5599 14416 5607
rect 14382 5573 14416 5599
rect 14478 6517 14512 6543
rect 14478 6509 14512 6517
rect 14478 6449 14512 6471
rect 14478 6437 14512 6449
rect 14478 6381 14512 6399
rect 14478 6365 14512 6381
rect 14478 6313 14512 6327
rect 14478 6293 14512 6313
rect 14478 6245 14512 6255
rect 14478 6221 14512 6245
rect 14478 6177 14512 6183
rect 14478 6149 14512 6177
rect 14478 6109 14512 6111
rect 14478 6077 14512 6109
rect 14478 6007 14512 6039
rect 14478 6005 14512 6007
rect 14478 5939 14512 5967
rect 14478 5933 14512 5939
rect 14478 5871 14512 5895
rect 14478 5861 14512 5871
rect 14478 5803 14512 5823
rect 14478 5789 14512 5803
rect 14478 5735 14512 5751
rect 14478 5717 14512 5735
rect 14478 5667 14512 5679
rect 14478 5645 14512 5667
rect 14478 5599 14512 5607
rect 14478 5573 14512 5599
rect 14574 6517 14608 6543
rect 14574 6509 14608 6517
rect 14574 6449 14608 6471
rect 14574 6437 14608 6449
rect 14574 6381 14608 6399
rect 14574 6365 14608 6381
rect 14574 6313 14608 6327
rect 14574 6293 14608 6313
rect 14574 6245 14608 6255
rect 14574 6221 14608 6245
rect 14574 6177 14608 6183
rect 14574 6149 14608 6177
rect 14574 6109 14608 6111
rect 14574 6077 14608 6109
rect 14574 6007 14608 6039
rect 14574 6005 14608 6007
rect 14574 5939 14608 5967
rect 14574 5933 14608 5939
rect 14574 5871 14608 5895
rect 14574 5861 14608 5871
rect 14574 5803 14608 5823
rect 14574 5789 14608 5803
rect 14574 5735 14608 5751
rect 14574 5717 14608 5735
rect 14574 5667 14608 5679
rect 14574 5645 14608 5667
rect 14574 5599 14608 5607
rect 14574 5573 14608 5599
rect 14670 6517 14704 6543
rect 14670 6509 14704 6517
rect 14670 6449 14704 6471
rect 14670 6437 14704 6449
rect 14670 6381 14704 6399
rect 14670 6365 14704 6381
rect 14670 6313 14704 6327
rect 14670 6293 14704 6313
rect 14670 6245 14704 6255
rect 14670 6221 14704 6245
rect 14670 6177 14704 6183
rect 14670 6149 14704 6177
rect 14670 6109 14704 6111
rect 14670 6077 14704 6109
rect 14670 6007 14704 6039
rect 14670 6005 14704 6007
rect 14670 5939 14704 5967
rect 14670 5933 14704 5939
rect 14670 5871 14704 5895
rect 14670 5861 14704 5871
rect 14670 5803 14704 5823
rect 14670 5789 14704 5803
rect 14670 5735 14704 5751
rect 14670 5717 14704 5735
rect 14670 5667 14704 5679
rect 14670 5645 14704 5667
rect 14670 5599 14704 5607
rect 14670 5573 14704 5599
rect 14766 6517 14800 6543
rect 14766 6509 14800 6517
rect 14766 6449 14800 6471
rect 14766 6437 14800 6449
rect 14766 6381 14800 6399
rect 14766 6365 14800 6381
rect 14766 6313 14800 6327
rect 14766 6293 14800 6313
rect 14766 6245 14800 6255
rect 14766 6221 14800 6245
rect 14766 6177 14800 6183
rect 14766 6149 14800 6177
rect 14766 6109 14800 6111
rect 14766 6077 14800 6109
rect 14766 6007 14800 6039
rect 14766 6005 14800 6007
rect 14766 5939 14800 5967
rect 14766 5933 14800 5939
rect 14766 5871 14800 5895
rect 14766 5861 14800 5871
rect 14766 5803 14800 5823
rect 14766 5789 14800 5803
rect 14766 5735 14800 5751
rect 14766 5717 14800 5735
rect 14766 5667 14800 5679
rect 14766 5645 14800 5667
rect 14766 5599 14800 5607
rect 14766 5573 14800 5599
rect 14862 6517 14896 6543
rect 14862 6509 14896 6517
rect 14862 6449 14896 6471
rect 14862 6437 14896 6449
rect 14862 6381 14896 6399
rect 14862 6365 14896 6381
rect 14862 6313 14896 6327
rect 14862 6293 14896 6313
rect 14862 6245 14896 6255
rect 14862 6221 14896 6245
rect 14862 6177 14896 6183
rect 14862 6149 14896 6177
rect 14862 6109 14896 6111
rect 14862 6077 14896 6109
rect 14862 6007 14896 6039
rect 14862 6005 14896 6007
rect 14862 5939 14896 5967
rect 14862 5933 14896 5939
rect 14862 5871 14896 5895
rect 14862 5861 14896 5871
rect 14862 5803 14896 5823
rect 14862 5789 14896 5803
rect 14862 5735 14896 5751
rect 14862 5717 14896 5735
rect 14862 5667 14896 5679
rect 14862 5645 14896 5667
rect 14862 5599 14896 5607
rect 14862 5573 14896 5599
rect 14958 6517 14992 6543
rect 14958 6509 14992 6517
rect 14958 6449 14992 6471
rect 14958 6437 14992 6449
rect 14958 6381 14992 6399
rect 14958 6365 14992 6381
rect 14958 6313 14992 6327
rect 14958 6293 14992 6313
rect 14958 6245 14992 6255
rect 14958 6221 14992 6245
rect 14958 6177 14992 6183
rect 14958 6149 14992 6177
rect 14958 6109 14992 6111
rect 14958 6077 14992 6109
rect 14958 6007 14992 6039
rect 15614 6148 15648 6182
rect 14958 6005 14992 6007
rect 14958 5939 14992 5967
rect 14958 5933 14992 5939
rect 14958 5871 14992 5895
rect 14958 5861 14992 5871
rect 14958 5803 14992 5823
rect 14958 5789 14992 5803
rect 14958 5735 14992 5751
rect 14958 5717 14992 5735
rect 14958 5667 14992 5679
rect 14958 5645 14992 5667
rect 14958 5599 14992 5607
rect 14958 5573 14992 5599
rect 15518 5861 15552 5879
rect 15518 5845 15552 5861
rect 15518 5793 15552 5807
rect 15518 5773 15552 5793
rect 15518 5725 15552 5735
rect 15518 5701 15552 5725
rect 15518 5657 15552 5663
rect 15518 5629 15552 5657
rect 15518 5589 15552 5591
rect 15518 5557 15552 5589
rect 11354 5352 11456 5398
rect 15518 5487 15552 5519
rect 15518 5485 15552 5487
rect -868 5311 -834 5317
rect 13094 5320 13196 5366
rect 14510 5326 14612 5372
rect 15518 5419 15552 5447
rect 15518 5413 15552 5419
rect 15518 5351 15552 5375
rect 15518 5341 15552 5351
rect -868 5249 -834 5273
rect -868 5239 -834 5249
rect -868 5181 -834 5201
rect -868 5167 -834 5181
rect -868 5113 -834 5129
rect 15518 5283 15552 5303
rect 15518 5269 15552 5283
rect 15518 5215 15552 5231
rect 15518 5197 15552 5215
rect 15518 5147 15552 5159
rect 15518 5125 15552 5147
rect -868 5095 -834 5113
rect -868 5045 -834 5057
rect -868 5023 -834 5045
rect 1580 5090 1614 5124
rect 4536 5074 4570 5108
rect 7566 5074 7600 5108
rect 10654 5072 10688 5106
rect -868 4977 -834 4985
rect -868 4951 -834 4977
rect 1484 4903 1518 4929
rect 1484 4895 1518 4903
rect -22950 4673 -22772 4779
rect -20936 4665 -20758 4771
rect -18939 4666 -18761 4772
rect -16317 4683 -16139 4789
rect -14320 4672 -14142 4778
rect -12320 4676 -12142 4782
rect -9969 4679 -9791 4785
rect -7976 4671 -7798 4777
rect -5972 4672 -5794 4778
rect 1484 4835 1518 4857
rect 1484 4823 1518 4835
rect -1067 4735 -1033 4769
rect 1484 4767 1518 4785
rect 1484 4751 1518 4767
rect 1484 4699 1518 4713
rect 1484 4679 1518 4699
rect 1484 4631 1518 4641
rect -23586 4401 -23552 4427
rect -23586 4393 -23552 4401
rect -23586 4333 -23552 4355
rect -23586 4321 -23552 4333
rect -23586 4265 -23552 4283
rect -23586 4249 -23552 4265
rect -23586 4197 -23552 4211
rect -23586 4177 -23552 4197
rect -23586 4129 -23552 4139
rect -23586 4105 -23552 4129
rect -23586 4061 -23552 4067
rect -23586 4033 -23552 4061
rect -23586 3993 -23552 3995
rect -23586 3961 -23552 3993
rect -23586 3891 -23552 3923
rect -23586 3889 -23552 3891
rect -23586 3823 -23552 3851
rect -23586 3817 -23552 3823
rect -23586 3755 -23552 3779
rect -23586 3745 -23552 3755
rect -23586 3687 -23552 3707
rect -23586 3673 -23552 3687
rect -23586 3619 -23552 3635
rect -23586 3601 -23552 3619
rect -23586 3551 -23552 3563
rect -23586 3529 -23552 3551
rect -23586 3483 -23552 3491
rect -23586 3457 -23552 3483
rect -23490 4401 -23456 4427
rect -23490 4393 -23456 4401
rect -23490 4333 -23456 4355
rect -23490 4321 -23456 4333
rect -23490 4265 -23456 4283
rect -23490 4249 -23456 4265
rect -23490 4197 -23456 4211
rect -23490 4177 -23456 4197
rect -23490 4129 -23456 4139
rect -23490 4105 -23456 4129
rect -23490 4061 -23456 4067
rect -23490 4033 -23456 4061
rect -23490 3993 -23456 3995
rect -23490 3961 -23456 3993
rect -23490 3891 -23456 3923
rect -23490 3889 -23456 3891
rect -23490 3823 -23456 3851
rect -23490 3817 -23456 3823
rect -23490 3755 -23456 3779
rect -23490 3745 -23456 3755
rect -23490 3687 -23456 3707
rect -23490 3673 -23456 3687
rect -23490 3619 -23456 3635
rect -23490 3601 -23456 3619
rect -23490 3551 -23456 3563
rect -23490 3529 -23456 3551
rect -23490 3483 -23456 3491
rect -23490 3457 -23456 3483
rect -23394 4401 -23360 4427
rect -23394 4393 -23360 4401
rect -23394 4333 -23360 4355
rect -23394 4321 -23360 4333
rect -23394 4265 -23360 4283
rect -23394 4249 -23360 4265
rect -23394 4197 -23360 4211
rect -23394 4177 -23360 4197
rect -23394 4129 -23360 4139
rect -23394 4105 -23360 4129
rect -23394 4061 -23360 4067
rect -23394 4033 -23360 4061
rect -23394 3993 -23360 3995
rect -23394 3961 -23360 3993
rect -23394 3891 -23360 3923
rect -23394 3889 -23360 3891
rect -23394 3823 -23360 3851
rect -23394 3817 -23360 3823
rect -23394 3755 -23360 3779
rect -23394 3745 -23360 3755
rect -23394 3687 -23360 3707
rect -23394 3673 -23360 3687
rect -23394 3619 -23360 3635
rect -23394 3601 -23360 3619
rect -23394 3551 -23360 3563
rect -23394 3529 -23360 3551
rect -23394 3483 -23360 3491
rect -23394 3457 -23360 3483
rect -23298 4401 -23264 4427
rect -23298 4393 -23264 4401
rect -23298 4333 -23264 4355
rect -23298 4321 -23264 4333
rect -23298 4265 -23264 4283
rect -23298 4249 -23264 4265
rect -23298 4197 -23264 4211
rect -23298 4177 -23264 4197
rect -23298 4129 -23264 4139
rect -23298 4105 -23264 4129
rect -23298 4061 -23264 4067
rect -23298 4033 -23264 4061
rect -23298 3993 -23264 3995
rect -23298 3961 -23264 3993
rect -23298 3891 -23264 3923
rect -23298 3889 -23264 3891
rect -23298 3823 -23264 3851
rect -23298 3817 -23264 3823
rect -23298 3755 -23264 3779
rect -23298 3745 -23264 3755
rect -23298 3687 -23264 3707
rect -23298 3673 -23264 3687
rect -23298 3619 -23264 3635
rect -23298 3601 -23264 3619
rect -23298 3551 -23264 3563
rect -23298 3529 -23264 3551
rect -23298 3483 -23264 3491
rect -23298 3457 -23264 3483
rect -23202 4401 -23168 4427
rect -23202 4393 -23168 4401
rect -23202 4333 -23168 4355
rect -23202 4321 -23168 4333
rect -23202 4265 -23168 4283
rect -23202 4249 -23168 4265
rect -23202 4197 -23168 4211
rect -23202 4177 -23168 4197
rect -23202 4129 -23168 4139
rect -23202 4105 -23168 4129
rect -23202 4061 -23168 4067
rect -23202 4033 -23168 4061
rect -23202 3993 -23168 3995
rect -23202 3961 -23168 3993
rect -23202 3891 -23168 3923
rect -23202 3889 -23168 3891
rect -23202 3823 -23168 3851
rect -23202 3817 -23168 3823
rect -23202 3755 -23168 3779
rect -23202 3745 -23168 3755
rect -23202 3687 -23168 3707
rect -23202 3673 -23168 3687
rect -23202 3619 -23168 3635
rect -23202 3601 -23168 3619
rect -23202 3551 -23168 3563
rect -23202 3529 -23168 3551
rect -23202 3483 -23168 3491
rect -23202 3457 -23168 3483
rect -23106 4401 -23072 4427
rect -23106 4393 -23072 4401
rect -23106 4333 -23072 4355
rect -23106 4321 -23072 4333
rect -23106 4265 -23072 4283
rect -23106 4249 -23072 4265
rect -23106 4197 -23072 4211
rect -23106 4177 -23072 4197
rect -23106 4129 -23072 4139
rect -23106 4105 -23072 4129
rect -23106 4061 -23072 4067
rect -23106 4033 -23072 4061
rect -23106 3993 -23072 3995
rect -23106 3961 -23072 3993
rect -23106 3891 -23072 3923
rect -23106 3889 -23072 3891
rect -23106 3823 -23072 3851
rect -23106 3817 -23072 3823
rect -23106 3755 -23072 3779
rect -23106 3745 -23072 3755
rect -23106 3687 -23072 3707
rect -23106 3673 -23072 3687
rect -23106 3619 -23072 3635
rect -23106 3601 -23072 3619
rect -23106 3551 -23072 3563
rect -23106 3529 -23072 3551
rect -23106 3483 -23072 3491
rect -23106 3457 -23072 3483
rect -23010 4401 -22976 4427
rect -23010 4393 -22976 4401
rect -23010 4333 -22976 4355
rect -23010 4321 -22976 4333
rect -23010 4265 -22976 4283
rect -23010 4249 -22976 4265
rect -23010 4197 -22976 4211
rect -23010 4177 -22976 4197
rect -23010 4129 -22976 4139
rect -23010 4105 -22976 4129
rect -23010 4061 -22976 4067
rect -23010 4033 -22976 4061
rect -23010 3993 -22976 3995
rect -23010 3961 -22976 3993
rect -23010 3891 -22976 3923
rect -23010 3889 -22976 3891
rect -23010 3823 -22976 3851
rect -23010 3817 -22976 3823
rect -23010 3755 -22976 3779
rect -23010 3745 -22976 3755
rect -23010 3687 -22976 3707
rect -23010 3673 -22976 3687
rect -23010 3619 -22976 3635
rect -23010 3601 -22976 3619
rect -23010 3551 -22976 3563
rect -23010 3529 -22976 3551
rect -23010 3483 -22976 3491
rect -23010 3457 -22976 3483
rect -22914 4401 -22880 4427
rect -22914 4393 -22880 4401
rect -22914 4333 -22880 4355
rect -22914 4321 -22880 4333
rect -22914 4265 -22880 4283
rect -22914 4249 -22880 4265
rect -22914 4197 -22880 4211
rect -22914 4177 -22880 4197
rect -22914 4129 -22880 4139
rect -22914 4105 -22880 4129
rect -22914 4061 -22880 4067
rect -22914 4033 -22880 4061
rect -22914 3993 -22880 3995
rect -22914 3961 -22880 3993
rect -22914 3891 -22880 3923
rect -22914 3889 -22880 3891
rect -22914 3823 -22880 3851
rect -22914 3817 -22880 3823
rect -22914 3755 -22880 3779
rect -22914 3745 -22880 3755
rect -22914 3687 -22880 3707
rect -22914 3673 -22880 3687
rect -22914 3619 -22880 3635
rect -22914 3601 -22880 3619
rect -22914 3551 -22880 3563
rect -22914 3529 -22880 3551
rect -22914 3483 -22880 3491
rect -22914 3457 -22880 3483
rect -22818 4401 -22784 4427
rect -22818 4393 -22784 4401
rect -22818 4333 -22784 4355
rect -22818 4321 -22784 4333
rect -22818 4265 -22784 4283
rect -22818 4249 -22784 4265
rect -22818 4197 -22784 4211
rect -22818 4177 -22784 4197
rect -22818 4129 -22784 4139
rect -22818 4105 -22784 4129
rect -22818 4061 -22784 4067
rect -22818 4033 -22784 4061
rect -22818 3993 -22784 3995
rect -22818 3961 -22784 3993
rect -22818 3891 -22784 3923
rect -22818 3889 -22784 3891
rect -22818 3823 -22784 3851
rect -22818 3817 -22784 3823
rect -22818 3755 -22784 3779
rect -22818 3745 -22784 3755
rect -22818 3687 -22784 3707
rect -22818 3673 -22784 3687
rect -22818 3619 -22784 3635
rect -22818 3601 -22784 3619
rect -22818 3551 -22784 3563
rect -22818 3529 -22784 3551
rect -22818 3483 -22784 3491
rect -22818 3457 -22784 3483
rect -22722 4401 -22688 4427
rect -22722 4393 -22688 4401
rect -22722 4333 -22688 4355
rect -22722 4321 -22688 4333
rect -22722 4265 -22688 4283
rect -22722 4249 -22688 4265
rect -22722 4197 -22688 4211
rect -22722 4177 -22688 4197
rect -22722 4129 -22688 4139
rect -22722 4105 -22688 4129
rect -22722 4061 -22688 4067
rect -22722 4033 -22688 4061
rect -22722 3993 -22688 3995
rect -22722 3961 -22688 3993
rect -22722 3891 -22688 3923
rect -22722 3889 -22688 3891
rect -22722 3823 -22688 3851
rect -22722 3817 -22688 3823
rect -22722 3755 -22688 3779
rect -22722 3745 -22688 3755
rect -22722 3687 -22688 3707
rect -22722 3673 -22688 3687
rect -22722 3619 -22688 3635
rect -22722 3601 -22688 3619
rect -22722 3551 -22688 3563
rect -22722 3529 -22688 3551
rect -22722 3483 -22688 3491
rect -22722 3457 -22688 3483
rect -22626 4401 -22592 4427
rect -22626 4393 -22592 4401
rect -22626 4333 -22592 4355
rect -22626 4321 -22592 4333
rect -22626 4265 -22592 4283
rect -22626 4249 -22592 4265
rect -22626 4197 -22592 4211
rect -22626 4177 -22592 4197
rect -22626 4129 -22592 4139
rect -22626 4105 -22592 4129
rect -22626 4061 -22592 4067
rect -22626 4033 -22592 4061
rect -22626 3993 -22592 3995
rect -22626 3961 -22592 3993
rect -22626 3891 -22592 3923
rect -22626 3889 -22592 3891
rect -22626 3823 -22592 3851
rect -22626 3817 -22592 3823
rect -22626 3755 -22592 3779
rect -22626 3745 -22592 3755
rect -22626 3687 -22592 3707
rect -22626 3673 -22592 3687
rect -22626 3619 -22592 3635
rect -22626 3601 -22592 3619
rect -22626 3551 -22592 3563
rect -22626 3529 -22592 3551
rect -22626 3483 -22592 3491
rect -22626 3457 -22592 3483
rect -22530 4401 -22496 4427
rect -22530 4393 -22496 4401
rect -22530 4333 -22496 4355
rect -22530 4321 -22496 4333
rect -22530 4265 -22496 4283
rect -22530 4249 -22496 4265
rect -22530 4197 -22496 4211
rect -22530 4177 -22496 4197
rect -22530 4129 -22496 4139
rect -22530 4105 -22496 4129
rect -22530 4061 -22496 4067
rect -22530 4033 -22496 4061
rect -22530 3993 -22496 3995
rect -22530 3961 -22496 3993
rect -22530 3891 -22496 3923
rect -22530 3889 -22496 3891
rect -22530 3823 -22496 3851
rect -22530 3817 -22496 3823
rect -22530 3755 -22496 3779
rect -22530 3745 -22496 3755
rect -22530 3687 -22496 3707
rect -22530 3673 -22496 3687
rect -22530 3619 -22496 3635
rect -22530 3601 -22496 3619
rect -22530 3551 -22496 3563
rect -22530 3529 -22496 3551
rect -22530 3483 -22496 3491
rect -22530 3457 -22496 3483
rect -22434 4401 -22400 4427
rect -22434 4393 -22400 4401
rect -22434 4333 -22400 4355
rect -22434 4321 -22400 4333
rect -22434 4265 -22400 4283
rect -22434 4249 -22400 4265
rect -22434 4197 -22400 4211
rect -22434 4177 -22400 4197
rect -22434 4129 -22400 4139
rect -22434 4105 -22400 4129
rect -22434 4061 -22400 4067
rect -22434 4033 -22400 4061
rect -22434 3993 -22400 3995
rect -22434 3961 -22400 3993
rect -22434 3891 -22400 3923
rect -22434 3889 -22400 3891
rect -22434 3823 -22400 3851
rect -22434 3817 -22400 3823
rect -22434 3755 -22400 3779
rect -22434 3745 -22400 3755
rect -22434 3687 -22400 3707
rect -22434 3673 -22400 3687
rect -22434 3619 -22400 3635
rect -22434 3601 -22400 3619
rect -22434 3551 -22400 3563
rect -22434 3529 -22400 3551
rect -22434 3483 -22400 3491
rect -22434 3457 -22400 3483
rect -22338 4401 -22304 4427
rect -22338 4393 -22304 4401
rect -22338 4333 -22304 4355
rect -22338 4321 -22304 4333
rect -22338 4265 -22304 4283
rect -22338 4249 -22304 4265
rect -22338 4197 -22304 4211
rect -22338 4177 -22304 4197
rect -22338 4129 -22304 4139
rect -22338 4105 -22304 4129
rect -22338 4061 -22304 4067
rect -22338 4033 -22304 4061
rect -22338 3993 -22304 3995
rect -22338 3961 -22304 3993
rect -22338 3891 -22304 3923
rect -22338 3889 -22304 3891
rect -22338 3823 -22304 3851
rect -22338 3817 -22304 3823
rect -22338 3755 -22304 3779
rect -22338 3745 -22304 3755
rect -22338 3687 -22304 3707
rect -22338 3673 -22304 3687
rect -22338 3619 -22304 3635
rect -22338 3601 -22304 3619
rect -22338 3551 -22304 3563
rect -22338 3529 -22304 3551
rect -22338 3483 -22304 3491
rect -22338 3457 -22304 3483
rect -22242 4401 -22208 4427
rect -22242 4393 -22208 4401
rect -22242 4333 -22208 4355
rect -22242 4321 -22208 4333
rect -22242 4265 -22208 4283
rect -22242 4249 -22208 4265
rect -22242 4197 -22208 4211
rect -22242 4177 -22208 4197
rect -22242 4129 -22208 4139
rect -22242 4105 -22208 4129
rect -22242 4061 -22208 4067
rect -22242 4033 -22208 4061
rect -22242 3993 -22208 3995
rect -22242 3961 -22208 3993
rect -22242 3891 -22208 3923
rect -22242 3889 -22208 3891
rect -22242 3823 -22208 3851
rect -22242 3817 -22208 3823
rect -22242 3755 -22208 3779
rect -22242 3745 -22208 3755
rect -22242 3687 -22208 3707
rect -22242 3673 -22208 3687
rect -22242 3619 -22208 3635
rect -22242 3601 -22208 3619
rect -22242 3551 -22208 3563
rect -22242 3529 -22208 3551
rect -22242 3483 -22208 3491
rect -22242 3457 -22208 3483
rect -22146 4401 -22112 4427
rect -22146 4393 -22112 4401
rect -22146 4333 -22112 4355
rect -22146 4321 -22112 4333
rect -22146 4265 -22112 4283
rect -22146 4249 -22112 4265
rect -22146 4197 -22112 4211
rect -22146 4177 -22112 4197
rect -22146 4129 -22112 4139
rect -22146 4105 -22112 4129
rect -22146 4061 -22112 4067
rect -22146 4033 -22112 4061
rect -22146 3993 -22112 3995
rect -22146 3961 -22112 3993
rect -22146 3891 -22112 3923
rect -22146 3889 -22112 3891
rect -22146 3823 -22112 3851
rect -22146 3817 -22112 3823
rect -22146 3755 -22112 3779
rect -22146 3745 -22112 3755
rect -22146 3687 -22112 3707
rect -22146 3673 -22112 3687
rect -22146 3619 -22112 3635
rect -22146 3601 -22112 3619
rect -22146 3551 -22112 3563
rect -22146 3529 -22112 3551
rect -22146 3483 -22112 3491
rect -22146 3457 -22112 3483
rect -22050 4401 -22016 4427
rect -22050 4393 -22016 4401
rect -22050 4333 -22016 4355
rect -22050 4321 -22016 4333
rect -22050 4265 -22016 4283
rect -22050 4249 -22016 4265
rect -22050 4197 -22016 4211
rect -22050 4177 -22016 4197
rect -22050 4129 -22016 4139
rect -22050 4105 -22016 4129
rect -22050 4061 -22016 4067
rect -22050 4033 -22016 4061
rect -22050 3993 -22016 3995
rect -22050 3961 -22016 3993
rect -22050 3891 -22016 3923
rect -22050 3889 -22016 3891
rect -22050 3823 -22016 3851
rect -22050 3817 -22016 3823
rect -22050 3755 -22016 3779
rect -22050 3745 -22016 3755
rect -22050 3687 -22016 3707
rect -22050 3673 -22016 3687
rect -22050 3619 -22016 3635
rect -22050 3601 -22016 3619
rect -22050 3551 -22016 3563
rect -22050 3529 -22016 3551
rect -22050 3483 -22016 3491
rect -22050 3457 -22016 3483
rect -21954 4401 -21920 4427
rect -21954 4393 -21920 4401
rect -21954 4333 -21920 4355
rect -21954 4321 -21920 4333
rect -21954 4265 -21920 4283
rect -21954 4249 -21920 4265
rect -21954 4197 -21920 4211
rect -21954 4177 -21920 4197
rect -21954 4129 -21920 4139
rect -21954 4105 -21920 4129
rect -21954 4061 -21920 4067
rect -21954 4033 -21920 4061
rect -21954 3993 -21920 3995
rect -21954 3961 -21920 3993
rect -21954 3891 -21920 3923
rect -21954 3889 -21920 3891
rect -21954 3823 -21920 3851
rect -21954 3817 -21920 3823
rect -21954 3755 -21920 3779
rect -21954 3745 -21920 3755
rect -21954 3687 -21920 3707
rect -21954 3673 -21920 3687
rect -21954 3619 -21920 3635
rect -21954 3601 -21920 3619
rect -21954 3551 -21920 3563
rect -21954 3529 -21920 3551
rect -21954 3483 -21920 3491
rect -21954 3457 -21920 3483
rect -21858 4401 -21824 4427
rect -21858 4393 -21824 4401
rect -21858 4333 -21824 4355
rect -21858 4321 -21824 4333
rect -21858 4265 -21824 4283
rect -21858 4249 -21824 4265
rect -21858 4197 -21824 4211
rect -21858 4177 -21824 4197
rect -21858 4129 -21824 4139
rect -21858 4105 -21824 4129
rect -21858 4061 -21824 4067
rect -21858 4033 -21824 4061
rect -21858 3993 -21824 3995
rect -21858 3961 -21824 3993
rect -21858 3891 -21824 3923
rect -21858 3889 -21824 3891
rect -21858 3823 -21824 3851
rect -21858 3817 -21824 3823
rect -21858 3755 -21824 3779
rect -21858 3745 -21824 3755
rect -21858 3687 -21824 3707
rect -21858 3673 -21824 3687
rect -21858 3619 -21824 3635
rect -21858 3601 -21824 3619
rect -21858 3551 -21824 3563
rect -21858 3529 -21824 3551
rect -21858 3483 -21824 3491
rect -21858 3457 -21824 3483
rect -21762 4401 -21728 4427
rect -21762 4393 -21728 4401
rect -21762 4333 -21728 4355
rect -21762 4321 -21728 4333
rect -21762 4265 -21728 4283
rect -21762 4249 -21728 4265
rect -21762 4197 -21728 4211
rect -21762 4177 -21728 4197
rect -21762 4129 -21728 4139
rect -21762 4105 -21728 4129
rect -21762 4061 -21728 4067
rect -21762 4033 -21728 4061
rect -21762 3993 -21728 3995
rect -21762 3961 -21728 3993
rect -21762 3891 -21728 3923
rect -21762 3889 -21728 3891
rect -21762 3823 -21728 3851
rect -21762 3817 -21728 3823
rect -21762 3755 -21728 3779
rect -21762 3745 -21728 3755
rect -21762 3687 -21728 3707
rect -21762 3673 -21728 3687
rect -21762 3619 -21728 3635
rect -21762 3601 -21728 3619
rect -21762 3551 -21728 3563
rect -21762 3529 -21728 3551
rect -21762 3483 -21728 3491
rect -21762 3457 -21728 3483
rect -21666 4401 -21632 4427
rect -21666 4393 -21632 4401
rect -21666 4333 -21632 4355
rect -21666 4321 -21632 4333
rect -21666 4265 -21632 4283
rect -21666 4249 -21632 4265
rect -21666 4197 -21632 4211
rect -21666 4177 -21632 4197
rect -21666 4129 -21632 4139
rect -21666 4105 -21632 4129
rect -21666 4061 -21632 4067
rect -21666 4033 -21632 4061
rect -21666 3993 -21632 3995
rect -21666 3961 -21632 3993
rect -21666 3891 -21632 3923
rect -21666 3889 -21632 3891
rect -21666 3823 -21632 3851
rect -21666 3817 -21632 3823
rect -21666 3755 -21632 3779
rect -21666 3745 -21632 3755
rect -21666 3687 -21632 3707
rect -21666 3673 -21632 3687
rect -21666 3619 -21632 3635
rect -21666 3601 -21632 3619
rect -21666 3551 -21632 3563
rect -21666 3529 -21632 3551
rect -21666 3483 -21632 3491
rect -21666 3457 -21632 3483
rect -21442 4407 -21408 4433
rect -21442 4399 -21408 4407
rect -21442 4339 -21408 4361
rect -21442 4327 -21408 4339
rect -21442 4271 -21408 4289
rect -21442 4255 -21408 4271
rect -21442 4203 -21408 4217
rect -21442 4183 -21408 4203
rect -21442 4135 -21408 4145
rect -21442 4111 -21408 4135
rect -21442 4067 -21408 4073
rect -21442 4039 -21408 4067
rect -21442 3999 -21408 4001
rect -21442 3967 -21408 3999
rect -21442 3897 -21408 3929
rect -21442 3895 -21408 3897
rect -21442 3829 -21408 3857
rect -21442 3823 -21408 3829
rect -21442 3761 -21408 3785
rect -21442 3751 -21408 3761
rect -21442 3693 -21408 3713
rect -21442 3679 -21408 3693
rect -21442 3625 -21408 3641
rect -21442 3607 -21408 3625
rect -21442 3557 -21408 3569
rect -21442 3535 -21408 3557
rect -21442 3489 -21408 3497
rect -21442 3463 -21408 3489
rect -21346 4407 -21312 4433
rect -21346 4399 -21312 4407
rect -21346 4339 -21312 4361
rect -21346 4327 -21312 4339
rect -21346 4271 -21312 4289
rect -21346 4255 -21312 4271
rect -21346 4203 -21312 4217
rect -21346 4183 -21312 4203
rect -21346 4135 -21312 4145
rect -21346 4111 -21312 4135
rect -21346 4067 -21312 4073
rect -21346 4039 -21312 4067
rect -21346 3999 -21312 4001
rect -21346 3967 -21312 3999
rect -21346 3897 -21312 3929
rect -21346 3895 -21312 3897
rect -21346 3829 -21312 3857
rect -21346 3823 -21312 3829
rect -21346 3761 -21312 3785
rect -21346 3751 -21312 3761
rect -21346 3693 -21312 3713
rect -21346 3679 -21312 3693
rect -21346 3625 -21312 3641
rect -21346 3607 -21312 3625
rect -21346 3557 -21312 3569
rect -21346 3535 -21312 3557
rect -21346 3489 -21312 3497
rect -21346 3463 -21312 3489
rect -21250 4407 -21216 4433
rect -21250 4399 -21216 4407
rect -21250 4339 -21216 4361
rect -21250 4327 -21216 4339
rect -21250 4271 -21216 4289
rect -21250 4255 -21216 4271
rect -21250 4203 -21216 4217
rect -21250 4183 -21216 4203
rect -21250 4135 -21216 4145
rect -21250 4111 -21216 4135
rect -21250 4067 -21216 4073
rect -21250 4039 -21216 4067
rect -21250 3999 -21216 4001
rect -21250 3967 -21216 3999
rect -21250 3897 -21216 3929
rect -21250 3895 -21216 3897
rect -21250 3829 -21216 3857
rect -21250 3823 -21216 3829
rect -21250 3761 -21216 3785
rect -21250 3751 -21216 3761
rect -21250 3693 -21216 3713
rect -21250 3679 -21216 3693
rect -21250 3625 -21216 3641
rect -21250 3607 -21216 3625
rect -21250 3557 -21216 3569
rect -21250 3535 -21216 3557
rect -21250 3489 -21216 3497
rect -21250 3463 -21216 3489
rect -21154 4407 -21120 4433
rect -21154 4399 -21120 4407
rect -21154 4339 -21120 4361
rect -21154 4327 -21120 4339
rect -21154 4271 -21120 4289
rect -21154 4255 -21120 4271
rect -21154 4203 -21120 4217
rect -21154 4183 -21120 4203
rect -21154 4135 -21120 4145
rect -21154 4111 -21120 4135
rect -21154 4067 -21120 4073
rect -21154 4039 -21120 4067
rect -21154 3999 -21120 4001
rect -21154 3967 -21120 3999
rect -21154 3897 -21120 3929
rect -21154 3895 -21120 3897
rect -21154 3829 -21120 3857
rect -21154 3823 -21120 3829
rect -21154 3761 -21120 3785
rect -21154 3751 -21120 3761
rect -21154 3693 -21120 3713
rect -21154 3679 -21120 3693
rect -21154 3625 -21120 3641
rect -21154 3607 -21120 3625
rect -21154 3557 -21120 3569
rect -21154 3535 -21120 3557
rect -21154 3489 -21120 3497
rect -21154 3463 -21120 3489
rect -21058 4407 -21024 4433
rect -21058 4399 -21024 4407
rect -21058 4339 -21024 4361
rect -21058 4327 -21024 4339
rect -21058 4271 -21024 4289
rect -21058 4255 -21024 4271
rect -21058 4203 -21024 4217
rect -21058 4183 -21024 4203
rect -21058 4135 -21024 4145
rect -21058 4111 -21024 4135
rect -21058 4067 -21024 4073
rect -21058 4039 -21024 4067
rect -21058 3999 -21024 4001
rect -21058 3967 -21024 3999
rect -21058 3897 -21024 3929
rect -21058 3895 -21024 3897
rect -21058 3829 -21024 3857
rect -21058 3823 -21024 3829
rect -21058 3761 -21024 3785
rect -21058 3751 -21024 3761
rect -21058 3693 -21024 3713
rect -21058 3679 -21024 3693
rect -21058 3625 -21024 3641
rect -21058 3607 -21024 3625
rect -21058 3557 -21024 3569
rect -21058 3535 -21024 3557
rect -21058 3489 -21024 3497
rect -21058 3463 -21024 3489
rect -20962 4407 -20928 4433
rect -20962 4399 -20928 4407
rect -20962 4339 -20928 4361
rect -20962 4327 -20928 4339
rect -20962 4271 -20928 4289
rect -20962 4255 -20928 4271
rect -20962 4203 -20928 4217
rect -20962 4183 -20928 4203
rect -20962 4135 -20928 4145
rect -20962 4111 -20928 4135
rect -20962 4067 -20928 4073
rect -20962 4039 -20928 4067
rect -20962 3999 -20928 4001
rect -20962 3967 -20928 3999
rect -20962 3897 -20928 3929
rect -20962 3895 -20928 3897
rect -20962 3829 -20928 3857
rect -20962 3823 -20928 3829
rect -20962 3761 -20928 3785
rect -20962 3751 -20928 3761
rect -20962 3693 -20928 3713
rect -20962 3679 -20928 3693
rect -20962 3625 -20928 3641
rect -20962 3607 -20928 3625
rect -20962 3557 -20928 3569
rect -20962 3535 -20928 3557
rect -20962 3489 -20928 3497
rect -20962 3463 -20928 3489
rect -20866 4407 -20832 4433
rect -20866 4399 -20832 4407
rect -20866 4339 -20832 4361
rect -20866 4327 -20832 4339
rect -20866 4271 -20832 4289
rect -20866 4255 -20832 4271
rect -20866 4203 -20832 4217
rect -20866 4183 -20832 4203
rect -20866 4135 -20832 4145
rect -20866 4111 -20832 4135
rect -20866 4067 -20832 4073
rect -20866 4039 -20832 4067
rect -20866 3999 -20832 4001
rect -20866 3967 -20832 3999
rect -20866 3897 -20832 3929
rect -20866 3895 -20832 3897
rect -20866 3829 -20832 3857
rect -20866 3823 -20832 3829
rect -20866 3761 -20832 3785
rect -20866 3751 -20832 3761
rect -20866 3693 -20832 3713
rect -20866 3679 -20832 3693
rect -20866 3625 -20832 3641
rect -20866 3607 -20832 3625
rect -20866 3557 -20832 3569
rect -20866 3535 -20832 3557
rect -20866 3489 -20832 3497
rect -20866 3463 -20832 3489
rect -20770 4407 -20736 4433
rect -20770 4399 -20736 4407
rect -20770 4339 -20736 4361
rect -20770 4327 -20736 4339
rect -20770 4271 -20736 4289
rect -20770 4255 -20736 4271
rect -20770 4203 -20736 4217
rect -20770 4183 -20736 4203
rect -20770 4135 -20736 4145
rect -20770 4111 -20736 4135
rect -20770 4067 -20736 4073
rect -20770 4039 -20736 4067
rect -20770 3999 -20736 4001
rect -20770 3967 -20736 3999
rect -20770 3897 -20736 3929
rect -20770 3895 -20736 3897
rect -20770 3829 -20736 3857
rect -20770 3823 -20736 3829
rect -20770 3761 -20736 3785
rect -20770 3751 -20736 3761
rect -20770 3693 -20736 3713
rect -20770 3679 -20736 3693
rect -20770 3625 -20736 3641
rect -20770 3607 -20736 3625
rect -20770 3557 -20736 3569
rect -20770 3535 -20736 3557
rect -20770 3489 -20736 3497
rect -20770 3463 -20736 3489
rect -20674 4407 -20640 4433
rect -20674 4399 -20640 4407
rect -20674 4339 -20640 4361
rect -20674 4327 -20640 4339
rect -20674 4271 -20640 4289
rect -20674 4255 -20640 4271
rect -20674 4203 -20640 4217
rect -20674 4183 -20640 4203
rect -20674 4135 -20640 4145
rect -20674 4111 -20640 4135
rect -20674 4067 -20640 4073
rect -20674 4039 -20640 4067
rect -20674 3999 -20640 4001
rect -20674 3967 -20640 3999
rect -20674 3897 -20640 3929
rect -20674 3895 -20640 3897
rect -20674 3829 -20640 3857
rect -20674 3823 -20640 3829
rect -20674 3761 -20640 3785
rect -20674 3751 -20640 3761
rect -20674 3693 -20640 3713
rect -20674 3679 -20640 3693
rect -20674 3625 -20640 3641
rect -20674 3607 -20640 3625
rect -20674 3557 -20640 3569
rect -20674 3535 -20640 3557
rect -20674 3489 -20640 3497
rect -20674 3463 -20640 3489
rect -20578 4407 -20544 4433
rect -20578 4399 -20544 4407
rect -20578 4339 -20544 4361
rect -20578 4327 -20544 4339
rect -20578 4271 -20544 4289
rect -20578 4255 -20544 4271
rect -20578 4203 -20544 4217
rect -20578 4183 -20544 4203
rect -20578 4135 -20544 4145
rect -20578 4111 -20544 4135
rect -20578 4067 -20544 4073
rect -20578 4039 -20544 4067
rect -20578 3999 -20544 4001
rect -20578 3967 -20544 3999
rect -20578 3897 -20544 3929
rect -20578 3895 -20544 3897
rect -20578 3829 -20544 3857
rect -20578 3823 -20544 3829
rect -20578 3761 -20544 3785
rect -20578 3751 -20544 3761
rect -20578 3693 -20544 3713
rect -20578 3679 -20544 3693
rect -20578 3625 -20544 3641
rect -20578 3607 -20544 3625
rect -20578 3557 -20544 3569
rect -20578 3535 -20544 3557
rect -20578 3489 -20544 3497
rect -20578 3463 -20544 3489
rect -20482 4407 -20448 4433
rect -20482 4399 -20448 4407
rect -20482 4339 -20448 4361
rect -20482 4327 -20448 4339
rect -20482 4271 -20448 4289
rect -20482 4255 -20448 4271
rect -20482 4203 -20448 4217
rect -20482 4183 -20448 4203
rect -20482 4135 -20448 4145
rect -20482 4111 -20448 4135
rect -20482 4067 -20448 4073
rect -20482 4039 -20448 4067
rect -20482 3999 -20448 4001
rect -20482 3967 -20448 3999
rect -20482 3897 -20448 3929
rect -20482 3895 -20448 3897
rect -20482 3829 -20448 3857
rect -20482 3823 -20448 3829
rect -20482 3761 -20448 3785
rect -20482 3751 -20448 3761
rect -20482 3693 -20448 3713
rect -20482 3679 -20448 3693
rect -20482 3625 -20448 3641
rect -20482 3607 -20448 3625
rect -20482 3557 -20448 3569
rect -20482 3535 -20448 3557
rect -20482 3489 -20448 3497
rect -20482 3463 -20448 3489
rect -20386 4407 -20352 4433
rect -20386 4399 -20352 4407
rect -20386 4339 -20352 4361
rect -20386 4327 -20352 4339
rect -20386 4271 -20352 4289
rect -20386 4255 -20352 4271
rect -20386 4203 -20352 4217
rect -20386 4183 -20352 4203
rect -20386 4135 -20352 4145
rect -20386 4111 -20352 4135
rect -20386 4067 -20352 4073
rect -20386 4039 -20352 4067
rect -20386 3999 -20352 4001
rect -20386 3967 -20352 3999
rect -20386 3897 -20352 3929
rect -20386 3895 -20352 3897
rect -20386 3829 -20352 3857
rect -20386 3823 -20352 3829
rect -20386 3761 -20352 3785
rect -20386 3751 -20352 3761
rect -20386 3693 -20352 3713
rect -20386 3679 -20352 3693
rect -20386 3625 -20352 3641
rect -20386 3607 -20352 3625
rect -20386 3557 -20352 3569
rect -20386 3535 -20352 3557
rect -20386 3489 -20352 3497
rect -20386 3463 -20352 3489
rect -20290 4407 -20256 4433
rect -20290 4399 -20256 4407
rect -20290 4339 -20256 4361
rect -20290 4327 -20256 4339
rect -20290 4271 -20256 4289
rect -20290 4255 -20256 4271
rect -20290 4203 -20256 4217
rect -20290 4183 -20256 4203
rect -20290 4135 -20256 4145
rect -20290 4111 -20256 4135
rect -20290 4067 -20256 4073
rect -20290 4039 -20256 4067
rect -20290 3999 -20256 4001
rect -20290 3967 -20256 3999
rect -20290 3897 -20256 3929
rect -20290 3895 -20256 3897
rect -20290 3829 -20256 3857
rect -20290 3823 -20256 3829
rect -20290 3761 -20256 3785
rect -20290 3751 -20256 3761
rect -20290 3693 -20256 3713
rect -20290 3679 -20256 3693
rect -20290 3625 -20256 3641
rect -20290 3607 -20256 3625
rect -20290 3557 -20256 3569
rect -20290 3535 -20256 3557
rect -20290 3489 -20256 3497
rect -20290 3463 -20256 3489
rect -20194 4407 -20160 4433
rect -20194 4399 -20160 4407
rect -20194 4339 -20160 4361
rect -20194 4327 -20160 4339
rect -20194 4271 -20160 4289
rect -20194 4255 -20160 4271
rect -20194 4203 -20160 4217
rect -20194 4183 -20160 4203
rect -20194 4135 -20160 4145
rect -20194 4111 -20160 4135
rect -20194 4067 -20160 4073
rect -20194 4039 -20160 4067
rect -20194 3999 -20160 4001
rect -20194 3967 -20160 3999
rect -20194 3897 -20160 3929
rect -20194 3895 -20160 3897
rect -20194 3829 -20160 3857
rect -20194 3823 -20160 3829
rect -20194 3761 -20160 3785
rect -20194 3751 -20160 3761
rect -20194 3693 -20160 3713
rect -20194 3679 -20160 3693
rect -20194 3625 -20160 3641
rect -20194 3607 -20160 3625
rect -20194 3557 -20160 3569
rect -20194 3535 -20160 3557
rect -20194 3489 -20160 3497
rect -20194 3463 -20160 3489
rect -20098 4407 -20064 4433
rect -20098 4399 -20064 4407
rect -20098 4339 -20064 4361
rect -20098 4327 -20064 4339
rect -20098 4271 -20064 4289
rect -20098 4255 -20064 4271
rect -20098 4203 -20064 4217
rect -20098 4183 -20064 4203
rect -20098 4135 -20064 4145
rect -20098 4111 -20064 4135
rect -20098 4067 -20064 4073
rect -20098 4039 -20064 4067
rect -20098 3999 -20064 4001
rect -20098 3967 -20064 3999
rect -20098 3897 -20064 3929
rect -20098 3895 -20064 3897
rect -20098 3829 -20064 3857
rect -20098 3823 -20064 3829
rect -20098 3761 -20064 3785
rect -20098 3751 -20064 3761
rect -20098 3693 -20064 3713
rect -20098 3679 -20064 3693
rect -20098 3625 -20064 3641
rect -20098 3607 -20064 3625
rect -20098 3557 -20064 3569
rect -20098 3535 -20064 3557
rect -20098 3489 -20064 3497
rect -20098 3463 -20064 3489
rect -20002 4407 -19968 4433
rect -20002 4399 -19968 4407
rect -20002 4339 -19968 4361
rect -20002 4327 -19968 4339
rect -20002 4271 -19968 4289
rect -20002 4255 -19968 4271
rect -20002 4203 -19968 4217
rect -20002 4183 -19968 4203
rect -20002 4135 -19968 4145
rect -20002 4111 -19968 4135
rect -20002 4067 -19968 4073
rect -20002 4039 -19968 4067
rect -20002 3999 -19968 4001
rect -20002 3967 -19968 3999
rect -20002 3897 -19968 3929
rect -20002 3895 -19968 3897
rect -20002 3829 -19968 3857
rect -20002 3823 -19968 3829
rect -20002 3761 -19968 3785
rect -20002 3751 -19968 3761
rect -20002 3693 -19968 3713
rect -20002 3679 -19968 3693
rect -20002 3625 -19968 3641
rect -20002 3607 -19968 3625
rect -20002 3557 -19968 3569
rect -20002 3535 -19968 3557
rect -20002 3489 -19968 3497
rect -20002 3463 -19968 3489
rect -19758 4413 -19724 4439
rect -19758 4405 -19724 4413
rect -19758 4345 -19724 4367
rect -19758 4333 -19724 4345
rect -19758 4277 -19724 4295
rect -19758 4261 -19724 4277
rect -19758 4209 -19724 4223
rect -19758 4189 -19724 4209
rect -19758 4141 -19724 4151
rect -19758 4117 -19724 4141
rect -19758 4073 -19724 4079
rect -19758 4045 -19724 4073
rect -19758 4005 -19724 4007
rect -19758 3973 -19724 4005
rect -19758 3903 -19724 3935
rect -19758 3901 -19724 3903
rect -19758 3835 -19724 3863
rect -19758 3829 -19724 3835
rect -19758 3767 -19724 3791
rect -19758 3757 -19724 3767
rect -19758 3699 -19724 3719
rect -19758 3685 -19724 3699
rect -19758 3631 -19724 3647
rect -19758 3613 -19724 3631
rect -19758 3563 -19724 3575
rect -19758 3541 -19724 3563
rect -19758 3495 -19724 3503
rect -19758 3469 -19724 3495
rect -19662 4413 -19628 4439
rect -19662 4405 -19628 4413
rect -19662 4345 -19628 4367
rect -19662 4333 -19628 4345
rect -19662 4277 -19628 4295
rect -19662 4261 -19628 4277
rect -19662 4209 -19628 4223
rect -19662 4189 -19628 4209
rect -19662 4141 -19628 4151
rect -19662 4117 -19628 4141
rect -19662 4073 -19628 4079
rect -19662 4045 -19628 4073
rect -19662 4005 -19628 4007
rect -19662 3973 -19628 4005
rect -19662 3903 -19628 3935
rect -19662 3901 -19628 3903
rect -19662 3835 -19628 3863
rect -19662 3829 -19628 3835
rect -19662 3767 -19628 3791
rect -19662 3757 -19628 3767
rect -19662 3699 -19628 3719
rect -19662 3685 -19628 3699
rect -19662 3631 -19628 3647
rect -19662 3613 -19628 3631
rect -19662 3563 -19628 3575
rect -19662 3541 -19628 3563
rect -19662 3495 -19628 3503
rect -19662 3469 -19628 3495
rect -19566 4413 -19532 4439
rect -19566 4405 -19532 4413
rect -19566 4345 -19532 4367
rect -19566 4333 -19532 4345
rect -19566 4277 -19532 4295
rect -19566 4261 -19532 4277
rect -19566 4209 -19532 4223
rect -19566 4189 -19532 4209
rect -19566 4141 -19532 4151
rect -19566 4117 -19532 4141
rect -19566 4073 -19532 4079
rect -19566 4045 -19532 4073
rect -19566 4005 -19532 4007
rect -19566 3973 -19532 4005
rect -19566 3903 -19532 3935
rect -19566 3901 -19532 3903
rect -19566 3835 -19532 3863
rect -19566 3829 -19532 3835
rect -19566 3767 -19532 3791
rect -19566 3757 -19532 3767
rect -19566 3699 -19532 3719
rect -19566 3685 -19532 3699
rect -19566 3631 -19532 3647
rect -19566 3613 -19532 3631
rect -19566 3563 -19532 3575
rect -19566 3541 -19532 3563
rect -19566 3495 -19532 3503
rect -19566 3469 -19532 3495
rect -19470 4413 -19436 4439
rect -19470 4405 -19436 4413
rect -19470 4345 -19436 4367
rect -19470 4333 -19436 4345
rect -19470 4277 -19436 4295
rect -19470 4261 -19436 4277
rect -19470 4209 -19436 4223
rect -19470 4189 -19436 4209
rect -19470 4141 -19436 4151
rect -19470 4117 -19436 4141
rect -19470 4073 -19436 4079
rect -19470 4045 -19436 4073
rect -19470 4005 -19436 4007
rect -19470 3973 -19436 4005
rect -19470 3903 -19436 3935
rect -19470 3901 -19436 3903
rect -19470 3835 -19436 3863
rect -19470 3829 -19436 3835
rect -19470 3767 -19436 3791
rect -19470 3757 -19436 3767
rect -19470 3699 -19436 3719
rect -19470 3685 -19436 3699
rect -19470 3631 -19436 3647
rect -19470 3613 -19436 3631
rect -19470 3563 -19436 3575
rect -19470 3541 -19436 3563
rect -19470 3495 -19436 3503
rect -19470 3469 -19436 3495
rect -19374 4413 -19340 4439
rect -19374 4405 -19340 4413
rect -19374 4345 -19340 4367
rect -19374 4333 -19340 4345
rect -19374 4277 -19340 4295
rect -19374 4261 -19340 4277
rect -19374 4209 -19340 4223
rect -19374 4189 -19340 4209
rect -19374 4141 -19340 4151
rect -19374 4117 -19340 4141
rect -19374 4073 -19340 4079
rect -19374 4045 -19340 4073
rect -19374 4005 -19340 4007
rect -19374 3973 -19340 4005
rect -19374 3903 -19340 3935
rect -19374 3901 -19340 3903
rect -19374 3835 -19340 3863
rect -19374 3829 -19340 3835
rect -19374 3767 -19340 3791
rect -19374 3757 -19340 3767
rect -19374 3699 -19340 3719
rect -19374 3685 -19340 3699
rect -19374 3631 -19340 3647
rect -19374 3613 -19340 3631
rect -19374 3563 -19340 3575
rect -19374 3541 -19340 3563
rect -19374 3495 -19340 3503
rect -19374 3469 -19340 3495
rect -19278 4413 -19244 4439
rect -19278 4405 -19244 4413
rect -19278 4345 -19244 4367
rect -19278 4333 -19244 4345
rect -19278 4277 -19244 4295
rect -19278 4261 -19244 4277
rect -19278 4209 -19244 4223
rect -19278 4189 -19244 4209
rect -19278 4141 -19244 4151
rect -19278 4117 -19244 4141
rect -19278 4073 -19244 4079
rect -19278 4045 -19244 4073
rect -19278 4005 -19244 4007
rect -19278 3973 -19244 4005
rect -19278 3903 -19244 3935
rect -19278 3901 -19244 3903
rect -19278 3835 -19244 3863
rect -19278 3829 -19244 3835
rect -19278 3767 -19244 3791
rect -19278 3757 -19244 3767
rect -19278 3699 -19244 3719
rect -19278 3685 -19244 3699
rect -19278 3631 -19244 3647
rect -19278 3613 -19244 3631
rect -19278 3563 -19244 3575
rect -19278 3541 -19244 3563
rect -19278 3495 -19244 3503
rect -19278 3469 -19244 3495
rect -19182 4413 -19148 4439
rect -19182 4405 -19148 4413
rect -19182 4345 -19148 4367
rect -19182 4333 -19148 4345
rect -19182 4277 -19148 4295
rect -19182 4261 -19148 4277
rect -19182 4209 -19148 4223
rect -19182 4189 -19148 4209
rect -19182 4141 -19148 4151
rect -19182 4117 -19148 4141
rect -19182 4073 -19148 4079
rect -19182 4045 -19148 4073
rect -19182 4005 -19148 4007
rect -19182 3973 -19148 4005
rect -19182 3903 -19148 3935
rect -19182 3901 -19148 3903
rect -19182 3835 -19148 3863
rect -19182 3829 -19148 3835
rect -19182 3767 -19148 3791
rect -19182 3757 -19148 3767
rect -19182 3699 -19148 3719
rect -19182 3685 -19148 3699
rect -19182 3631 -19148 3647
rect -19182 3613 -19148 3631
rect -19182 3563 -19148 3575
rect -19182 3541 -19148 3563
rect -19182 3495 -19148 3503
rect -19182 3469 -19148 3495
rect -19086 4413 -19052 4439
rect -19086 4405 -19052 4413
rect -19086 4345 -19052 4367
rect -19086 4333 -19052 4345
rect -19086 4277 -19052 4295
rect -19086 4261 -19052 4277
rect -19086 4209 -19052 4223
rect -19086 4189 -19052 4209
rect -19086 4141 -19052 4151
rect -19086 4117 -19052 4141
rect -19086 4073 -19052 4079
rect -19086 4045 -19052 4073
rect -19086 4005 -19052 4007
rect -19086 3973 -19052 4005
rect -19086 3903 -19052 3935
rect -19086 3901 -19052 3903
rect -19086 3835 -19052 3863
rect -19086 3829 -19052 3835
rect -19086 3767 -19052 3791
rect -19086 3757 -19052 3767
rect -19086 3699 -19052 3719
rect -19086 3685 -19052 3699
rect -19086 3631 -19052 3647
rect -19086 3613 -19052 3631
rect -19086 3563 -19052 3575
rect -19086 3541 -19052 3563
rect -19086 3495 -19052 3503
rect -19086 3469 -19052 3495
rect -18990 4413 -18956 4439
rect -18990 4405 -18956 4413
rect -18990 4345 -18956 4367
rect -18990 4333 -18956 4345
rect -18990 4277 -18956 4295
rect -18990 4261 -18956 4277
rect -18990 4209 -18956 4223
rect -18990 4189 -18956 4209
rect -18990 4141 -18956 4151
rect -18990 4117 -18956 4141
rect -18990 4073 -18956 4079
rect -18990 4045 -18956 4073
rect -18990 4005 -18956 4007
rect -18990 3973 -18956 4005
rect -18990 3903 -18956 3935
rect -18990 3901 -18956 3903
rect -18990 3835 -18956 3863
rect -18990 3829 -18956 3835
rect -18990 3767 -18956 3791
rect -18990 3757 -18956 3767
rect -18990 3699 -18956 3719
rect -18990 3685 -18956 3699
rect -18990 3631 -18956 3647
rect -18990 3613 -18956 3631
rect -18990 3563 -18956 3575
rect -18990 3541 -18956 3563
rect -18990 3495 -18956 3503
rect -18990 3469 -18956 3495
rect -18894 4413 -18860 4439
rect -18894 4405 -18860 4413
rect -18894 4345 -18860 4367
rect -18894 4333 -18860 4345
rect -18894 4277 -18860 4295
rect -18894 4261 -18860 4277
rect -18894 4209 -18860 4223
rect -18894 4189 -18860 4209
rect -18894 4141 -18860 4151
rect -18894 4117 -18860 4141
rect -18894 4073 -18860 4079
rect -18894 4045 -18860 4073
rect -18894 4005 -18860 4007
rect -18894 3973 -18860 4005
rect -18894 3903 -18860 3935
rect -18894 3901 -18860 3903
rect -18894 3835 -18860 3863
rect -18894 3829 -18860 3835
rect -18894 3767 -18860 3791
rect -18894 3757 -18860 3767
rect -18894 3699 -18860 3719
rect -18894 3685 -18860 3699
rect -18894 3631 -18860 3647
rect -18894 3613 -18860 3631
rect -18894 3563 -18860 3575
rect -18894 3541 -18860 3563
rect -18894 3495 -18860 3503
rect -18894 3469 -18860 3495
rect -18798 4413 -18764 4439
rect -18798 4405 -18764 4413
rect -18798 4345 -18764 4367
rect -18798 4333 -18764 4345
rect -18798 4277 -18764 4295
rect -18798 4261 -18764 4277
rect -18798 4209 -18764 4223
rect -18798 4189 -18764 4209
rect -18798 4141 -18764 4151
rect -18798 4117 -18764 4141
rect -18798 4073 -18764 4079
rect -18798 4045 -18764 4073
rect -18798 4005 -18764 4007
rect -18798 3973 -18764 4005
rect -18798 3903 -18764 3935
rect -18798 3901 -18764 3903
rect -18798 3835 -18764 3863
rect -18798 3829 -18764 3835
rect -18798 3767 -18764 3791
rect -18798 3757 -18764 3767
rect -18798 3699 -18764 3719
rect -18798 3685 -18764 3699
rect -18798 3631 -18764 3647
rect -18798 3613 -18764 3631
rect -18798 3563 -18764 3575
rect -18798 3541 -18764 3563
rect -18798 3495 -18764 3503
rect -18798 3469 -18764 3495
rect -18590 4415 -18556 4441
rect -18590 4407 -18556 4415
rect -18590 4347 -18556 4369
rect -18590 4335 -18556 4347
rect -18590 4279 -18556 4297
rect -18590 4263 -18556 4279
rect -18590 4211 -18556 4225
rect -18590 4191 -18556 4211
rect -18590 4143 -18556 4153
rect -18590 4119 -18556 4143
rect -18590 4075 -18556 4081
rect -18590 4047 -18556 4075
rect -18590 4007 -18556 4009
rect -18590 3975 -18556 4007
rect -18590 3905 -18556 3937
rect -18590 3903 -18556 3905
rect -18590 3837 -18556 3865
rect -18590 3831 -18556 3837
rect -18590 3769 -18556 3793
rect -18590 3759 -18556 3769
rect -18590 3701 -18556 3721
rect -18590 3687 -18556 3701
rect -18590 3633 -18556 3649
rect -18590 3615 -18556 3633
rect -18590 3565 -18556 3577
rect -18590 3543 -18556 3565
rect -18590 3497 -18556 3505
rect -18590 3471 -18556 3497
rect -18494 4415 -18460 4441
rect -18494 4407 -18460 4415
rect -18494 4347 -18460 4369
rect -18494 4335 -18460 4347
rect -18494 4279 -18460 4297
rect -18494 4263 -18460 4279
rect -18494 4211 -18460 4225
rect -18494 4191 -18460 4211
rect -18494 4143 -18460 4153
rect -18494 4119 -18460 4143
rect -18494 4075 -18460 4081
rect -18494 4047 -18460 4075
rect -18494 4007 -18460 4009
rect -18494 3975 -18460 4007
rect -18494 3905 -18460 3937
rect -18494 3903 -18460 3905
rect -18494 3837 -18460 3865
rect -18494 3831 -18460 3837
rect -18494 3769 -18460 3793
rect -18494 3759 -18460 3769
rect -18494 3701 -18460 3721
rect -18494 3687 -18460 3701
rect -18494 3633 -18460 3649
rect -18494 3615 -18460 3633
rect -18494 3565 -18460 3577
rect -18494 3543 -18460 3565
rect -18494 3497 -18460 3505
rect -18494 3471 -18460 3497
rect -18398 4415 -18364 4441
rect -18398 4407 -18364 4415
rect -18398 4347 -18364 4369
rect -18398 4335 -18364 4347
rect -18398 4279 -18364 4297
rect -18398 4263 -18364 4279
rect -18398 4211 -18364 4225
rect -18398 4191 -18364 4211
rect -18398 4143 -18364 4153
rect -18398 4119 -18364 4143
rect -18398 4075 -18364 4081
rect -18398 4047 -18364 4075
rect -18398 4007 -18364 4009
rect -18398 3975 -18364 4007
rect -18398 3905 -18364 3937
rect -18398 3903 -18364 3905
rect -18398 3837 -18364 3865
rect -18398 3831 -18364 3837
rect -18398 3769 -18364 3793
rect -18398 3759 -18364 3769
rect -18398 3701 -18364 3721
rect -18398 3687 -18364 3701
rect -18398 3633 -18364 3649
rect -18398 3615 -18364 3633
rect -18398 3565 -18364 3577
rect -18398 3543 -18364 3565
rect -18398 3497 -18364 3505
rect -18398 3471 -18364 3497
rect -18302 4415 -18268 4441
rect -18302 4407 -18268 4415
rect -18302 4347 -18268 4369
rect -18302 4335 -18268 4347
rect -18302 4279 -18268 4297
rect -18302 4263 -18268 4279
rect -18302 4211 -18268 4225
rect -18302 4191 -18268 4211
rect -18302 4143 -18268 4153
rect -18302 4119 -18268 4143
rect -18302 4075 -18268 4081
rect -18302 4047 -18268 4075
rect -18302 4007 -18268 4009
rect -18302 3975 -18268 4007
rect -18302 3905 -18268 3937
rect -18302 3903 -18268 3905
rect -18302 3837 -18268 3865
rect -18302 3831 -18268 3837
rect -18302 3769 -18268 3793
rect -18302 3759 -18268 3769
rect -18302 3701 -18268 3721
rect -18302 3687 -18268 3701
rect -18302 3633 -18268 3649
rect -18302 3615 -18268 3633
rect -18302 3565 -18268 3577
rect -18302 3543 -18268 3565
rect -18302 3497 -18268 3505
rect -18302 3471 -18268 3497
rect -18206 4415 -18172 4441
rect -18206 4407 -18172 4415
rect -18206 4347 -18172 4369
rect -18206 4335 -18172 4347
rect -18206 4279 -18172 4297
rect -18206 4263 -18172 4279
rect -18206 4211 -18172 4225
rect -18206 4191 -18172 4211
rect -18206 4143 -18172 4153
rect -18206 4119 -18172 4143
rect -18206 4075 -18172 4081
rect -18206 4047 -18172 4075
rect -18206 4007 -18172 4009
rect -18206 3975 -18172 4007
rect -18206 3905 -18172 3937
rect -18206 3903 -18172 3905
rect -18206 3837 -18172 3865
rect -18206 3831 -18172 3837
rect -18206 3769 -18172 3793
rect -18206 3759 -18172 3769
rect -18206 3701 -18172 3721
rect -18206 3687 -18172 3701
rect -18206 3633 -18172 3649
rect -18206 3615 -18172 3633
rect -18206 3565 -18172 3577
rect -18206 3543 -18172 3565
rect -18206 3497 -18172 3505
rect -18206 3471 -18172 3497
rect -18110 4415 -18076 4441
rect -18110 4407 -18076 4415
rect -18110 4347 -18076 4369
rect -18110 4335 -18076 4347
rect -18110 4279 -18076 4297
rect -18110 4263 -18076 4279
rect -18110 4211 -18076 4225
rect -18110 4191 -18076 4211
rect -18110 4143 -18076 4153
rect -18110 4119 -18076 4143
rect -18110 4075 -18076 4081
rect -18110 4047 -18076 4075
rect -18110 4007 -18076 4009
rect -18110 3975 -18076 4007
rect -18110 3905 -18076 3937
rect -18110 3903 -18076 3905
rect -18110 3837 -18076 3865
rect -18110 3831 -18076 3837
rect -18110 3769 -18076 3793
rect -18110 3759 -18076 3769
rect -18110 3701 -18076 3721
rect -18110 3687 -18076 3701
rect -18110 3633 -18076 3649
rect -18110 3615 -18076 3633
rect -18110 3565 -18076 3577
rect -18110 3543 -18076 3565
rect -18110 3497 -18076 3505
rect -18110 3471 -18076 3497
rect 1484 4607 1518 4631
rect 1484 4563 1518 4569
rect -16756 4413 -16722 4439
rect -16756 4405 -16722 4413
rect -16756 4345 -16722 4367
rect -16756 4333 -16722 4345
rect -16756 4277 -16722 4295
rect -16756 4261 -16722 4277
rect -16756 4209 -16722 4223
rect -16756 4189 -16722 4209
rect -16756 4141 -16722 4151
rect -16756 4117 -16722 4141
rect -16756 4073 -16722 4079
rect -16756 4045 -16722 4073
rect -16756 4005 -16722 4007
rect -16756 3973 -16722 4005
rect -16756 3903 -16722 3935
rect -16756 3901 -16722 3903
rect -16756 3835 -16722 3863
rect -16756 3829 -16722 3835
rect -16756 3767 -16722 3791
rect -16756 3757 -16722 3767
rect -16756 3699 -16722 3719
rect -16756 3685 -16722 3699
rect -16756 3631 -16722 3647
rect -16756 3613 -16722 3631
rect -16756 3563 -16722 3575
rect -16756 3541 -16722 3563
rect -16756 3495 -16722 3503
rect -16756 3469 -16722 3495
rect -16660 4413 -16626 4439
rect -16660 4405 -16626 4413
rect -16660 4345 -16626 4367
rect -16660 4333 -16626 4345
rect -16660 4277 -16626 4295
rect -16660 4261 -16626 4277
rect -16660 4209 -16626 4223
rect -16660 4189 -16626 4209
rect -16660 4141 -16626 4151
rect -16660 4117 -16626 4141
rect -16660 4073 -16626 4079
rect -16660 4045 -16626 4073
rect -16660 4005 -16626 4007
rect -16660 3973 -16626 4005
rect -16660 3903 -16626 3935
rect -16660 3901 -16626 3903
rect -16660 3835 -16626 3863
rect -16660 3829 -16626 3835
rect -16660 3767 -16626 3791
rect -16660 3757 -16626 3767
rect -16660 3699 -16626 3719
rect -16660 3685 -16626 3699
rect -16660 3631 -16626 3647
rect -16660 3613 -16626 3631
rect -16660 3563 -16626 3575
rect -16660 3541 -16626 3563
rect -16660 3495 -16626 3503
rect -16660 3469 -16626 3495
rect -16564 4413 -16530 4439
rect -16564 4405 -16530 4413
rect -16564 4345 -16530 4367
rect -16564 4333 -16530 4345
rect -16564 4277 -16530 4295
rect -16564 4261 -16530 4277
rect -16564 4209 -16530 4223
rect -16564 4189 -16530 4209
rect -16564 4141 -16530 4151
rect -16564 4117 -16530 4141
rect -16564 4073 -16530 4079
rect -16564 4045 -16530 4073
rect -16564 4005 -16530 4007
rect -16564 3973 -16530 4005
rect -16564 3903 -16530 3935
rect -16564 3901 -16530 3903
rect -16564 3835 -16530 3863
rect -16564 3829 -16530 3835
rect -16564 3767 -16530 3791
rect -16564 3757 -16530 3767
rect -16564 3699 -16530 3719
rect -16564 3685 -16530 3699
rect -16564 3631 -16530 3647
rect -16564 3613 -16530 3631
rect -16564 3563 -16530 3575
rect -16564 3541 -16530 3563
rect -16564 3495 -16530 3503
rect -16564 3469 -16530 3495
rect -16468 4413 -16434 4439
rect -16468 4405 -16434 4413
rect -16468 4345 -16434 4367
rect -16468 4333 -16434 4345
rect -16468 4277 -16434 4295
rect -16468 4261 -16434 4277
rect -16468 4209 -16434 4223
rect -16468 4189 -16434 4209
rect -16468 4141 -16434 4151
rect -16468 4117 -16434 4141
rect -16468 4073 -16434 4079
rect -16468 4045 -16434 4073
rect -16468 4005 -16434 4007
rect -16468 3973 -16434 4005
rect -16468 3903 -16434 3935
rect -16468 3901 -16434 3903
rect -16468 3835 -16434 3863
rect -16468 3829 -16434 3835
rect -16468 3767 -16434 3791
rect -16468 3757 -16434 3767
rect -16468 3699 -16434 3719
rect -16468 3685 -16434 3699
rect -16468 3631 -16434 3647
rect -16468 3613 -16434 3631
rect -16468 3563 -16434 3575
rect -16468 3541 -16434 3563
rect -16468 3495 -16434 3503
rect -16468 3469 -16434 3495
rect -16372 4413 -16338 4439
rect -16372 4405 -16338 4413
rect -16372 4345 -16338 4367
rect -16372 4333 -16338 4345
rect -16372 4277 -16338 4295
rect -16372 4261 -16338 4277
rect -16372 4209 -16338 4223
rect -16372 4189 -16338 4209
rect -16372 4141 -16338 4151
rect -16372 4117 -16338 4141
rect -16372 4073 -16338 4079
rect -16372 4045 -16338 4073
rect -16372 4005 -16338 4007
rect -16372 3973 -16338 4005
rect -16372 3903 -16338 3935
rect -16372 3901 -16338 3903
rect -16372 3835 -16338 3863
rect -16372 3829 -16338 3835
rect -16372 3767 -16338 3791
rect -16372 3757 -16338 3767
rect -16372 3699 -16338 3719
rect -16372 3685 -16338 3699
rect -16372 3631 -16338 3647
rect -16372 3613 -16338 3631
rect -16372 3563 -16338 3575
rect -16372 3541 -16338 3563
rect -16372 3495 -16338 3503
rect -16372 3469 -16338 3495
rect -16276 4413 -16242 4439
rect -16276 4405 -16242 4413
rect -16276 4345 -16242 4367
rect -16276 4333 -16242 4345
rect -16276 4277 -16242 4295
rect -16276 4261 -16242 4277
rect -16276 4209 -16242 4223
rect -16276 4189 -16242 4209
rect -16276 4141 -16242 4151
rect -16276 4117 -16242 4141
rect -16276 4073 -16242 4079
rect -16276 4045 -16242 4073
rect -16276 4005 -16242 4007
rect -16276 3973 -16242 4005
rect -16276 3903 -16242 3935
rect -16276 3901 -16242 3903
rect -16276 3835 -16242 3863
rect -16276 3829 -16242 3835
rect -16276 3767 -16242 3791
rect -16276 3757 -16242 3767
rect -16276 3699 -16242 3719
rect -16276 3685 -16242 3699
rect -16276 3631 -16242 3647
rect -16276 3613 -16242 3631
rect -16276 3563 -16242 3575
rect -16276 3541 -16242 3563
rect -16276 3495 -16242 3503
rect -16276 3469 -16242 3495
rect -16180 4413 -16146 4439
rect -16180 4405 -16146 4413
rect -16180 4345 -16146 4367
rect -16180 4333 -16146 4345
rect -16180 4277 -16146 4295
rect -16180 4261 -16146 4277
rect -16180 4209 -16146 4223
rect -16180 4189 -16146 4209
rect -16180 4141 -16146 4151
rect -16180 4117 -16146 4141
rect -16180 4073 -16146 4079
rect -16180 4045 -16146 4073
rect -16180 4005 -16146 4007
rect -16180 3973 -16146 4005
rect -16180 3903 -16146 3935
rect -16180 3901 -16146 3903
rect -16180 3835 -16146 3863
rect -16180 3829 -16146 3835
rect -16180 3767 -16146 3791
rect -16180 3757 -16146 3767
rect -16180 3699 -16146 3719
rect -16180 3685 -16146 3699
rect -16180 3631 -16146 3647
rect -16180 3613 -16146 3631
rect -16180 3563 -16146 3575
rect -16180 3541 -16146 3563
rect -16180 3495 -16146 3503
rect -16180 3469 -16146 3495
rect -16084 4413 -16050 4439
rect -16084 4405 -16050 4413
rect -16084 4345 -16050 4367
rect -16084 4333 -16050 4345
rect -16084 4277 -16050 4295
rect -16084 4261 -16050 4277
rect -16084 4209 -16050 4223
rect -16084 4189 -16050 4209
rect -16084 4141 -16050 4151
rect -16084 4117 -16050 4141
rect -16084 4073 -16050 4079
rect -16084 4045 -16050 4073
rect -16084 4005 -16050 4007
rect -16084 3973 -16050 4005
rect -16084 3903 -16050 3935
rect -16084 3901 -16050 3903
rect -16084 3835 -16050 3863
rect -16084 3829 -16050 3835
rect -16084 3767 -16050 3791
rect -16084 3757 -16050 3767
rect -16084 3699 -16050 3719
rect -16084 3685 -16050 3699
rect -16084 3631 -16050 3647
rect -16084 3613 -16050 3631
rect -16084 3563 -16050 3575
rect -16084 3541 -16050 3563
rect -16084 3495 -16050 3503
rect -16084 3469 -16050 3495
rect -15988 4413 -15954 4439
rect -15988 4405 -15954 4413
rect -15988 4345 -15954 4367
rect -15988 4333 -15954 4345
rect -15988 4277 -15954 4295
rect -15988 4261 -15954 4277
rect -15988 4209 -15954 4223
rect -15988 4189 -15954 4209
rect -15988 4141 -15954 4151
rect -15988 4117 -15954 4141
rect -15988 4073 -15954 4079
rect -15988 4045 -15954 4073
rect -15988 4005 -15954 4007
rect -15988 3973 -15954 4005
rect -15988 3903 -15954 3935
rect -15988 3901 -15954 3903
rect -15988 3835 -15954 3863
rect -15988 3829 -15954 3835
rect -15988 3767 -15954 3791
rect -15988 3757 -15954 3767
rect -15988 3699 -15954 3719
rect -15988 3685 -15954 3699
rect -15988 3631 -15954 3647
rect -15988 3613 -15954 3631
rect -15988 3563 -15954 3575
rect -15988 3541 -15954 3563
rect -15988 3495 -15954 3503
rect -15988 3469 -15954 3495
rect -15892 4413 -15858 4439
rect -15892 4405 -15858 4413
rect -15892 4345 -15858 4367
rect -15892 4333 -15858 4345
rect -15892 4277 -15858 4295
rect -15892 4261 -15858 4277
rect -15892 4209 -15858 4223
rect -15892 4189 -15858 4209
rect -15892 4141 -15858 4151
rect -15892 4117 -15858 4141
rect -15892 4073 -15858 4079
rect -15892 4045 -15858 4073
rect -15892 4005 -15858 4007
rect -15892 3973 -15858 4005
rect -15892 3903 -15858 3935
rect -15892 3901 -15858 3903
rect -15892 3835 -15858 3863
rect -15892 3829 -15858 3835
rect -15892 3767 -15858 3791
rect -15892 3757 -15858 3767
rect -15892 3699 -15858 3719
rect -15892 3685 -15858 3699
rect -15892 3631 -15858 3647
rect -15892 3613 -15858 3631
rect -15892 3563 -15858 3575
rect -15892 3541 -15858 3563
rect -15892 3495 -15858 3503
rect -15892 3469 -15858 3495
rect -15796 4413 -15762 4439
rect -15796 4405 -15762 4413
rect -15796 4345 -15762 4367
rect -15796 4333 -15762 4345
rect -15796 4277 -15762 4295
rect -15796 4261 -15762 4277
rect -15796 4209 -15762 4223
rect -15796 4189 -15762 4209
rect -15796 4141 -15762 4151
rect -15796 4117 -15762 4141
rect -15796 4073 -15762 4079
rect -15796 4045 -15762 4073
rect -15796 4005 -15762 4007
rect -15796 3973 -15762 4005
rect -15796 3903 -15762 3935
rect -15796 3901 -15762 3903
rect -15796 3835 -15762 3863
rect -15796 3829 -15762 3835
rect -15796 3767 -15762 3791
rect -15796 3757 -15762 3767
rect -15796 3699 -15762 3719
rect -15796 3685 -15762 3699
rect -15796 3631 -15762 3647
rect -15796 3613 -15762 3631
rect -15796 3563 -15762 3575
rect -15796 3541 -15762 3563
rect -15796 3495 -15762 3503
rect -15796 3469 -15762 3495
rect -15700 4413 -15666 4439
rect -15700 4405 -15666 4413
rect -15700 4345 -15666 4367
rect -15700 4333 -15666 4345
rect -15700 4277 -15666 4295
rect -15700 4261 -15666 4277
rect -15700 4209 -15666 4223
rect -15700 4189 -15666 4209
rect -15700 4141 -15666 4151
rect -15700 4117 -15666 4141
rect -15700 4073 -15666 4079
rect -15700 4045 -15666 4073
rect -15700 4005 -15666 4007
rect -15700 3973 -15666 4005
rect -15700 3903 -15666 3935
rect -15700 3901 -15666 3903
rect -15700 3835 -15666 3863
rect -15700 3829 -15666 3835
rect -15700 3767 -15666 3791
rect -15700 3757 -15666 3767
rect -15700 3699 -15666 3719
rect -15700 3685 -15666 3699
rect -15700 3631 -15666 3647
rect -15700 3613 -15666 3631
rect -15700 3563 -15666 3575
rect -15700 3541 -15666 3563
rect -15700 3495 -15666 3503
rect -15700 3469 -15666 3495
rect -15604 4413 -15570 4439
rect -15604 4405 -15570 4413
rect -15604 4345 -15570 4367
rect -15604 4333 -15570 4345
rect -15604 4277 -15570 4295
rect -15604 4261 -15570 4277
rect -15604 4209 -15570 4223
rect -15604 4189 -15570 4209
rect -15604 4141 -15570 4151
rect -15604 4117 -15570 4141
rect -15604 4073 -15570 4079
rect -15604 4045 -15570 4073
rect -15604 4005 -15570 4007
rect -15604 3973 -15570 4005
rect -15604 3903 -15570 3935
rect -15604 3901 -15570 3903
rect -15604 3835 -15570 3863
rect -15604 3829 -15570 3835
rect -15604 3767 -15570 3791
rect -15604 3757 -15570 3767
rect -15604 3699 -15570 3719
rect -15604 3685 -15570 3699
rect -15604 3631 -15570 3647
rect -15604 3613 -15570 3631
rect -15604 3563 -15570 3575
rect -15604 3541 -15570 3563
rect -15604 3495 -15570 3503
rect -15604 3469 -15570 3495
rect -15508 4413 -15474 4439
rect -15508 4405 -15474 4413
rect -15508 4345 -15474 4367
rect -15508 4333 -15474 4345
rect -15508 4277 -15474 4295
rect -15508 4261 -15474 4277
rect -15508 4209 -15474 4223
rect -15508 4189 -15474 4209
rect -15508 4141 -15474 4151
rect -15508 4117 -15474 4141
rect -15508 4073 -15474 4079
rect -15508 4045 -15474 4073
rect -15508 4005 -15474 4007
rect -15508 3973 -15474 4005
rect -15508 3903 -15474 3935
rect -15508 3901 -15474 3903
rect -15508 3835 -15474 3863
rect -15508 3829 -15474 3835
rect -15508 3767 -15474 3791
rect -15508 3757 -15474 3767
rect -15508 3699 -15474 3719
rect -15508 3685 -15474 3699
rect -15508 3631 -15474 3647
rect -15508 3613 -15474 3631
rect -15508 3563 -15474 3575
rect -15508 3541 -15474 3563
rect -15508 3495 -15474 3503
rect -15508 3469 -15474 3495
rect -15412 4413 -15378 4439
rect -15412 4405 -15378 4413
rect -15412 4345 -15378 4367
rect -15412 4333 -15378 4345
rect -15412 4277 -15378 4295
rect -15412 4261 -15378 4277
rect -15412 4209 -15378 4223
rect -15412 4189 -15378 4209
rect -15412 4141 -15378 4151
rect -15412 4117 -15378 4141
rect -15412 4073 -15378 4079
rect -15412 4045 -15378 4073
rect -15412 4005 -15378 4007
rect -15412 3973 -15378 4005
rect -15412 3903 -15378 3935
rect -15412 3901 -15378 3903
rect -15412 3835 -15378 3863
rect -15412 3829 -15378 3835
rect -15412 3767 -15378 3791
rect -15412 3757 -15378 3767
rect -15412 3699 -15378 3719
rect -15412 3685 -15378 3699
rect -15412 3631 -15378 3647
rect -15412 3613 -15378 3631
rect -15412 3563 -15378 3575
rect -15412 3541 -15378 3563
rect -15412 3495 -15378 3503
rect -15412 3469 -15378 3495
rect -15316 4413 -15282 4439
rect -15316 4405 -15282 4413
rect -15316 4345 -15282 4367
rect -15316 4333 -15282 4345
rect -15316 4277 -15282 4295
rect -15316 4261 -15282 4277
rect -15316 4209 -15282 4223
rect -15316 4189 -15282 4209
rect -15316 4141 -15282 4151
rect -15316 4117 -15282 4141
rect -15316 4073 -15282 4079
rect -15316 4045 -15282 4073
rect -15316 4005 -15282 4007
rect -15316 3973 -15282 4005
rect -15316 3903 -15282 3935
rect -15316 3901 -15282 3903
rect -15316 3835 -15282 3863
rect -15316 3829 -15282 3835
rect -15316 3767 -15282 3791
rect -15316 3757 -15282 3767
rect -15316 3699 -15282 3719
rect -15316 3685 -15282 3699
rect -15316 3631 -15282 3647
rect -15316 3613 -15282 3631
rect -15316 3563 -15282 3575
rect -15316 3541 -15282 3563
rect -15316 3495 -15282 3503
rect -15316 3469 -15282 3495
rect -15220 4413 -15186 4439
rect -15220 4405 -15186 4413
rect -15220 4345 -15186 4367
rect -15220 4333 -15186 4345
rect -15220 4277 -15186 4295
rect -15220 4261 -15186 4277
rect -15220 4209 -15186 4223
rect -15220 4189 -15186 4209
rect -15220 4141 -15186 4151
rect -15220 4117 -15186 4141
rect -15220 4073 -15186 4079
rect -15220 4045 -15186 4073
rect -15220 4005 -15186 4007
rect -15220 3973 -15186 4005
rect -15220 3903 -15186 3935
rect -15220 3901 -15186 3903
rect -15220 3835 -15186 3863
rect -15220 3829 -15186 3835
rect -15220 3767 -15186 3791
rect -15220 3757 -15186 3767
rect -15220 3699 -15186 3719
rect -15220 3685 -15186 3699
rect -15220 3631 -15186 3647
rect -15220 3613 -15186 3631
rect -15220 3563 -15186 3575
rect -15220 3541 -15186 3563
rect -15220 3495 -15186 3503
rect -15220 3469 -15186 3495
rect -15124 4413 -15090 4439
rect -15124 4405 -15090 4413
rect -15124 4345 -15090 4367
rect -15124 4333 -15090 4345
rect -15124 4277 -15090 4295
rect -15124 4261 -15090 4277
rect -15124 4209 -15090 4223
rect -15124 4189 -15090 4209
rect -15124 4141 -15090 4151
rect -15124 4117 -15090 4141
rect -15124 4073 -15090 4079
rect -15124 4045 -15090 4073
rect -15124 4005 -15090 4007
rect -15124 3973 -15090 4005
rect -15124 3903 -15090 3935
rect -15124 3901 -15090 3903
rect -15124 3835 -15090 3863
rect -15124 3829 -15090 3835
rect -15124 3767 -15090 3791
rect -15124 3757 -15090 3767
rect -15124 3699 -15090 3719
rect -15124 3685 -15090 3699
rect -15124 3631 -15090 3647
rect -15124 3613 -15090 3631
rect -15124 3563 -15090 3575
rect -15124 3541 -15090 3563
rect -15124 3495 -15090 3503
rect -15124 3469 -15090 3495
rect -15028 4413 -14994 4439
rect -15028 4405 -14994 4413
rect -15028 4345 -14994 4367
rect -15028 4333 -14994 4345
rect -15028 4277 -14994 4295
rect -15028 4261 -14994 4277
rect -15028 4209 -14994 4223
rect -15028 4189 -14994 4209
rect -15028 4141 -14994 4151
rect -15028 4117 -14994 4141
rect -15028 4073 -14994 4079
rect -15028 4045 -14994 4073
rect -15028 4005 -14994 4007
rect -15028 3973 -14994 4005
rect -15028 3903 -14994 3935
rect -15028 3901 -14994 3903
rect -15028 3835 -14994 3863
rect -15028 3829 -14994 3835
rect -15028 3767 -14994 3791
rect -15028 3757 -14994 3767
rect -15028 3699 -14994 3719
rect -15028 3685 -14994 3699
rect -15028 3631 -14994 3647
rect -15028 3613 -14994 3631
rect -15028 3563 -14994 3575
rect -15028 3541 -14994 3563
rect -15028 3495 -14994 3503
rect -15028 3469 -14994 3495
rect -14932 4413 -14898 4439
rect -14932 4405 -14898 4413
rect -14932 4345 -14898 4367
rect -14932 4333 -14898 4345
rect -14932 4277 -14898 4295
rect -14932 4261 -14898 4277
rect -14932 4209 -14898 4223
rect -14932 4189 -14898 4209
rect -14932 4141 -14898 4151
rect -14932 4117 -14898 4141
rect -14932 4073 -14898 4079
rect -14932 4045 -14898 4073
rect -14932 4005 -14898 4007
rect -14932 3973 -14898 4005
rect -14932 3903 -14898 3935
rect -14932 3901 -14898 3903
rect -14932 3835 -14898 3863
rect -14932 3829 -14898 3835
rect -14932 3767 -14898 3791
rect -14932 3757 -14898 3767
rect -14932 3699 -14898 3719
rect -14932 3685 -14898 3699
rect -14932 3631 -14898 3647
rect -14932 3613 -14898 3631
rect -14932 3563 -14898 3575
rect -14932 3541 -14898 3563
rect -14932 3495 -14898 3503
rect -14932 3469 -14898 3495
rect -14836 4413 -14802 4439
rect -14836 4405 -14802 4413
rect -14836 4345 -14802 4367
rect -14836 4333 -14802 4345
rect -14836 4277 -14802 4295
rect -14836 4261 -14802 4277
rect -14836 4209 -14802 4223
rect -14836 4189 -14802 4209
rect -14836 4141 -14802 4151
rect -14836 4117 -14802 4141
rect -14836 4073 -14802 4079
rect -14836 4045 -14802 4073
rect -14836 4005 -14802 4007
rect -14836 3973 -14802 4005
rect -14836 3903 -14802 3935
rect -14836 3901 -14802 3903
rect -14836 3835 -14802 3863
rect -14836 3829 -14802 3835
rect -14836 3767 -14802 3791
rect -14836 3757 -14802 3767
rect -14836 3699 -14802 3719
rect -14836 3685 -14802 3699
rect -14836 3631 -14802 3647
rect -14836 3613 -14802 3631
rect -14836 3563 -14802 3575
rect -14836 3541 -14802 3563
rect -14836 3495 -14802 3503
rect -14836 3469 -14802 3495
rect -14612 4419 -14578 4445
rect -14612 4411 -14578 4419
rect -14612 4351 -14578 4373
rect -14612 4339 -14578 4351
rect -14612 4283 -14578 4301
rect -14612 4267 -14578 4283
rect -14612 4215 -14578 4229
rect -14612 4195 -14578 4215
rect -14612 4147 -14578 4157
rect -14612 4123 -14578 4147
rect -14612 4079 -14578 4085
rect -14612 4051 -14578 4079
rect -14612 4011 -14578 4013
rect -14612 3979 -14578 4011
rect -14612 3909 -14578 3941
rect -14612 3907 -14578 3909
rect -14612 3841 -14578 3869
rect -14612 3835 -14578 3841
rect -14612 3773 -14578 3797
rect -14612 3763 -14578 3773
rect -14612 3705 -14578 3725
rect -14612 3691 -14578 3705
rect -14612 3637 -14578 3653
rect -14612 3619 -14578 3637
rect -14612 3569 -14578 3581
rect -14612 3547 -14578 3569
rect -14612 3501 -14578 3509
rect -14612 3475 -14578 3501
rect -14516 4419 -14482 4445
rect -14516 4411 -14482 4419
rect -14516 4351 -14482 4373
rect -14516 4339 -14482 4351
rect -14516 4283 -14482 4301
rect -14516 4267 -14482 4283
rect -14516 4215 -14482 4229
rect -14516 4195 -14482 4215
rect -14516 4147 -14482 4157
rect -14516 4123 -14482 4147
rect -14516 4079 -14482 4085
rect -14516 4051 -14482 4079
rect -14516 4011 -14482 4013
rect -14516 3979 -14482 4011
rect -14516 3909 -14482 3941
rect -14516 3907 -14482 3909
rect -14516 3841 -14482 3869
rect -14516 3835 -14482 3841
rect -14516 3773 -14482 3797
rect -14516 3763 -14482 3773
rect -14516 3705 -14482 3725
rect -14516 3691 -14482 3705
rect -14516 3637 -14482 3653
rect -14516 3619 -14482 3637
rect -14516 3569 -14482 3581
rect -14516 3547 -14482 3569
rect -14516 3501 -14482 3509
rect -14516 3475 -14482 3501
rect -14420 4419 -14386 4445
rect -14420 4411 -14386 4419
rect -14420 4351 -14386 4373
rect -14420 4339 -14386 4351
rect -14420 4283 -14386 4301
rect -14420 4267 -14386 4283
rect -14420 4215 -14386 4229
rect -14420 4195 -14386 4215
rect -14420 4147 -14386 4157
rect -14420 4123 -14386 4147
rect -14420 4079 -14386 4085
rect -14420 4051 -14386 4079
rect -14420 4011 -14386 4013
rect -14420 3979 -14386 4011
rect -14420 3909 -14386 3941
rect -14420 3907 -14386 3909
rect -14420 3841 -14386 3869
rect -14420 3835 -14386 3841
rect -14420 3773 -14386 3797
rect -14420 3763 -14386 3773
rect -14420 3705 -14386 3725
rect -14420 3691 -14386 3705
rect -14420 3637 -14386 3653
rect -14420 3619 -14386 3637
rect -14420 3569 -14386 3581
rect -14420 3547 -14386 3569
rect -14420 3501 -14386 3509
rect -14420 3475 -14386 3501
rect -14324 4419 -14290 4445
rect -14324 4411 -14290 4419
rect -14324 4351 -14290 4373
rect -14324 4339 -14290 4351
rect -14324 4283 -14290 4301
rect -14324 4267 -14290 4283
rect -14324 4215 -14290 4229
rect -14324 4195 -14290 4215
rect -14324 4147 -14290 4157
rect -14324 4123 -14290 4147
rect -14324 4079 -14290 4085
rect -14324 4051 -14290 4079
rect -14324 4011 -14290 4013
rect -14324 3979 -14290 4011
rect -14324 3909 -14290 3941
rect -14324 3907 -14290 3909
rect -14324 3841 -14290 3869
rect -14324 3835 -14290 3841
rect -14324 3773 -14290 3797
rect -14324 3763 -14290 3773
rect -14324 3705 -14290 3725
rect -14324 3691 -14290 3705
rect -14324 3637 -14290 3653
rect -14324 3619 -14290 3637
rect -14324 3569 -14290 3581
rect -14324 3547 -14290 3569
rect -14324 3501 -14290 3509
rect -14324 3475 -14290 3501
rect -14228 4419 -14194 4445
rect -14228 4411 -14194 4419
rect -14228 4351 -14194 4373
rect -14228 4339 -14194 4351
rect -14228 4283 -14194 4301
rect -14228 4267 -14194 4283
rect -14228 4215 -14194 4229
rect -14228 4195 -14194 4215
rect -14228 4147 -14194 4157
rect -14228 4123 -14194 4147
rect -14228 4079 -14194 4085
rect -14228 4051 -14194 4079
rect -14228 4011 -14194 4013
rect -14228 3979 -14194 4011
rect -14228 3909 -14194 3941
rect -14228 3907 -14194 3909
rect -14228 3841 -14194 3869
rect -14228 3835 -14194 3841
rect -14228 3773 -14194 3797
rect -14228 3763 -14194 3773
rect -14228 3705 -14194 3725
rect -14228 3691 -14194 3705
rect -14228 3637 -14194 3653
rect -14228 3619 -14194 3637
rect -14228 3569 -14194 3581
rect -14228 3547 -14194 3569
rect -14228 3501 -14194 3509
rect -14228 3475 -14194 3501
rect -14132 4419 -14098 4445
rect -14132 4411 -14098 4419
rect -14132 4351 -14098 4373
rect -14132 4339 -14098 4351
rect -14132 4283 -14098 4301
rect -14132 4267 -14098 4283
rect -14132 4215 -14098 4229
rect -14132 4195 -14098 4215
rect -14132 4147 -14098 4157
rect -14132 4123 -14098 4147
rect -14132 4079 -14098 4085
rect -14132 4051 -14098 4079
rect -14132 4011 -14098 4013
rect -14132 3979 -14098 4011
rect -14132 3909 -14098 3941
rect -14132 3907 -14098 3909
rect -14132 3841 -14098 3869
rect -14132 3835 -14098 3841
rect -14132 3773 -14098 3797
rect -14132 3763 -14098 3773
rect -14132 3705 -14098 3725
rect -14132 3691 -14098 3705
rect -14132 3637 -14098 3653
rect -14132 3619 -14098 3637
rect -14132 3569 -14098 3581
rect -14132 3547 -14098 3569
rect -14132 3501 -14098 3509
rect -14132 3475 -14098 3501
rect -14036 4419 -14002 4445
rect -14036 4411 -14002 4419
rect -14036 4351 -14002 4373
rect -14036 4339 -14002 4351
rect -14036 4283 -14002 4301
rect -14036 4267 -14002 4283
rect -14036 4215 -14002 4229
rect -14036 4195 -14002 4215
rect -14036 4147 -14002 4157
rect -14036 4123 -14002 4147
rect -14036 4079 -14002 4085
rect -14036 4051 -14002 4079
rect -14036 4011 -14002 4013
rect -14036 3979 -14002 4011
rect -14036 3909 -14002 3941
rect -14036 3907 -14002 3909
rect -14036 3841 -14002 3869
rect -14036 3835 -14002 3841
rect -14036 3773 -14002 3797
rect -14036 3763 -14002 3773
rect -14036 3705 -14002 3725
rect -14036 3691 -14002 3705
rect -14036 3637 -14002 3653
rect -14036 3619 -14002 3637
rect -14036 3569 -14002 3581
rect -14036 3547 -14002 3569
rect -14036 3501 -14002 3509
rect -14036 3475 -14002 3501
rect -13940 4419 -13906 4445
rect -13940 4411 -13906 4419
rect -13940 4351 -13906 4373
rect -13940 4339 -13906 4351
rect -13940 4283 -13906 4301
rect -13940 4267 -13906 4283
rect -13940 4215 -13906 4229
rect -13940 4195 -13906 4215
rect -13940 4147 -13906 4157
rect -13940 4123 -13906 4147
rect -13940 4079 -13906 4085
rect -13940 4051 -13906 4079
rect -13940 4011 -13906 4013
rect -13940 3979 -13906 4011
rect -13940 3909 -13906 3941
rect -13940 3907 -13906 3909
rect -13940 3841 -13906 3869
rect -13940 3835 -13906 3841
rect -13940 3773 -13906 3797
rect -13940 3763 -13906 3773
rect -13940 3705 -13906 3725
rect -13940 3691 -13906 3705
rect -13940 3637 -13906 3653
rect -13940 3619 -13906 3637
rect -13940 3569 -13906 3581
rect -13940 3547 -13906 3569
rect -13940 3501 -13906 3509
rect -13940 3475 -13906 3501
rect -13844 4419 -13810 4445
rect -13844 4411 -13810 4419
rect -13844 4351 -13810 4373
rect -13844 4339 -13810 4351
rect -13844 4283 -13810 4301
rect -13844 4267 -13810 4283
rect -13844 4215 -13810 4229
rect -13844 4195 -13810 4215
rect -13844 4147 -13810 4157
rect -13844 4123 -13810 4147
rect -13844 4079 -13810 4085
rect -13844 4051 -13810 4079
rect -13844 4011 -13810 4013
rect -13844 3979 -13810 4011
rect -13844 3909 -13810 3941
rect -13844 3907 -13810 3909
rect -13844 3841 -13810 3869
rect -13844 3835 -13810 3841
rect -13844 3773 -13810 3797
rect -13844 3763 -13810 3773
rect -13844 3705 -13810 3725
rect -13844 3691 -13810 3705
rect -13844 3637 -13810 3653
rect -13844 3619 -13810 3637
rect -13844 3569 -13810 3581
rect -13844 3547 -13810 3569
rect -13844 3501 -13810 3509
rect -13844 3475 -13810 3501
rect -13748 4419 -13714 4445
rect -13748 4411 -13714 4419
rect -13748 4351 -13714 4373
rect -13748 4339 -13714 4351
rect -13748 4283 -13714 4301
rect -13748 4267 -13714 4283
rect -13748 4215 -13714 4229
rect -13748 4195 -13714 4215
rect -13748 4147 -13714 4157
rect -13748 4123 -13714 4147
rect -13748 4079 -13714 4085
rect -13748 4051 -13714 4079
rect -13748 4011 -13714 4013
rect -13748 3979 -13714 4011
rect -13748 3909 -13714 3941
rect -13748 3907 -13714 3909
rect -13748 3841 -13714 3869
rect -13748 3835 -13714 3841
rect -13748 3773 -13714 3797
rect -13748 3763 -13714 3773
rect -13748 3705 -13714 3725
rect -13748 3691 -13714 3705
rect -13748 3637 -13714 3653
rect -13748 3619 -13714 3637
rect -13748 3569 -13714 3581
rect -13748 3547 -13714 3569
rect -13748 3501 -13714 3509
rect -13748 3475 -13714 3501
rect -13652 4419 -13618 4445
rect -13652 4411 -13618 4419
rect -13652 4351 -13618 4373
rect -13652 4339 -13618 4351
rect -13652 4283 -13618 4301
rect -13652 4267 -13618 4283
rect -13652 4215 -13618 4229
rect -13652 4195 -13618 4215
rect -13652 4147 -13618 4157
rect -13652 4123 -13618 4147
rect -13652 4079 -13618 4085
rect -13652 4051 -13618 4079
rect -13652 4011 -13618 4013
rect -13652 3979 -13618 4011
rect -13652 3909 -13618 3941
rect -13652 3907 -13618 3909
rect -13652 3841 -13618 3869
rect -13652 3835 -13618 3841
rect -13652 3773 -13618 3797
rect -13652 3763 -13618 3773
rect -13652 3705 -13618 3725
rect -13652 3691 -13618 3705
rect -13652 3637 -13618 3653
rect -13652 3619 -13618 3637
rect -13652 3569 -13618 3581
rect -13652 3547 -13618 3569
rect -13652 3501 -13618 3509
rect -13652 3475 -13618 3501
rect -13556 4419 -13522 4445
rect -13556 4411 -13522 4419
rect -13556 4351 -13522 4373
rect -13556 4339 -13522 4351
rect -13556 4283 -13522 4301
rect -13556 4267 -13522 4283
rect -13556 4215 -13522 4229
rect -13556 4195 -13522 4215
rect -13556 4147 -13522 4157
rect -13556 4123 -13522 4147
rect -13556 4079 -13522 4085
rect -13556 4051 -13522 4079
rect -13556 4011 -13522 4013
rect -13556 3979 -13522 4011
rect -13556 3909 -13522 3941
rect -13556 3907 -13522 3909
rect -13556 3841 -13522 3869
rect -13556 3835 -13522 3841
rect -13556 3773 -13522 3797
rect -13556 3763 -13522 3773
rect -13556 3705 -13522 3725
rect -13556 3691 -13522 3705
rect -13556 3637 -13522 3653
rect -13556 3619 -13522 3637
rect -13556 3569 -13522 3581
rect -13556 3547 -13522 3569
rect -13556 3501 -13522 3509
rect -13556 3475 -13522 3501
rect -13460 4419 -13426 4445
rect -13460 4411 -13426 4419
rect -13460 4351 -13426 4373
rect -13460 4339 -13426 4351
rect -13460 4283 -13426 4301
rect -13460 4267 -13426 4283
rect -13460 4215 -13426 4229
rect -13460 4195 -13426 4215
rect -13460 4147 -13426 4157
rect -13460 4123 -13426 4147
rect -13460 4079 -13426 4085
rect -13460 4051 -13426 4079
rect -13460 4011 -13426 4013
rect -13460 3979 -13426 4011
rect -13460 3909 -13426 3941
rect -13460 3907 -13426 3909
rect -13460 3841 -13426 3869
rect -13460 3835 -13426 3841
rect -13460 3773 -13426 3797
rect -13460 3763 -13426 3773
rect -13460 3705 -13426 3725
rect -13460 3691 -13426 3705
rect -13460 3637 -13426 3653
rect -13460 3619 -13426 3637
rect -13460 3569 -13426 3581
rect -13460 3547 -13426 3569
rect -13460 3501 -13426 3509
rect -13460 3475 -13426 3501
rect -13364 4419 -13330 4445
rect -13364 4411 -13330 4419
rect -13364 4351 -13330 4373
rect -13364 4339 -13330 4351
rect -13364 4283 -13330 4301
rect -13364 4267 -13330 4283
rect -13364 4215 -13330 4229
rect -13364 4195 -13330 4215
rect -13364 4147 -13330 4157
rect -13364 4123 -13330 4147
rect -13364 4079 -13330 4085
rect -13364 4051 -13330 4079
rect -13364 4011 -13330 4013
rect -13364 3979 -13330 4011
rect -13364 3909 -13330 3941
rect -13364 3907 -13330 3909
rect -13364 3841 -13330 3869
rect -13364 3835 -13330 3841
rect -13364 3773 -13330 3797
rect -13364 3763 -13330 3773
rect -13364 3705 -13330 3725
rect -13364 3691 -13330 3705
rect -13364 3637 -13330 3653
rect -13364 3619 -13330 3637
rect -13364 3569 -13330 3581
rect -13364 3547 -13330 3569
rect -13364 3501 -13330 3509
rect -13364 3475 -13330 3501
rect -13268 4419 -13234 4445
rect -13268 4411 -13234 4419
rect -13268 4351 -13234 4373
rect -13268 4339 -13234 4351
rect -13268 4283 -13234 4301
rect -13268 4267 -13234 4283
rect -13268 4215 -13234 4229
rect -13268 4195 -13234 4215
rect -13268 4147 -13234 4157
rect -13268 4123 -13234 4147
rect -13268 4079 -13234 4085
rect -13268 4051 -13234 4079
rect -13268 4011 -13234 4013
rect -13268 3979 -13234 4011
rect -13268 3909 -13234 3941
rect -13268 3907 -13234 3909
rect -13268 3841 -13234 3869
rect -13268 3835 -13234 3841
rect -13268 3773 -13234 3797
rect -13268 3763 -13234 3773
rect -13268 3705 -13234 3725
rect -13268 3691 -13234 3705
rect -13268 3637 -13234 3653
rect -13268 3619 -13234 3637
rect -13268 3569 -13234 3581
rect -13268 3547 -13234 3569
rect -13268 3501 -13234 3509
rect -13268 3475 -13234 3501
rect -13172 4419 -13138 4445
rect -13172 4411 -13138 4419
rect -13172 4351 -13138 4373
rect -13172 4339 -13138 4351
rect -13172 4283 -13138 4301
rect -13172 4267 -13138 4283
rect -13172 4215 -13138 4229
rect -13172 4195 -13138 4215
rect -13172 4147 -13138 4157
rect -13172 4123 -13138 4147
rect -13172 4079 -13138 4085
rect -13172 4051 -13138 4079
rect -13172 4011 -13138 4013
rect -13172 3979 -13138 4011
rect -13172 3909 -13138 3941
rect -13172 3907 -13138 3909
rect -13172 3841 -13138 3869
rect -13172 3835 -13138 3841
rect -13172 3773 -13138 3797
rect -13172 3763 -13138 3773
rect -13172 3705 -13138 3725
rect -13172 3691 -13138 3705
rect -13172 3637 -13138 3653
rect -13172 3619 -13138 3637
rect -13172 3569 -13138 3581
rect -13172 3547 -13138 3569
rect -13172 3501 -13138 3509
rect -13172 3475 -13138 3501
rect -12928 4425 -12894 4451
rect -12928 4417 -12894 4425
rect -12928 4357 -12894 4379
rect -12928 4345 -12894 4357
rect -12928 4289 -12894 4307
rect -12928 4273 -12894 4289
rect -12928 4221 -12894 4235
rect -12928 4201 -12894 4221
rect -12928 4153 -12894 4163
rect -12928 4129 -12894 4153
rect -12928 4085 -12894 4091
rect -12928 4057 -12894 4085
rect -12928 4017 -12894 4019
rect -12928 3985 -12894 4017
rect -12928 3915 -12894 3947
rect -12928 3913 -12894 3915
rect -12928 3847 -12894 3875
rect -12928 3841 -12894 3847
rect -12928 3779 -12894 3803
rect -12928 3769 -12894 3779
rect -12928 3711 -12894 3731
rect -12928 3697 -12894 3711
rect -12928 3643 -12894 3659
rect -12928 3625 -12894 3643
rect -12928 3575 -12894 3587
rect -12928 3553 -12894 3575
rect -12928 3507 -12894 3515
rect -12928 3481 -12894 3507
rect -12832 4425 -12798 4451
rect -12832 4417 -12798 4425
rect -12832 4357 -12798 4379
rect -12832 4345 -12798 4357
rect -12832 4289 -12798 4307
rect -12832 4273 -12798 4289
rect -12832 4221 -12798 4235
rect -12832 4201 -12798 4221
rect -12832 4153 -12798 4163
rect -12832 4129 -12798 4153
rect -12832 4085 -12798 4091
rect -12832 4057 -12798 4085
rect -12832 4017 -12798 4019
rect -12832 3985 -12798 4017
rect -12832 3915 -12798 3947
rect -12832 3913 -12798 3915
rect -12832 3847 -12798 3875
rect -12832 3841 -12798 3847
rect -12832 3779 -12798 3803
rect -12832 3769 -12798 3779
rect -12832 3711 -12798 3731
rect -12832 3697 -12798 3711
rect -12832 3643 -12798 3659
rect -12832 3625 -12798 3643
rect -12832 3575 -12798 3587
rect -12832 3553 -12798 3575
rect -12832 3507 -12798 3515
rect -12832 3481 -12798 3507
rect -21714 3241 -21680 3275
rect -22974 3096 -22940 3130
rect -20050 3247 -20016 3281
rect -20771 3098 -20737 3132
rect -21716 2982 -21682 3016
rect -18846 3253 -18812 3287
rect -19118 3111 -19084 3145
rect -20048 2984 -20014 3018
rect -18158 3235 -18124 3269
rect -18302 3113 -18268 3147
rect -18850 3028 -18816 3062
rect -23492 2813 -23458 2839
rect -23492 2805 -23458 2813
rect -23492 2745 -23458 2767
rect -23492 2733 -23458 2745
rect -23492 2677 -23458 2695
rect -23492 2661 -23458 2677
rect -23492 2609 -23458 2623
rect -23492 2589 -23458 2609
rect -23492 2541 -23458 2551
rect -23492 2517 -23458 2541
rect -23492 2473 -23458 2479
rect -23492 2445 -23458 2473
rect -23492 2405 -23458 2407
rect -23492 2373 -23458 2405
rect -23492 2303 -23458 2335
rect -23492 2301 -23458 2303
rect -23492 2235 -23458 2263
rect -23492 2229 -23458 2235
rect -23492 2167 -23458 2191
rect -23492 2157 -23458 2167
rect -23492 2099 -23458 2119
rect -23492 2085 -23458 2099
rect -23492 2031 -23458 2047
rect -23492 2013 -23458 2031
rect -23492 1963 -23458 1975
rect -23492 1941 -23458 1963
rect -23492 1895 -23458 1903
rect -23492 1869 -23458 1895
rect -23396 2813 -23362 2839
rect -23396 2805 -23362 2813
rect -23396 2745 -23362 2767
rect -23396 2733 -23362 2745
rect -23396 2677 -23362 2695
rect -23396 2661 -23362 2677
rect -23396 2609 -23362 2623
rect -23396 2589 -23362 2609
rect -23396 2541 -23362 2551
rect -23396 2517 -23362 2541
rect -23396 2473 -23362 2479
rect -23396 2445 -23362 2473
rect -23396 2405 -23362 2407
rect -23396 2373 -23362 2405
rect -23396 2303 -23362 2335
rect -23396 2301 -23362 2303
rect -23396 2235 -23362 2263
rect -23396 2229 -23362 2235
rect -23396 2167 -23362 2191
rect -23396 2157 -23362 2167
rect -23396 2099 -23362 2119
rect -23396 2085 -23362 2099
rect -23396 2031 -23362 2047
rect -23396 2013 -23362 2031
rect -23396 1963 -23362 1975
rect -23396 1941 -23362 1963
rect -23396 1895 -23362 1903
rect -23396 1869 -23362 1895
rect -23300 2813 -23266 2839
rect -23300 2805 -23266 2813
rect -23300 2745 -23266 2767
rect -23300 2733 -23266 2745
rect -23300 2677 -23266 2695
rect -23300 2661 -23266 2677
rect -23300 2609 -23266 2623
rect -23300 2589 -23266 2609
rect -23300 2541 -23266 2551
rect -23300 2517 -23266 2541
rect -23300 2473 -23266 2479
rect -23300 2445 -23266 2473
rect -23300 2405 -23266 2407
rect -23300 2373 -23266 2405
rect -23300 2303 -23266 2335
rect -23300 2301 -23266 2303
rect -23300 2235 -23266 2263
rect -23300 2229 -23266 2235
rect -23300 2167 -23266 2191
rect -23300 2157 -23266 2167
rect -23300 2099 -23266 2119
rect -23300 2085 -23266 2099
rect -23300 2031 -23266 2047
rect -23300 2013 -23266 2031
rect -23300 1963 -23266 1975
rect -23300 1941 -23266 1963
rect -23300 1895 -23266 1903
rect -23300 1869 -23266 1895
rect -23204 2813 -23170 2839
rect -23204 2805 -23170 2813
rect -23204 2745 -23170 2767
rect -23204 2733 -23170 2745
rect -23204 2677 -23170 2695
rect -23204 2661 -23170 2677
rect -23204 2609 -23170 2623
rect -23204 2589 -23170 2609
rect -23204 2541 -23170 2551
rect -23204 2517 -23170 2541
rect -23204 2473 -23170 2479
rect -23204 2445 -23170 2473
rect -23204 2405 -23170 2407
rect -23204 2373 -23170 2405
rect -23204 2303 -23170 2335
rect -23204 2301 -23170 2303
rect -23204 2235 -23170 2263
rect -23204 2229 -23170 2235
rect -23204 2167 -23170 2191
rect -23204 2157 -23170 2167
rect -23204 2099 -23170 2119
rect -23204 2085 -23170 2099
rect -23204 2031 -23170 2047
rect -23204 2013 -23170 2031
rect -23204 1963 -23170 1975
rect -23204 1941 -23170 1963
rect -23204 1895 -23170 1903
rect -23204 1869 -23170 1895
rect -23108 2813 -23074 2839
rect -23108 2805 -23074 2813
rect -23108 2745 -23074 2767
rect -23108 2733 -23074 2745
rect -23108 2677 -23074 2695
rect -23108 2661 -23074 2677
rect -23108 2609 -23074 2623
rect -23108 2589 -23074 2609
rect -23108 2541 -23074 2551
rect -23108 2517 -23074 2541
rect -23108 2473 -23074 2479
rect -23108 2445 -23074 2473
rect -23108 2405 -23074 2407
rect -23108 2373 -23074 2405
rect -23108 2303 -23074 2335
rect -23108 2301 -23074 2303
rect -23108 2235 -23074 2263
rect -23108 2229 -23074 2235
rect -23108 2167 -23074 2191
rect -23108 2157 -23074 2167
rect -23108 2099 -23074 2119
rect -23108 2085 -23074 2099
rect -23108 2031 -23074 2047
rect -23108 2013 -23074 2031
rect -23108 1963 -23074 1975
rect -23108 1941 -23074 1963
rect -23108 1895 -23074 1903
rect -23108 1869 -23074 1895
rect -23012 2813 -22978 2839
rect -23012 2805 -22978 2813
rect -23012 2745 -22978 2767
rect -23012 2733 -22978 2745
rect -23012 2677 -22978 2695
rect -23012 2661 -22978 2677
rect -23012 2609 -22978 2623
rect -23012 2589 -22978 2609
rect -23012 2541 -22978 2551
rect -23012 2517 -22978 2541
rect -23012 2473 -22978 2479
rect -23012 2445 -22978 2473
rect -23012 2405 -22978 2407
rect -23012 2373 -22978 2405
rect -23012 2303 -22978 2335
rect -23012 2301 -22978 2303
rect -23012 2235 -22978 2263
rect -23012 2229 -22978 2235
rect -23012 2167 -22978 2191
rect -23012 2157 -22978 2167
rect -23012 2099 -22978 2119
rect -23012 2085 -22978 2099
rect -23012 2031 -22978 2047
rect -23012 2013 -22978 2031
rect -23012 1963 -22978 1975
rect -23012 1941 -22978 1963
rect -23012 1895 -22978 1903
rect -23012 1869 -22978 1895
rect -22916 2813 -22882 2839
rect -22916 2805 -22882 2813
rect -22916 2745 -22882 2767
rect -22916 2733 -22882 2745
rect -22916 2677 -22882 2695
rect -22916 2661 -22882 2677
rect -22916 2609 -22882 2623
rect -22916 2589 -22882 2609
rect -22916 2541 -22882 2551
rect -22916 2517 -22882 2541
rect -22916 2473 -22882 2479
rect -22916 2445 -22882 2473
rect -22916 2405 -22882 2407
rect -22916 2373 -22882 2405
rect -22916 2303 -22882 2335
rect -22916 2301 -22882 2303
rect -22916 2235 -22882 2263
rect -22916 2229 -22882 2235
rect -22916 2167 -22882 2191
rect -22916 2157 -22882 2167
rect -22916 2099 -22882 2119
rect -22916 2085 -22882 2099
rect -22916 2031 -22882 2047
rect -22916 2013 -22882 2031
rect -22916 1963 -22882 1975
rect -22916 1941 -22882 1963
rect -22916 1895 -22882 1903
rect -22916 1869 -22882 1895
rect -22820 2813 -22786 2839
rect -22820 2805 -22786 2813
rect -22820 2745 -22786 2767
rect -22820 2733 -22786 2745
rect -22820 2677 -22786 2695
rect -22820 2661 -22786 2677
rect -22820 2609 -22786 2623
rect -22820 2589 -22786 2609
rect -22820 2541 -22786 2551
rect -22820 2517 -22786 2541
rect -22820 2473 -22786 2479
rect -22820 2445 -22786 2473
rect -22820 2405 -22786 2407
rect -22820 2373 -22786 2405
rect -22820 2303 -22786 2335
rect -22820 2301 -22786 2303
rect -22820 2235 -22786 2263
rect -22820 2229 -22786 2235
rect -22820 2167 -22786 2191
rect -22820 2157 -22786 2167
rect -22820 2099 -22786 2119
rect -22820 2085 -22786 2099
rect -22820 2031 -22786 2047
rect -22820 2013 -22786 2031
rect -22820 1963 -22786 1975
rect -22820 1941 -22786 1963
rect -22820 1895 -22786 1903
rect -22820 1869 -22786 1895
rect -22724 2813 -22690 2839
rect -22724 2805 -22690 2813
rect -22724 2745 -22690 2767
rect -22724 2733 -22690 2745
rect -22724 2677 -22690 2695
rect -22724 2661 -22690 2677
rect -22724 2609 -22690 2623
rect -22724 2589 -22690 2609
rect -22724 2541 -22690 2551
rect -22724 2517 -22690 2541
rect -22724 2473 -22690 2479
rect -22724 2445 -22690 2473
rect -22724 2405 -22690 2407
rect -22724 2373 -22690 2405
rect -22724 2303 -22690 2335
rect -22724 2301 -22690 2303
rect -22724 2235 -22690 2263
rect -22724 2229 -22690 2235
rect -22724 2167 -22690 2191
rect -22724 2157 -22690 2167
rect -22724 2099 -22690 2119
rect -22724 2085 -22690 2099
rect -22724 2031 -22690 2047
rect -22724 2013 -22690 2031
rect -22724 1963 -22690 1975
rect -22724 1941 -22690 1963
rect -22724 1895 -22690 1903
rect -22724 1869 -22690 1895
rect -22628 2813 -22594 2839
rect -22628 2805 -22594 2813
rect -22628 2745 -22594 2767
rect -22628 2733 -22594 2745
rect -22628 2677 -22594 2695
rect -22628 2661 -22594 2677
rect -22628 2609 -22594 2623
rect -22628 2589 -22594 2609
rect -22628 2541 -22594 2551
rect -22628 2517 -22594 2541
rect -22628 2473 -22594 2479
rect -22628 2445 -22594 2473
rect -22628 2405 -22594 2407
rect -22628 2373 -22594 2405
rect -22628 2303 -22594 2335
rect -22628 2301 -22594 2303
rect -22628 2235 -22594 2263
rect -22628 2229 -22594 2235
rect -22628 2167 -22594 2191
rect -22628 2157 -22594 2167
rect -22628 2099 -22594 2119
rect -22628 2085 -22594 2099
rect -22628 2031 -22594 2047
rect -22628 2013 -22594 2031
rect -22628 1963 -22594 1975
rect -22628 1941 -22594 1963
rect -22628 1895 -22594 1903
rect -22628 1869 -22594 1895
rect -22532 2813 -22498 2839
rect -22532 2805 -22498 2813
rect -22532 2745 -22498 2767
rect -22532 2733 -22498 2745
rect -22532 2677 -22498 2695
rect -22532 2661 -22498 2677
rect -22532 2609 -22498 2623
rect -22532 2589 -22498 2609
rect -22532 2541 -22498 2551
rect -22532 2517 -22498 2541
rect -22532 2473 -22498 2479
rect -22532 2445 -22498 2473
rect -22532 2405 -22498 2407
rect -22532 2373 -22498 2405
rect -22532 2303 -22498 2335
rect -22532 2301 -22498 2303
rect -22532 2235 -22498 2263
rect -22532 2229 -22498 2235
rect -22532 2167 -22498 2191
rect -22532 2157 -22498 2167
rect -22532 2099 -22498 2119
rect -22532 2085 -22498 2099
rect -22532 2031 -22498 2047
rect -22532 2013 -22498 2031
rect -22532 1963 -22498 1975
rect -22532 1941 -22498 1963
rect -22532 1895 -22498 1903
rect -22532 1869 -22498 1895
rect -22436 2813 -22402 2839
rect -22436 2805 -22402 2813
rect -22436 2745 -22402 2767
rect -22436 2733 -22402 2745
rect -22436 2677 -22402 2695
rect -22436 2661 -22402 2677
rect -22436 2609 -22402 2623
rect -22436 2589 -22402 2609
rect -22436 2541 -22402 2551
rect -22436 2517 -22402 2541
rect -22436 2473 -22402 2479
rect -22436 2445 -22402 2473
rect -22436 2405 -22402 2407
rect -22436 2373 -22402 2405
rect -22436 2303 -22402 2335
rect -22436 2301 -22402 2303
rect -22436 2235 -22402 2263
rect -22436 2229 -22402 2235
rect -22436 2167 -22402 2191
rect -22436 2157 -22402 2167
rect -22436 2099 -22402 2119
rect -22436 2085 -22402 2099
rect -22436 2031 -22402 2047
rect -22436 2013 -22402 2031
rect -22436 1963 -22402 1975
rect -22436 1941 -22402 1963
rect -22436 1895 -22402 1903
rect -22436 1869 -22402 1895
rect -22340 2813 -22306 2839
rect -22340 2805 -22306 2813
rect -22340 2745 -22306 2767
rect -22340 2733 -22306 2745
rect -22340 2677 -22306 2695
rect -22340 2661 -22306 2677
rect -22340 2609 -22306 2623
rect -22340 2589 -22306 2609
rect -22340 2541 -22306 2551
rect -22340 2517 -22306 2541
rect -22340 2473 -22306 2479
rect -22340 2445 -22306 2473
rect -22340 2405 -22306 2407
rect -22340 2373 -22306 2405
rect -22340 2303 -22306 2335
rect -22340 2301 -22306 2303
rect -22340 2235 -22306 2263
rect -22340 2229 -22306 2235
rect -22340 2167 -22306 2191
rect -22340 2157 -22306 2167
rect -22340 2099 -22306 2119
rect -22340 2085 -22306 2099
rect -22340 2031 -22306 2047
rect -22340 2013 -22306 2031
rect -22340 1963 -22306 1975
rect -22340 1941 -22306 1963
rect -22340 1895 -22306 1903
rect -22340 1869 -22306 1895
rect -22244 2813 -22210 2839
rect -22244 2805 -22210 2813
rect -22244 2745 -22210 2767
rect -22244 2733 -22210 2745
rect -22244 2677 -22210 2695
rect -22244 2661 -22210 2677
rect -22244 2609 -22210 2623
rect -22244 2589 -22210 2609
rect -22244 2541 -22210 2551
rect -22244 2517 -22210 2541
rect -22244 2473 -22210 2479
rect -22244 2445 -22210 2473
rect -22244 2405 -22210 2407
rect -22244 2373 -22210 2405
rect -22244 2303 -22210 2335
rect -22244 2301 -22210 2303
rect -22244 2235 -22210 2263
rect -22244 2229 -22210 2235
rect -22244 2167 -22210 2191
rect -22244 2157 -22210 2167
rect -22244 2099 -22210 2119
rect -22244 2085 -22210 2099
rect -22244 2031 -22210 2047
rect -22244 2013 -22210 2031
rect -22244 1963 -22210 1975
rect -22244 1941 -22210 1963
rect -22244 1895 -22210 1903
rect -22244 1869 -22210 1895
rect -22148 2813 -22114 2839
rect -22148 2805 -22114 2813
rect -22148 2745 -22114 2767
rect -22148 2733 -22114 2745
rect -22148 2677 -22114 2695
rect -22148 2661 -22114 2677
rect -22148 2609 -22114 2623
rect -22148 2589 -22114 2609
rect -22148 2541 -22114 2551
rect -22148 2517 -22114 2541
rect -22148 2473 -22114 2479
rect -22148 2445 -22114 2473
rect -22148 2405 -22114 2407
rect -22148 2373 -22114 2405
rect -22148 2303 -22114 2335
rect -22148 2301 -22114 2303
rect -22148 2235 -22114 2263
rect -22148 2229 -22114 2235
rect -22148 2167 -22114 2191
rect -22148 2157 -22114 2167
rect -22148 2099 -22114 2119
rect -22148 2085 -22114 2099
rect -22148 2031 -22114 2047
rect -22148 2013 -22114 2031
rect -22148 1963 -22114 1975
rect -22148 1941 -22114 1963
rect -22148 1895 -22114 1903
rect -22148 1869 -22114 1895
rect -22052 2813 -22018 2839
rect -22052 2805 -22018 2813
rect -22052 2745 -22018 2767
rect -22052 2733 -22018 2745
rect -22052 2677 -22018 2695
rect -22052 2661 -22018 2677
rect -22052 2609 -22018 2623
rect -22052 2589 -22018 2609
rect -22052 2541 -22018 2551
rect -22052 2517 -22018 2541
rect -22052 2473 -22018 2479
rect -22052 2445 -22018 2473
rect -22052 2405 -22018 2407
rect -22052 2373 -22018 2405
rect -22052 2303 -22018 2335
rect -22052 2301 -22018 2303
rect -22052 2235 -22018 2263
rect -22052 2229 -22018 2235
rect -22052 2167 -22018 2191
rect -22052 2157 -22018 2167
rect -22052 2099 -22018 2119
rect -22052 2085 -22018 2099
rect -22052 2031 -22018 2047
rect -22052 2013 -22018 2031
rect -22052 1963 -22018 1975
rect -22052 1941 -22018 1963
rect -22052 1895 -22018 1903
rect -22052 1869 -22018 1895
rect -21956 2813 -21922 2839
rect -21956 2805 -21922 2813
rect -21956 2745 -21922 2767
rect -21956 2733 -21922 2745
rect -21956 2677 -21922 2695
rect -21956 2661 -21922 2677
rect -21956 2609 -21922 2623
rect -21956 2589 -21922 2609
rect -21956 2541 -21922 2551
rect -21956 2517 -21922 2541
rect -21956 2473 -21922 2479
rect -21956 2445 -21922 2473
rect -21956 2405 -21922 2407
rect -21956 2373 -21922 2405
rect -21956 2303 -21922 2335
rect -21956 2301 -21922 2303
rect -21956 2235 -21922 2263
rect -21956 2229 -21922 2235
rect -21956 2167 -21922 2191
rect -21956 2157 -21922 2167
rect -21956 2099 -21922 2119
rect -21956 2085 -21922 2099
rect -21956 2031 -21922 2047
rect -21956 2013 -21922 2031
rect -21956 1963 -21922 1975
rect -21956 1941 -21922 1963
rect -21956 1895 -21922 1903
rect -21956 1869 -21922 1895
rect -21860 2813 -21826 2839
rect -21860 2805 -21826 2813
rect -21860 2745 -21826 2767
rect -21860 2733 -21826 2745
rect -21860 2677 -21826 2695
rect -21860 2661 -21826 2677
rect -21860 2609 -21826 2623
rect -21860 2589 -21826 2609
rect -21860 2541 -21826 2551
rect -21860 2517 -21826 2541
rect -21860 2473 -21826 2479
rect -21860 2445 -21826 2473
rect -21860 2405 -21826 2407
rect -21860 2373 -21826 2405
rect -21860 2303 -21826 2335
rect -21860 2301 -21826 2303
rect -21860 2235 -21826 2263
rect -21860 2229 -21826 2235
rect -21860 2167 -21826 2191
rect -21860 2157 -21826 2167
rect -21860 2099 -21826 2119
rect -21860 2085 -21826 2099
rect -21860 2031 -21826 2047
rect -21860 2013 -21826 2031
rect -21860 1963 -21826 1975
rect -21860 1941 -21826 1963
rect -21860 1895 -21826 1903
rect -21860 1869 -21826 1895
rect -21764 2813 -21730 2839
rect -21764 2805 -21730 2813
rect -21764 2745 -21730 2767
rect -21764 2733 -21730 2745
rect -21764 2677 -21730 2695
rect -21764 2661 -21730 2677
rect -21764 2609 -21730 2623
rect -21764 2589 -21730 2609
rect -21764 2541 -21730 2551
rect -21764 2517 -21730 2541
rect -21764 2473 -21730 2479
rect -21764 2445 -21730 2473
rect -21764 2405 -21730 2407
rect -21764 2373 -21730 2405
rect -21764 2303 -21730 2335
rect -21764 2301 -21730 2303
rect -21764 2235 -21730 2263
rect -21764 2229 -21730 2235
rect -21764 2167 -21730 2191
rect -21764 2157 -21730 2167
rect -21764 2099 -21730 2119
rect -21764 2085 -21730 2099
rect -21764 2031 -21730 2047
rect -21764 2013 -21730 2031
rect -21764 1963 -21730 1975
rect -21764 1941 -21730 1963
rect -21764 1895 -21730 1903
rect -21764 1869 -21730 1895
rect -21668 2813 -21634 2839
rect -21668 2805 -21634 2813
rect -21668 2745 -21634 2767
rect -21668 2733 -21634 2745
rect -21668 2677 -21634 2695
rect -21668 2661 -21634 2677
rect -21668 2609 -21634 2623
rect -21668 2589 -21634 2609
rect -21668 2541 -21634 2551
rect -21668 2517 -21634 2541
rect -21668 2473 -21634 2479
rect -21668 2445 -21634 2473
rect -21668 2405 -21634 2407
rect -21668 2373 -21634 2405
rect -21668 2303 -21634 2335
rect -21668 2301 -21634 2303
rect -21668 2235 -21634 2263
rect -21668 2229 -21634 2235
rect -21668 2167 -21634 2191
rect -21668 2157 -21634 2167
rect -21668 2099 -21634 2119
rect -21668 2085 -21634 2099
rect -21668 2031 -21634 2047
rect -21668 2013 -21634 2031
rect -21668 1963 -21634 1975
rect -21668 1941 -21634 1963
rect -21668 1895 -21634 1903
rect -21668 1869 -21634 1895
rect -21572 2813 -21538 2839
rect -21572 2805 -21538 2813
rect -21572 2745 -21538 2767
rect -21572 2733 -21538 2745
rect -21572 2677 -21538 2695
rect -21572 2661 -21538 2677
rect -21572 2609 -21538 2623
rect -21572 2589 -21538 2609
rect -21572 2541 -21538 2551
rect -21572 2517 -21538 2541
rect -21572 2473 -21538 2479
rect -21572 2445 -21538 2473
rect -21572 2405 -21538 2407
rect -21572 2373 -21538 2405
rect -21572 2303 -21538 2335
rect -21572 2301 -21538 2303
rect -21572 2235 -21538 2263
rect -21572 2229 -21538 2235
rect -21572 2167 -21538 2191
rect -21572 2157 -21538 2167
rect -21572 2099 -21538 2119
rect -21572 2085 -21538 2099
rect -21572 2031 -21538 2047
rect -21572 2013 -21538 2031
rect -21572 1963 -21538 1975
rect -21572 1941 -21538 1963
rect -21572 1895 -21538 1903
rect -21572 1869 -21538 1895
rect -21344 2805 -21310 2831
rect -21344 2797 -21310 2805
rect -21344 2737 -21310 2759
rect -21344 2725 -21310 2737
rect -21344 2669 -21310 2687
rect -21344 2653 -21310 2669
rect -21344 2601 -21310 2615
rect -21344 2581 -21310 2601
rect -21344 2533 -21310 2543
rect -21344 2509 -21310 2533
rect -21344 2465 -21310 2471
rect -21344 2437 -21310 2465
rect -21344 2397 -21310 2399
rect -21344 2365 -21310 2397
rect -21344 2295 -21310 2327
rect -21344 2293 -21310 2295
rect -21344 2227 -21310 2255
rect -21344 2221 -21310 2227
rect -21344 2159 -21310 2183
rect -21344 2149 -21310 2159
rect -21344 2091 -21310 2111
rect -21344 2077 -21310 2091
rect -21344 2023 -21310 2039
rect -21344 2005 -21310 2023
rect -21344 1955 -21310 1967
rect -21344 1933 -21310 1955
rect -21344 1887 -21310 1895
rect -21344 1861 -21310 1887
rect -21248 2805 -21214 2831
rect -21248 2797 -21214 2805
rect -21248 2737 -21214 2759
rect -21248 2725 -21214 2737
rect -21248 2669 -21214 2687
rect -21248 2653 -21214 2669
rect -21248 2601 -21214 2615
rect -21248 2581 -21214 2601
rect -21248 2533 -21214 2543
rect -21248 2509 -21214 2533
rect -21248 2465 -21214 2471
rect -21248 2437 -21214 2465
rect -21248 2397 -21214 2399
rect -21248 2365 -21214 2397
rect -21248 2295 -21214 2327
rect -21248 2293 -21214 2295
rect -21248 2227 -21214 2255
rect -21248 2221 -21214 2227
rect -21248 2159 -21214 2183
rect -21248 2149 -21214 2159
rect -21248 2091 -21214 2111
rect -21248 2077 -21214 2091
rect -21248 2023 -21214 2039
rect -21248 2005 -21214 2023
rect -21248 1955 -21214 1967
rect -21248 1933 -21214 1955
rect -21248 1887 -21214 1895
rect -21248 1861 -21214 1887
rect -21152 2805 -21118 2831
rect -21152 2797 -21118 2805
rect -21152 2737 -21118 2759
rect -21152 2725 -21118 2737
rect -21152 2669 -21118 2687
rect -21152 2653 -21118 2669
rect -21152 2601 -21118 2615
rect -21152 2581 -21118 2601
rect -21152 2533 -21118 2543
rect -21152 2509 -21118 2533
rect -21152 2465 -21118 2471
rect -21152 2437 -21118 2465
rect -21152 2397 -21118 2399
rect -21152 2365 -21118 2397
rect -21152 2295 -21118 2327
rect -21152 2293 -21118 2295
rect -21152 2227 -21118 2255
rect -21152 2221 -21118 2227
rect -21152 2159 -21118 2183
rect -21152 2149 -21118 2159
rect -21152 2091 -21118 2111
rect -21152 2077 -21118 2091
rect -21152 2023 -21118 2039
rect -21152 2005 -21118 2023
rect -21152 1955 -21118 1967
rect -21152 1933 -21118 1955
rect -21152 1887 -21118 1895
rect -21152 1861 -21118 1887
rect -21056 2805 -21022 2831
rect -21056 2797 -21022 2805
rect -21056 2737 -21022 2759
rect -21056 2725 -21022 2737
rect -21056 2669 -21022 2687
rect -21056 2653 -21022 2669
rect -21056 2601 -21022 2615
rect -21056 2581 -21022 2601
rect -21056 2533 -21022 2543
rect -21056 2509 -21022 2533
rect -21056 2465 -21022 2471
rect -21056 2437 -21022 2465
rect -21056 2397 -21022 2399
rect -21056 2365 -21022 2397
rect -21056 2295 -21022 2327
rect -21056 2293 -21022 2295
rect -21056 2227 -21022 2255
rect -21056 2221 -21022 2227
rect -21056 2159 -21022 2183
rect -21056 2149 -21022 2159
rect -21056 2091 -21022 2111
rect -21056 2077 -21022 2091
rect -21056 2023 -21022 2039
rect -21056 2005 -21022 2023
rect -21056 1955 -21022 1967
rect -21056 1933 -21022 1955
rect -21056 1887 -21022 1895
rect -21056 1861 -21022 1887
rect -20960 2805 -20926 2831
rect -20960 2797 -20926 2805
rect -20960 2737 -20926 2759
rect -20960 2725 -20926 2737
rect -20960 2669 -20926 2687
rect -20960 2653 -20926 2669
rect -20960 2601 -20926 2615
rect -20960 2581 -20926 2601
rect -20960 2533 -20926 2543
rect -20960 2509 -20926 2533
rect -20960 2465 -20926 2471
rect -20960 2437 -20926 2465
rect -20960 2397 -20926 2399
rect -20960 2365 -20926 2397
rect -20960 2295 -20926 2327
rect -20960 2293 -20926 2295
rect -20960 2227 -20926 2255
rect -20960 2221 -20926 2227
rect -20960 2159 -20926 2183
rect -20960 2149 -20926 2159
rect -20960 2091 -20926 2111
rect -20960 2077 -20926 2091
rect -20960 2023 -20926 2039
rect -20960 2005 -20926 2023
rect -20960 1955 -20926 1967
rect -20960 1933 -20926 1955
rect -20960 1887 -20926 1895
rect -20960 1861 -20926 1887
rect -20864 2805 -20830 2831
rect -20864 2797 -20830 2805
rect -20864 2737 -20830 2759
rect -20864 2725 -20830 2737
rect -20864 2669 -20830 2687
rect -20864 2653 -20830 2669
rect -20864 2601 -20830 2615
rect -20864 2581 -20830 2601
rect -20864 2533 -20830 2543
rect -20864 2509 -20830 2533
rect -20864 2465 -20830 2471
rect -20864 2437 -20830 2465
rect -20864 2397 -20830 2399
rect -20864 2365 -20830 2397
rect -20864 2295 -20830 2327
rect -20864 2293 -20830 2295
rect -20864 2227 -20830 2255
rect -20864 2221 -20830 2227
rect -20864 2159 -20830 2183
rect -20864 2149 -20830 2159
rect -20864 2091 -20830 2111
rect -20864 2077 -20830 2091
rect -20864 2023 -20830 2039
rect -20864 2005 -20830 2023
rect -20864 1955 -20830 1967
rect -20864 1933 -20830 1955
rect -20864 1887 -20830 1895
rect -20864 1861 -20830 1887
rect -20768 2805 -20734 2831
rect -20768 2797 -20734 2805
rect -20768 2737 -20734 2759
rect -20768 2725 -20734 2737
rect -20768 2669 -20734 2687
rect -20768 2653 -20734 2669
rect -20768 2601 -20734 2615
rect -20768 2581 -20734 2601
rect -20768 2533 -20734 2543
rect -20768 2509 -20734 2533
rect -20768 2465 -20734 2471
rect -20768 2437 -20734 2465
rect -20768 2397 -20734 2399
rect -20768 2365 -20734 2397
rect -20768 2295 -20734 2327
rect -20768 2293 -20734 2295
rect -20768 2227 -20734 2255
rect -20768 2221 -20734 2227
rect -20768 2159 -20734 2183
rect -20768 2149 -20734 2159
rect -20768 2091 -20734 2111
rect -20768 2077 -20734 2091
rect -20768 2023 -20734 2039
rect -20768 2005 -20734 2023
rect -20768 1955 -20734 1967
rect -20768 1933 -20734 1955
rect -20768 1887 -20734 1895
rect -20768 1861 -20734 1887
rect -20672 2805 -20638 2831
rect -20672 2797 -20638 2805
rect -20672 2737 -20638 2759
rect -20672 2725 -20638 2737
rect -20672 2669 -20638 2687
rect -20672 2653 -20638 2669
rect -20672 2601 -20638 2615
rect -20672 2581 -20638 2601
rect -20672 2533 -20638 2543
rect -20672 2509 -20638 2533
rect -20672 2465 -20638 2471
rect -20672 2437 -20638 2465
rect -20672 2397 -20638 2399
rect -20672 2365 -20638 2397
rect -20672 2295 -20638 2327
rect -20672 2293 -20638 2295
rect -20672 2227 -20638 2255
rect -20672 2221 -20638 2227
rect -20672 2159 -20638 2183
rect -20672 2149 -20638 2159
rect -20672 2091 -20638 2111
rect -20672 2077 -20638 2091
rect -20672 2023 -20638 2039
rect -20672 2005 -20638 2023
rect -20672 1955 -20638 1967
rect -20672 1933 -20638 1955
rect -20672 1887 -20638 1895
rect -20672 1861 -20638 1887
rect -20576 2805 -20542 2831
rect -20576 2797 -20542 2805
rect -20576 2737 -20542 2759
rect -20576 2725 -20542 2737
rect -20576 2669 -20542 2687
rect -20576 2653 -20542 2669
rect -20576 2601 -20542 2615
rect -20576 2581 -20542 2601
rect -20576 2533 -20542 2543
rect -20576 2509 -20542 2533
rect -20576 2465 -20542 2471
rect -20576 2437 -20542 2465
rect -20576 2397 -20542 2399
rect -20576 2365 -20542 2397
rect -20576 2295 -20542 2327
rect -20576 2293 -20542 2295
rect -20576 2227 -20542 2255
rect -20576 2221 -20542 2227
rect -20576 2159 -20542 2183
rect -20576 2149 -20542 2159
rect -20576 2091 -20542 2111
rect -20576 2077 -20542 2091
rect -20576 2023 -20542 2039
rect -20576 2005 -20542 2023
rect -20576 1955 -20542 1967
rect -20576 1933 -20542 1955
rect -20576 1887 -20542 1895
rect -20576 1861 -20542 1887
rect -20480 2805 -20446 2831
rect -20480 2797 -20446 2805
rect -20480 2737 -20446 2759
rect -20480 2725 -20446 2737
rect -20480 2669 -20446 2687
rect -20480 2653 -20446 2669
rect -20480 2601 -20446 2615
rect -20480 2581 -20446 2601
rect -20480 2533 -20446 2543
rect -20480 2509 -20446 2533
rect -20480 2465 -20446 2471
rect -20480 2437 -20446 2465
rect -20480 2397 -20446 2399
rect -20480 2365 -20446 2397
rect -20480 2295 -20446 2327
rect -20480 2293 -20446 2295
rect -20480 2227 -20446 2255
rect -20480 2221 -20446 2227
rect -20480 2159 -20446 2183
rect -20480 2149 -20446 2159
rect -20480 2091 -20446 2111
rect -20480 2077 -20446 2091
rect -20480 2023 -20446 2039
rect -20480 2005 -20446 2023
rect -20480 1955 -20446 1967
rect -20480 1933 -20446 1955
rect -20480 1887 -20446 1895
rect -20480 1861 -20446 1887
rect -20384 2805 -20350 2831
rect -20384 2797 -20350 2805
rect -20384 2737 -20350 2759
rect -20384 2725 -20350 2737
rect -20384 2669 -20350 2687
rect -20384 2653 -20350 2669
rect -20384 2601 -20350 2615
rect -20384 2581 -20350 2601
rect -20384 2533 -20350 2543
rect -20384 2509 -20350 2533
rect -20384 2465 -20350 2471
rect -20384 2437 -20350 2465
rect -20384 2397 -20350 2399
rect -20384 2365 -20350 2397
rect -20384 2295 -20350 2327
rect -20384 2293 -20350 2295
rect -20384 2227 -20350 2255
rect -20384 2221 -20350 2227
rect -20384 2159 -20350 2183
rect -20384 2149 -20350 2159
rect -20384 2091 -20350 2111
rect -20384 2077 -20350 2091
rect -20384 2023 -20350 2039
rect -20384 2005 -20350 2023
rect -20384 1955 -20350 1967
rect -20384 1933 -20350 1955
rect -20384 1887 -20350 1895
rect -20384 1861 -20350 1887
rect -20288 2805 -20254 2831
rect -20288 2797 -20254 2805
rect -20288 2737 -20254 2759
rect -20288 2725 -20254 2737
rect -20288 2669 -20254 2687
rect -20288 2653 -20254 2669
rect -20288 2601 -20254 2615
rect -20288 2581 -20254 2601
rect -20288 2533 -20254 2543
rect -20288 2509 -20254 2533
rect -20288 2465 -20254 2471
rect -20288 2437 -20254 2465
rect -20288 2397 -20254 2399
rect -20288 2365 -20254 2397
rect -20288 2295 -20254 2327
rect -20288 2293 -20254 2295
rect -20288 2227 -20254 2255
rect -20288 2221 -20254 2227
rect -20288 2159 -20254 2183
rect -20288 2149 -20254 2159
rect -20288 2091 -20254 2111
rect -20288 2077 -20254 2091
rect -20288 2023 -20254 2039
rect -20288 2005 -20254 2023
rect -20288 1955 -20254 1967
rect -20288 1933 -20254 1955
rect -20288 1887 -20254 1895
rect -20288 1861 -20254 1887
rect -20192 2805 -20158 2831
rect -20192 2797 -20158 2805
rect -20192 2737 -20158 2759
rect -20192 2725 -20158 2737
rect -20192 2669 -20158 2687
rect -20192 2653 -20158 2669
rect -20192 2601 -20158 2615
rect -20192 2581 -20158 2601
rect -20192 2533 -20158 2543
rect -20192 2509 -20158 2533
rect -20192 2465 -20158 2471
rect -20192 2437 -20158 2465
rect -20192 2397 -20158 2399
rect -20192 2365 -20158 2397
rect -20192 2295 -20158 2327
rect -20192 2293 -20158 2295
rect -20192 2227 -20158 2255
rect -20192 2221 -20158 2227
rect -20192 2159 -20158 2183
rect -20192 2149 -20158 2159
rect -20192 2091 -20158 2111
rect -20192 2077 -20158 2091
rect -20192 2023 -20158 2039
rect -20192 2005 -20158 2023
rect -20192 1955 -20158 1967
rect -20192 1933 -20158 1955
rect -20192 1887 -20158 1895
rect -20192 1861 -20158 1887
rect -20096 2805 -20062 2831
rect -20096 2797 -20062 2805
rect -20096 2737 -20062 2759
rect -20096 2725 -20062 2737
rect -20096 2669 -20062 2687
rect -20096 2653 -20062 2669
rect -20096 2601 -20062 2615
rect -20096 2581 -20062 2601
rect -20096 2533 -20062 2543
rect -20096 2509 -20062 2533
rect -20096 2465 -20062 2471
rect -20096 2437 -20062 2465
rect -20096 2397 -20062 2399
rect -20096 2365 -20062 2397
rect -20096 2295 -20062 2327
rect -20096 2293 -20062 2295
rect -20096 2227 -20062 2255
rect -20096 2221 -20062 2227
rect -20096 2159 -20062 2183
rect -20096 2149 -20062 2159
rect -20096 2091 -20062 2111
rect -20096 2077 -20062 2091
rect -20096 2023 -20062 2039
rect -20096 2005 -20062 2023
rect -20096 1955 -20062 1967
rect -20096 1933 -20062 1955
rect -20096 1887 -20062 1895
rect -20096 1861 -20062 1887
rect -12736 4425 -12702 4451
rect -12736 4417 -12702 4425
rect -12736 4357 -12702 4379
rect -12736 4345 -12702 4357
rect -12736 4289 -12702 4307
rect -12736 4273 -12702 4289
rect -12736 4221 -12702 4235
rect -12736 4201 -12702 4221
rect -12736 4153 -12702 4163
rect -12736 4129 -12702 4153
rect -12736 4085 -12702 4091
rect -12736 4057 -12702 4085
rect -12736 4017 -12702 4019
rect -12736 3985 -12702 4017
rect -12736 3915 -12702 3947
rect -12736 3913 -12702 3915
rect -12736 3847 -12702 3875
rect -12736 3841 -12702 3847
rect -12736 3779 -12702 3803
rect -12736 3769 -12702 3779
rect -12736 3711 -12702 3731
rect -12736 3697 -12702 3711
rect -12736 3643 -12702 3659
rect -12736 3625 -12702 3643
rect -12736 3575 -12702 3587
rect -12736 3553 -12702 3575
rect -12736 3507 -12702 3515
rect -12736 3481 -12702 3507
rect -12640 4425 -12606 4451
rect -12640 4417 -12606 4425
rect -12640 4357 -12606 4379
rect -12640 4345 -12606 4357
rect -12640 4289 -12606 4307
rect -12640 4273 -12606 4289
rect -12640 4221 -12606 4235
rect -12640 4201 -12606 4221
rect -12640 4153 -12606 4163
rect -12640 4129 -12606 4153
rect -12640 4085 -12606 4091
rect -12640 4057 -12606 4085
rect -12640 4017 -12606 4019
rect -12640 3985 -12606 4017
rect -12640 3915 -12606 3947
rect -12640 3913 -12606 3915
rect -12640 3847 -12606 3875
rect -12640 3841 -12606 3847
rect -12640 3779 -12606 3803
rect -12640 3769 -12606 3779
rect -12640 3711 -12606 3731
rect -12640 3697 -12606 3711
rect -12640 3643 -12606 3659
rect -12640 3625 -12606 3643
rect -12640 3575 -12606 3587
rect -12640 3553 -12606 3575
rect -12640 3507 -12606 3515
rect -12640 3481 -12606 3507
rect -12544 4425 -12510 4451
rect -12544 4417 -12510 4425
rect -12544 4357 -12510 4379
rect -12544 4345 -12510 4357
rect -12544 4289 -12510 4307
rect -12544 4273 -12510 4289
rect -12544 4221 -12510 4235
rect -12544 4201 -12510 4221
rect -12544 4153 -12510 4163
rect -12544 4129 -12510 4153
rect -12544 4085 -12510 4091
rect -12544 4057 -12510 4085
rect -12544 4017 -12510 4019
rect -12544 3985 -12510 4017
rect -12544 3915 -12510 3947
rect -12544 3913 -12510 3915
rect -12544 3847 -12510 3875
rect -12544 3841 -12510 3847
rect -12544 3779 -12510 3803
rect -12544 3769 -12510 3779
rect -12544 3711 -12510 3731
rect -12544 3697 -12510 3711
rect -12544 3643 -12510 3659
rect -12544 3625 -12510 3643
rect -12544 3575 -12510 3587
rect -12544 3553 -12510 3575
rect -12544 3507 -12510 3515
rect -12544 3481 -12510 3507
rect -12448 4425 -12414 4451
rect -12448 4417 -12414 4425
rect -12448 4357 -12414 4379
rect -12448 4345 -12414 4357
rect -12448 4289 -12414 4307
rect -12448 4273 -12414 4289
rect -12448 4221 -12414 4235
rect -12448 4201 -12414 4221
rect -12448 4153 -12414 4163
rect -12448 4129 -12414 4153
rect -12448 4085 -12414 4091
rect -12448 4057 -12414 4085
rect -12448 4017 -12414 4019
rect -12448 3985 -12414 4017
rect -12448 3915 -12414 3947
rect -12448 3913 -12414 3915
rect -12448 3847 -12414 3875
rect -12448 3841 -12414 3847
rect -12448 3779 -12414 3803
rect -12448 3769 -12414 3779
rect -12448 3711 -12414 3731
rect -12448 3697 -12414 3711
rect -12448 3643 -12414 3659
rect -12448 3625 -12414 3643
rect -12448 3575 -12414 3587
rect -12448 3553 -12414 3575
rect -12448 3507 -12414 3515
rect -12448 3481 -12414 3507
rect -12352 4425 -12318 4451
rect -12352 4417 -12318 4425
rect -12352 4357 -12318 4379
rect -12352 4345 -12318 4357
rect -12352 4289 -12318 4307
rect -12352 4273 -12318 4289
rect -12352 4221 -12318 4235
rect -12352 4201 -12318 4221
rect -12352 4153 -12318 4163
rect -12352 4129 -12318 4153
rect -12352 4085 -12318 4091
rect -12352 4057 -12318 4085
rect -12352 4017 -12318 4019
rect -12352 3985 -12318 4017
rect -12352 3915 -12318 3947
rect -12352 3913 -12318 3915
rect -12352 3847 -12318 3875
rect -12352 3841 -12318 3847
rect -12352 3779 -12318 3803
rect -12352 3769 -12318 3779
rect -12352 3711 -12318 3731
rect -12352 3697 -12318 3711
rect -12352 3643 -12318 3659
rect -12352 3625 -12318 3643
rect -12352 3575 -12318 3587
rect -12352 3553 -12318 3575
rect -12352 3507 -12318 3515
rect -12352 3481 -12318 3507
rect -12256 4425 -12222 4451
rect -12256 4417 -12222 4425
rect -12256 4357 -12222 4379
rect -12256 4345 -12222 4357
rect -12256 4289 -12222 4307
rect -12256 4273 -12222 4289
rect -12256 4221 -12222 4235
rect -12256 4201 -12222 4221
rect -12256 4153 -12222 4163
rect -12256 4129 -12222 4153
rect -12256 4085 -12222 4091
rect -12256 4057 -12222 4085
rect -12256 4017 -12222 4019
rect -12256 3985 -12222 4017
rect -12256 3915 -12222 3947
rect -12256 3913 -12222 3915
rect -12256 3847 -12222 3875
rect -12256 3841 -12222 3847
rect -12256 3779 -12222 3803
rect -12256 3769 -12222 3779
rect -12256 3711 -12222 3731
rect -12256 3697 -12222 3711
rect -12256 3643 -12222 3659
rect -12256 3625 -12222 3643
rect -12256 3575 -12222 3587
rect -12256 3553 -12222 3575
rect -12256 3507 -12222 3515
rect -12256 3481 -12222 3507
rect -12160 4425 -12126 4451
rect -12160 4417 -12126 4425
rect -12160 4357 -12126 4379
rect -12160 4345 -12126 4357
rect -12160 4289 -12126 4307
rect -12160 4273 -12126 4289
rect -12160 4221 -12126 4235
rect -12160 4201 -12126 4221
rect -12160 4153 -12126 4163
rect -12160 4129 -12126 4153
rect -12160 4085 -12126 4091
rect -12160 4057 -12126 4085
rect -12160 4017 -12126 4019
rect -12160 3985 -12126 4017
rect -12160 3915 -12126 3947
rect -12160 3913 -12126 3915
rect -12160 3847 -12126 3875
rect -12160 3841 -12126 3847
rect -12160 3779 -12126 3803
rect -12160 3769 -12126 3779
rect -12160 3711 -12126 3731
rect -12160 3697 -12126 3711
rect -12160 3643 -12126 3659
rect -12160 3625 -12126 3643
rect -12160 3575 -12126 3587
rect -12160 3553 -12126 3575
rect -12160 3507 -12126 3515
rect -12160 3481 -12126 3507
rect -12064 4425 -12030 4451
rect -12064 4417 -12030 4425
rect -12064 4357 -12030 4379
rect -12064 4345 -12030 4357
rect -12064 4289 -12030 4307
rect -12064 4273 -12030 4289
rect -12064 4221 -12030 4235
rect -12064 4201 -12030 4221
rect -12064 4153 -12030 4163
rect -12064 4129 -12030 4153
rect -12064 4085 -12030 4091
rect -12064 4057 -12030 4085
rect -12064 4017 -12030 4019
rect -12064 3985 -12030 4017
rect -12064 3915 -12030 3947
rect -12064 3913 -12030 3915
rect -12064 3847 -12030 3875
rect -12064 3841 -12030 3847
rect -12064 3779 -12030 3803
rect -12064 3769 -12030 3779
rect -12064 3711 -12030 3731
rect -12064 3697 -12030 3711
rect -12064 3643 -12030 3659
rect -12064 3625 -12030 3643
rect -12064 3575 -12030 3587
rect -12064 3553 -12030 3575
rect -12064 3507 -12030 3515
rect -12064 3481 -12030 3507
rect -11968 4425 -11934 4451
rect -11968 4417 -11934 4425
rect -11968 4357 -11934 4379
rect -11968 4345 -11934 4357
rect -11968 4289 -11934 4307
rect -11968 4273 -11934 4289
rect -11968 4221 -11934 4235
rect -11968 4201 -11934 4221
rect -11968 4153 -11934 4163
rect -11968 4129 -11934 4153
rect -11968 4085 -11934 4091
rect -11968 4057 -11934 4085
rect -11968 4017 -11934 4019
rect -11968 3985 -11934 4017
rect -11968 3915 -11934 3947
rect -11968 3913 -11934 3915
rect -11968 3847 -11934 3875
rect -11968 3841 -11934 3847
rect -11968 3779 -11934 3803
rect -11968 3769 -11934 3779
rect -11968 3711 -11934 3731
rect -11968 3697 -11934 3711
rect -11968 3643 -11934 3659
rect -11968 3625 -11934 3643
rect -11968 3575 -11934 3587
rect -11968 3553 -11934 3575
rect -11968 3507 -11934 3515
rect -11968 3481 -11934 3507
rect -11760 4427 -11726 4453
rect -11760 4419 -11726 4427
rect -11760 4359 -11726 4381
rect -11760 4347 -11726 4359
rect -11760 4291 -11726 4309
rect -11760 4275 -11726 4291
rect -11760 4223 -11726 4237
rect -11760 4203 -11726 4223
rect -11760 4155 -11726 4165
rect -11760 4131 -11726 4155
rect -11760 4087 -11726 4093
rect -11760 4059 -11726 4087
rect -11760 4019 -11726 4021
rect -11760 3987 -11726 4019
rect -11760 3917 -11726 3949
rect -11760 3915 -11726 3917
rect -11760 3849 -11726 3877
rect -11760 3843 -11726 3849
rect -11760 3781 -11726 3805
rect -11760 3771 -11726 3781
rect -11760 3713 -11726 3733
rect -11760 3699 -11726 3713
rect -11760 3645 -11726 3661
rect -11760 3627 -11726 3645
rect -11760 3577 -11726 3589
rect -11760 3555 -11726 3577
rect -11760 3509 -11726 3517
rect -11760 3483 -11726 3509
rect -11664 4427 -11630 4453
rect -11664 4419 -11630 4427
rect -11664 4359 -11630 4381
rect -11664 4347 -11630 4359
rect -11664 4291 -11630 4309
rect -11664 4275 -11630 4291
rect -11664 4223 -11630 4237
rect -11664 4203 -11630 4223
rect -11664 4155 -11630 4165
rect -11664 4131 -11630 4155
rect -11664 4087 -11630 4093
rect -11664 4059 -11630 4087
rect -11664 4019 -11630 4021
rect -11664 3987 -11630 4019
rect -11664 3917 -11630 3949
rect -11664 3915 -11630 3917
rect -11664 3849 -11630 3877
rect -11664 3843 -11630 3849
rect -11664 3781 -11630 3805
rect -11664 3771 -11630 3781
rect -11664 3713 -11630 3733
rect -11664 3699 -11630 3713
rect -11664 3645 -11630 3661
rect -11664 3627 -11630 3645
rect -11664 3577 -11630 3589
rect -11664 3555 -11630 3577
rect -11664 3509 -11630 3517
rect -11664 3483 -11630 3509
rect -11568 4427 -11534 4453
rect -11568 4419 -11534 4427
rect -11568 4359 -11534 4381
rect -11568 4347 -11534 4359
rect -11568 4291 -11534 4309
rect -11568 4275 -11534 4291
rect -11568 4223 -11534 4237
rect -11568 4203 -11534 4223
rect -11568 4155 -11534 4165
rect -11568 4131 -11534 4155
rect -11568 4087 -11534 4093
rect -11568 4059 -11534 4087
rect -11568 4019 -11534 4021
rect -11568 3987 -11534 4019
rect -11568 3917 -11534 3949
rect -11568 3915 -11534 3917
rect -11568 3849 -11534 3877
rect -11568 3843 -11534 3849
rect -11568 3781 -11534 3805
rect -11568 3771 -11534 3781
rect -11568 3713 -11534 3733
rect -11568 3699 -11534 3713
rect -11568 3645 -11534 3661
rect -11568 3627 -11534 3645
rect -11568 3577 -11534 3589
rect -11568 3555 -11534 3577
rect -11568 3509 -11534 3517
rect -11568 3483 -11534 3509
rect -11472 4427 -11438 4453
rect -11472 4419 -11438 4427
rect -11472 4359 -11438 4381
rect -11472 4347 -11438 4359
rect -11472 4291 -11438 4309
rect -11472 4275 -11438 4291
rect -11472 4223 -11438 4237
rect -11472 4203 -11438 4223
rect -11472 4155 -11438 4165
rect -11472 4131 -11438 4155
rect -11472 4087 -11438 4093
rect -11472 4059 -11438 4087
rect -11472 4019 -11438 4021
rect -11472 3987 -11438 4019
rect -11472 3917 -11438 3949
rect -11472 3915 -11438 3917
rect -11472 3849 -11438 3877
rect -11472 3843 -11438 3849
rect -11472 3781 -11438 3805
rect -11472 3771 -11438 3781
rect -11472 3713 -11438 3733
rect -11472 3699 -11438 3713
rect -11472 3645 -11438 3661
rect -11472 3627 -11438 3645
rect -11472 3577 -11438 3589
rect -11472 3555 -11438 3577
rect -11472 3509 -11438 3517
rect -11472 3483 -11438 3509
rect -11376 4427 -11342 4453
rect -11376 4419 -11342 4427
rect -11376 4359 -11342 4381
rect -11376 4347 -11342 4359
rect -11376 4291 -11342 4309
rect -11376 4275 -11342 4291
rect -11376 4223 -11342 4237
rect -11376 4203 -11342 4223
rect -11376 4155 -11342 4165
rect -11376 4131 -11342 4155
rect -11376 4087 -11342 4093
rect -11376 4059 -11342 4087
rect -11376 4019 -11342 4021
rect -11376 3987 -11342 4019
rect -11376 3917 -11342 3949
rect -11376 3915 -11342 3917
rect -11376 3849 -11342 3877
rect -11376 3843 -11342 3849
rect -11376 3781 -11342 3805
rect -11376 3771 -11342 3781
rect -11376 3713 -11342 3733
rect -11376 3699 -11342 3713
rect -11376 3645 -11342 3661
rect -11376 3627 -11342 3645
rect -11376 3577 -11342 3589
rect -11376 3555 -11342 3577
rect -11376 3509 -11342 3517
rect -11376 3483 -11342 3509
rect -11280 4427 -11246 4453
rect -11280 4419 -11246 4427
rect -11280 4359 -11246 4381
rect -11280 4347 -11246 4359
rect -11280 4291 -11246 4309
rect -11280 4275 -11246 4291
rect -11280 4223 -11246 4237
rect -11280 4203 -11246 4223
rect -11280 4155 -11246 4165
rect -11280 4131 -11246 4155
rect -11280 4087 -11246 4093
rect -11280 4059 -11246 4087
rect -11280 4019 -11246 4021
rect -11280 3987 -11246 4019
rect -11280 3917 -11246 3949
rect -11280 3915 -11246 3917
rect -11280 3849 -11246 3877
rect -11280 3843 -11246 3849
rect -11280 3781 -11246 3805
rect -11280 3771 -11246 3781
rect -11280 3713 -11246 3733
rect -11280 3699 -11246 3713
rect -11280 3645 -11246 3661
rect -11280 3627 -11246 3645
rect -11280 3577 -11246 3589
rect -11280 3555 -11246 3577
rect -11280 3509 -11246 3517
rect -11280 3483 -11246 3509
rect -10290 4411 -10256 4437
rect -10290 4403 -10256 4411
rect -10290 4343 -10256 4365
rect -10290 4331 -10256 4343
rect -10290 4275 -10256 4293
rect -10290 4259 -10256 4275
rect -10290 4207 -10256 4221
rect -10290 4187 -10256 4207
rect -10290 4139 -10256 4149
rect -10290 4115 -10256 4139
rect -10290 4071 -10256 4077
rect -10290 4043 -10256 4071
rect -10290 4003 -10256 4005
rect -10290 3971 -10256 4003
rect -10290 3901 -10256 3933
rect -10290 3899 -10256 3901
rect -10290 3833 -10256 3861
rect -10290 3827 -10256 3833
rect -10290 3765 -10256 3789
rect -10290 3755 -10256 3765
rect -10290 3697 -10256 3717
rect -10290 3683 -10256 3697
rect -10290 3629 -10256 3645
rect -10290 3611 -10256 3629
rect -10290 3561 -10256 3573
rect -10290 3539 -10256 3561
rect -10290 3493 -10256 3501
rect -10290 3467 -10256 3493
rect -10194 4411 -10160 4437
rect -10194 4403 -10160 4411
rect -10194 4343 -10160 4365
rect -10194 4331 -10160 4343
rect -10194 4275 -10160 4293
rect -10194 4259 -10160 4275
rect -10194 4207 -10160 4221
rect -10194 4187 -10160 4207
rect -10194 4139 -10160 4149
rect -10194 4115 -10160 4139
rect -10194 4071 -10160 4077
rect -10194 4043 -10160 4071
rect -10194 4003 -10160 4005
rect -10194 3971 -10160 4003
rect -10194 3901 -10160 3933
rect -10194 3899 -10160 3901
rect -10194 3833 -10160 3861
rect -10194 3827 -10160 3833
rect -10194 3765 -10160 3789
rect -10194 3755 -10160 3765
rect -10194 3697 -10160 3717
rect -10194 3683 -10160 3697
rect -10194 3629 -10160 3645
rect -10194 3611 -10160 3629
rect -10194 3561 -10160 3573
rect -10194 3539 -10160 3561
rect -10194 3493 -10160 3501
rect -10194 3467 -10160 3493
rect -10098 4411 -10064 4437
rect -10098 4403 -10064 4411
rect -10098 4343 -10064 4365
rect -10098 4331 -10064 4343
rect -10098 4275 -10064 4293
rect -10098 4259 -10064 4275
rect -10098 4207 -10064 4221
rect -10098 4187 -10064 4207
rect -10098 4139 -10064 4149
rect -10098 4115 -10064 4139
rect -10098 4071 -10064 4077
rect -10098 4043 -10064 4071
rect -10098 4003 -10064 4005
rect -10098 3971 -10064 4003
rect -10098 3901 -10064 3933
rect -10098 3899 -10064 3901
rect -10098 3833 -10064 3861
rect -10098 3827 -10064 3833
rect -10098 3765 -10064 3789
rect -10098 3755 -10064 3765
rect -10098 3697 -10064 3717
rect -10098 3683 -10064 3697
rect -10098 3629 -10064 3645
rect -10098 3611 -10064 3629
rect -10098 3561 -10064 3573
rect -10098 3539 -10064 3561
rect -10098 3493 -10064 3501
rect -10098 3467 -10064 3493
rect -10002 4411 -9968 4437
rect -10002 4403 -9968 4411
rect -10002 4343 -9968 4365
rect -10002 4331 -9968 4343
rect -10002 4275 -9968 4293
rect -10002 4259 -9968 4275
rect -10002 4207 -9968 4221
rect -10002 4187 -9968 4207
rect -10002 4139 -9968 4149
rect -10002 4115 -9968 4139
rect -10002 4071 -9968 4077
rect -10002 4043 -9968 4071
rect -10002 4003 -9968 4005
rect -10002 3971 -9968 4003
rect -10002 3901 -9968 3933
rect -10002 3899 -9968 3901
rect -10002 3833 -9968 3861
rect -10002 3827 -9968 3833
rect -10002 3765 -9968 3789
rect -10002 3755 -9968 3765
rect -10002 3697 -9968 3717
rect -10002 3683 -9968 3697
rect -10002 3629 -9968 3645
rect -10002 3611 -9968 3629
rect -10002 3561 -9968 3573
rect -10002 3539 -9968 3561
rect -10002 3493 -9968 3501
rect -10002 3467 -9968 3493
rect -9906 4411 -9872 4437
rect -9906 4403 -9872 4411
rect -9906 4343 -9872 4365
rect -9906 4331 -9872 4343
rect -9906 4275 -9872 4293
rect -9906 4259 -9872 4275
rect -9906 4207 -9872 4221
rect -9906 4187 -9872 4207
rect -9906 4139 -9872 4149
rect -9906 4115 -9872 4139
rect -9906 4071 -9872 4077
rect -9906 4043 -9872 4071
rect -9906 4003 -9872 4005
rect -9906 3971 -9872 4003
rect -9906 3901 -9872 3933
rect -9906 3899 -9872 3901
rect -9906 3833 -9872 3861
rect -9906 3827 -9872 3833
rect -9906 3765 -9872 3789
rect -9906 3755 -9872 3765
rect -9906 3697 -9872 3717
rect -9906 3683 -9872 3697
rect -9906 3629 -9872 3645
rect -9906 3611 -9872 3629
rect -9906 3561 -9872 3573
rect -9906 3539 -9872 3561
rect -9906 3493 -9872 3501
rect -9906 3467 -9872 3493
rect -9810 4411 -9776 4437
rect -9810 4403 -9776 4411
rect -9810 4343 -9776 4365
rect -9810 4331 -9776 4343
rect -9810 4275 -9776 4293
rect -9810 4259 -9776 4275
rect -9810 4207 -9776 4221
rect -9810 4187 -9776 4207
rect -9810 4139 -9776 4149
rect -9810 4115 -9776 4139
rect -9810 4071 -9776 4077
rect -9810 4043 -9776 4071
rect -9810 4003 -9776 4005
rect -9810 3971 -9776 4003
rect -9810 3901 -9776 3933
rect -9810 3899 -9776 3901
rect -9810 3833 -9776 3861
rect -9810 3827 -9776 3833
rect -9810 3765 -9776 3789
rect -9810 3755 -9776 3765
rect -9810 3697 -9776 3717
rect -9810 3683 -9776 3697
rect -9810 3629 -9776 3645
rect -9810 3611 -9776 3629
rect -9810 3561 -9776 3573
rect -9810 3539 -9776 3561
rect -9810 3493 -9776 3501
rect -9810 3467 -9776 3493
rect -9714 4411 -9680 4437
rect -9714 4403 -9680 4411
rect -9714 4343 -9680 4365
rect -9714 4331 -9680 4343
rect -9714 4275 -9680 4293
rect -9714 4259 -9680 4275
rect -9714 4207 -9680 4221
rect -9714 4187 -9680 4207
rect -9714 4139 -9680 4149
rect -9714 4115 -9680 4139
rect -9714 4071 -9680 4077
rect -9714 4043 -9680 4071
rect -9714 4003 -9680 4005
rect -9714 3971 -9680 4003
rect -9714 3901 -9680 3933
rect -9714 3899 -9680 3901
rect -9714 3833 -9680 3861
rect -9714 3827 -9680 3833
rect -9714 3765 -9680 3789
rect -9714 3755 -9680 3765
rect -9714 3697 -9680 3717
rect -9714 3683 -9680 3697
rect -9714 3629 -9680 3645
rect -9714 3611 -9680 3629
rect -9714 3561 -9680 3573
rect -9714 3539 -9680 3561
rect -9714 3493 -9680 3501
rect -9714 3467 -9680 3493
rect -9618 4411 -9584 4437
rect -9618 4403 -9584 4411
rect -9618 4343 -9584 4365
rect -9618 4331 -9584 4343
rect -9618 4275 -9584 4293
rect -9618 4259 -9584 4275
rect -9618 4207 -9584 4221
rect -9618 4187 -9584 4207
rect -9618 4139 -9584 4149
rect -9618 4115 -9584 4139
rect -9618 4071 -9584 4077
rect -9618 4043 -9584 4071
rect -9618 4003 -9584 4005
rect -9618 3971 -9584 4003
rect -9618 3901 -9584 3933
rect -9618 3899 -9584 3901
rect -9618 3833 -9584 3861
rect -9618 3827 -9584 3833
rect -9618 3765 -9584 3789
rect -9618 3755 -9584 3765
rect -9618 3697 -9584 3717
rect -9618 3683 -9584 3697
rect -9618 3629 -9584 3645
rect -9618 3611 -9584 3629
rect -9618 3561 -9584 3573
rect -9618 3539 -9584 3561
rect -9618 3493 -9584 3501
rect -9618 3467 -9584 3493
rect -9522 4411 -9488 4437
rect -9522 4403 -9488 4411
rect -9522 4343 -9488 4365
rect -9522 4331 -9488 4343
rect -9522 4275 -9488 4293
rect -9522 4259 -9488 4275
rect -9522 4207 -9488 4221
rect -9522 4187 -9488 4207
rect -9522 4139 -9488 4149
rect -9522 4115 -9488 4139
rect -9522 4071 -9488 4077
rect -9522 4043 -9488 4071
rect -9522 4003 -9488 4005
rect -9522 3971 -9488 4003
rect -9522 3901 -9488 3933
rect -9522 3899 -9488 3901
rect -9522 3833 -9488 3861
rect -9522 3827 -9488 3833
rect -9522 3765 -9488 3789
rect -9522 3755 -9488 3765
rect -9522 3697 -9488 3717
rect -9522 3683 -9488 3697
rect -9522 3629 -9488 3645
rect -9522 3611 -9488 3629
rect -9522 3561 -9488 3573
rect -9522 3539 -9488 3561
rect -9522 3493 -9488 3501
rect -9522 3467 -9488 3493
rect -9426 4411 -9392 4437
rect -9426 4403 -9392 4411
rect -9426 4343 -9392 4365
rect -9426 4331 -9392 4343
rect -9426 4275 -9392 4293
rect -9426 4259 -9392 4275
rect -9426 4207 -9392 4221
rect -9426 4187 -9392 4207
rect -9426 4139 -9392 4149
rect -9426 4115 -9392 4139
rect -9426 4071 -9392 4077
rect -9426 4043 -9392 4071
rect -9426 4003 -9392 4005
rect -9426 3971 -9392 4003
rect -9426 3901 -9392 3933
rect -9426 3899 -9392 3901
rect -9426 3833 -9392 3861
rect -9426 3827 -9392 3833
rect -9426 3765 -9392 3789
rect -9426 3755 -9392 3765
rect -9426 3697 -9392 3717
rect -9426 3683 -9392 3697
rect -9426 3629 -9392 3645
rect -9426 3611 -9392 3629
rect -9426 3561 -9392 3573
rect -9426 3539 -9392 3561
rect -9426 3493 -9392 3501
rect -9426 3467 -9392 3493
rect -9330 4411 -9296 4437
rect -9330 4403 -9296 4411
rect -9330 4343 -9296 4365
rect -9330 4331 -9296 4343
rect -9330 4275 -9296 4293
rect -9330 4259 -9296 4275
rect -9330 4207 -9296 4221
rect -9330 4187 -9296 4207
rect -9330 4139 -9296 4149
rect -9330 4115 -9296 4139
rect -9330 4071 -9296 4077
rect -9330 4043 -9296 4071
rect -9330 4003 -9296 4005
rect -9330 3971 -9296 4003
rect -9330 3901 -9296 3933
rect -9330 3899 -9296 3901
rect -9330 3833 -9296 3861
rect -9330 3827 -9296 3833
rect -9330 3765 -9296 3789
rect -9330 3755 -9296 3765
rect -9330 3697 -9296 3717
rect -9330 3683 -9296 3697
rect -9330 3629 -9296 3645
rect -9330 3611 -9296 3629
rect -9330 3561 -9296 3573
rect -9330 3539 -9296 3561
rect -9330 3493 -9296 3501
rect -9330 3467 -9296 3493
rect -9234 4411 -9200 4437
rect -9234 4403 -9200 4411
rect -9234 4343 -9200 4365
rect -9234 4331 -9200 4343
rect -9234 4275 -9200 4293
rect -9234 4259 -9200 4275
rect -9234 4207 -9200 4221
rect -9234 4187 -9200 4207
rect -9234 4139 -9200 4149
rect -9234 4115 -9200 4139
rect -9234 4071 -9200 4077
rect -9234 4043 -9200 4071
rect -9234 4003 -9200 4005
rect -9234 3971 -9200 4003
rect -9234 3901 -9200 3933
rect -9234 3899 -9200 3901
rect -9234 3833 -9200 3861
rect -9234 3827 -9200 3833
rect -9234 3765 -9200 3789
rect -9234 3755 -9200 3765
rect -9234 3697 -9200 3717
rect -9234 3683 -9200 3697
rect -9234 3629 -9200 3645
rect -9234 3611 -9200 3629
rect -9234 3561 -9200 3573
rect -9234 3539 -9200 3561
rect -9234 3493 -9200 3501
rect -9234 3467 -9200 3493
rect -9138 4411 -9104 4437
rect -9138 4403 -9104 4411
rect -9138 4343 -9104 4365
rect -9138 4331 -9104 4343
rect -9138 4275 -9104 4293
rect -9138 4259 -9104 4275
rect -9138 4207 -9104 4221
rect -9138 4187 -9104 4207
rect -9138 4139 -9104 4149
rect -9138 4115 -9104 4139
rect -9138 4071 -9104 4077
rect -9138 4043 -9104 4071
rect -9138 4003 -9104 4005
rect -9138 3971 -9104 4003
rect -9138 3901 -9104 3933
rect -9138 3899 -9104 3901
rect -9138 3833 -9104 3861
rect -9138 3827 -9104 3833
rect -9138 3765 -9104 3789
rect -9138 3755 -9104 3765
rect -9138 3697 -9104 3717
rect -9138 3683 -9104 3697
rect -9138 3629 -9104 3645
rect -9138 3611 -9104 3629
rect -9138 3561 -9104 3573
rect -9138 3539 -9104 3561
rect -9138 3493 -9104 3501
rect -9138 3467 -9104 3493
rect -9042 4411 -9008 4437
rect -9042 4403 -9008 4411
rect -9042 4343 -9008 4365
rect -9042 4331 -9008 4343
rect -9042 4275 -9008 4293
rect -9042 4259 -9008 4275
rect -9042 4207 -9008 4221
rect -9042 4187 -9008 4207
rect -9042 4139 -9008 4149
rect -9042 4115 -9008 4139
rect -9042 4071 -9008 4077
rect -9042 4043 -9008 4071
rect -9042 4003 -9008 4005
rect -9042 3971 -9008 4003
rect -9042 3901 -9008 3933
rect -9042 3899 -9008 3901
rect -9042 3833 -9008 3861
rect -9042 3827 -9008 3833
rect -9042 3765 -9008 3789
rect -9042 3755 -9008 3765
rect -9042 3697 -9008 3717
rect -9042 3683 -9008 3697
rect -9042 3629 -9008 3645
rect -9042 3611 -9008 3629
rect -9042 3561 -9008 3573
rect -9042 3539 -9008 3561
rect -9042 3493 -9008 3501
rect -9042 3467 -9008 3493
rect -8946 4411 -8912 4437
rect -8946 4403 -8912 4411
rect -8946 4343 -8912 4365
rect -8946 4331 -8912 4343
rect -8946 4275 -8912 4293
rect -8946 4259 -8912 4275
rect -8946 4207 -8912 4221
rect -8946 4187 -8912 4207
rect -8946 4139 -8912 4149
rect -8946 4115 -8912 4139
rect -8946 4071 -8912 4077
rect -8946 4043 -8912 4071
rect -8946 4003 -8912 4005
rect -8946 3971 -8912 4003
rect -8946 3901 -8912 3933
rect -8946 3899 -8912 3901
rect -8946 3833 -8912 3861
rect -8946 3827 -8912 3833
rect -8946 3765 -8912 3789
rect -8946 3755 -8912 3765
rect -8946 3697 -8912 3717
rect -8946 3683 -8912 3697
rect -8946 3629 -8912 3645
rect -8946 3611 -8912 3629
rect -8946 3561 -8912 3573
rect -8946 3539 -8912 3561
rect -8946 3493 -8912 3501
rect -8946 3467 -8912 3493
rect -8850 4411 -8816 4437
rect -8850 4403 -8816 4411
rect -8850 4343 -8816 4365
rect -8850 4331 -8816 4343
rect -8850 4275 -8816 4293
rect -8850 4259 -8816 4275
rect -8850 4207 -8816 4221
rect -8850 4187 -8816 4207
rect -8850 4139 -8816 4149
rect -8850 4115 -8816 4139
rect -8850 4071 -8816 4077
rect -8850 4043 -8816 4071
rect -8850 4003 -8816 4005
rect -8850 3971 -8816 4003
rect -8850 3901 -8816 3933
rect -8850 3899 -8816 3901
rect -8850 3833 -8816 3861
rect -8850 3827 -8816 3833
rect -8850 3765 -8816 3789
rect -8850 3755 -8816 3765
rect -8850 3697 -8816 3717
rect -8850 3683 -8816 3697
rect -8850 3629 -8816 3645
rect -8850 3611 -8816 3629
rect -8850 3561 -8816 3573
rect -8850 3539 -8816 3561
rect -8850 3493 -8816 3501
rect -8850 3467 -8816 3493
rect -8754 4411 -8720 4437
rect -8754 4403 -8720 4411
rect -8754 4343 -8720 4365
rect -8754 4331 -8720 4343
rect -8754 4275 -8720 4293
rect -8754 4259 -8720 4275
rect -8754 4207 -8720 4221
rect -8754 4187 -8720 4207
rect -8754 4139 -8720 4149
rect -8754 4115 -8720 4139
rect -8754 4071 -8720 4077
rect -8754 4043 -8720 4071
rect -8754 4003 -8720 4005
rect -8754 3971 -8720 4003
rect -8754 3901 -8720 3933
rect -8754 3899 -8720 3901
rect -8754 3833 -8720 3861
rect -8754 3827 -8720 3833
rect -8754 3765 -8720 3789
rect -8754 3755 -8720 3765
rect -8754 3697 -8720 3717
rect -8754 3683 -8720 3697
rect -8754 3629 -8720 3645
rect -8754 3611 -8720 3629
rect -8754 3561 -8720 3573
rect -8754 3539 -8720 3561
rect -8754 3493 -8720 3501
rect -8754 3467 -8720 3493
rect -8658 4411 -8624 4437
rect -8658 4403 -8624 4411
rect -8658 4343 -8624 4365
rect -8658 4331 -8624 4343
rect -8658 4275 -8624 4293
rect -8658 4259 -8624 4275
rect -8658 4207 -8624 4221
rect -8658 4187 -8624 4207
rect -8658 4139 -8624 4149
rect -8658 4115 -8624 4139
rect -8658 4071 -8624 4077
rect -8658 4043 -8624 4071
rect -8658 4003 -8624 4005
rect -8658 3971 -8624 4003
rect -8658 3901 -8624 3933
rect -8658 3899 -8624 3901
rect -8658 3833 -8624 3861
rect -8658 3827 -8624 3833
rect -8658 3765 -8624 3789
rect -8658 3755 -8624 3765
rect -8658 3697 -8624 3717
rect -8658 3683 -8624 3697
rect -8658 3629 -8624 3645
rect -8658 3611 -8624 3629
rect -8658 3561 -8624 3573
rect -8658 3539 -8624 3561
rect -8658 3493 -8624 3501
rect -8658 3467 -8624 3493
rect -8562 4411 -8528 4437
rect -8562 4403 -8528 4411
rect -8562 4343 -8528 4365
rect -8562 4331 -8528 4343
rect -8562 4275 -8528 4293
rect -8562 4259 -8528 4275
rect -8562 4207 -8528 4221
rect -8562 4187 -8528 4207
rect -8562 4139 -8528 4149
rect -8562 4115 -8528 4139
rect -8562 4071 -8528 4077
rect -8562 4043 -8528 4071
rect -8562 4003 -8528 4005
rect -8562 3971 -8528 4003
rect -8562 3901 -8528 3933
rect -8562 3899 -8528 3901
rect -8562 3833 -8528 3861
rect -8562 3827 -8528 3833
rect -8562 3765 -8528 3789
rect -8562 3755 -8528 3765
rect -8562 3697 -8528 3717
rect -8562 3683 -8528 3697
rect -8562 3629 -8528 3645
rect -8562 3611 -8528 3629
rect -8562 3561 -8528 3573
rect -8562 3539 -8528 3561
rect -8562 3493 -8528 3501
rect -8562 3467 -8528 3493
rect -8466 4411 -8432 4437
rect -8466 4403 -8432 4411
rect -8466 4343 -8432 4365
rect -8466 4331 -8432 4343
rect -8466 4275 -8432 4293
rect -8466 4259 -8432 4275
rect -8466 4207 -8432 4221
rect -8466 4187 -8432 4207
rect -8466 4139 -8432 4149
rect -8466 4115 -8432 4139
rect -8466 4071 -8432 4077
rect -8466 4043 -8432 4071
rect -8466 4003 -8432 4005
rect -8466 3971 -8432 4003
rect -8466 3901 -8432 3933
rect -8466 3899 -8432 3901
rect -8466 3833 -8432 3861
rect -8466 3827 -8432 3833
rect -8466 3765 -8432 3789
rect -8466 3755 -8432 3765
rect -8466 3697 -8432 3717
rect -8466 3683 -8432 3697
rect -8466 3629 -8432 3645
rect -8466 3611 -8432 3629
rect -8466 3561 -8432 3573
rect -8466 3539 -8432 3561
rect -8466 3493 -8432 3501
rect -8466 3467 -8432 3493
rect -8370 4411 -8336 4437
rect -8370 4403 -8336 4411
rect -8370 4343 -8336 4365
rect -8370 4331 -8336 4343
rect -8370 4275 -8336 4293
rect -8370 4259 -8336 4275
rect -8370 4207 -8336 4221
rect -8370 4187 -8336 4207
rect -8370 4139 -8336 4149
rect -8370 4115 -8336 4139
rect -8370 4071 -8336 4077
rect -8370 4043 -8336 4071
rect -8370 4003 -8336 4005
rect -8370 3971 -8336 4003
rect -8370 3901 -8336 3933
rect -8370 3899 -8336 3901
rect -8370 3833 -8336 3861
rect -8370 3827 -8336 3833
rect -8370 3765 -8336 3789
rect -8370 3755 -8336 3765
rect -8370 3697 -8336 3717
rect -8370 3683 -8336 3697
rect -8370 3629 -8336 3645
rect -8370 3611 -8336 3629
rect -8370 3561 -8336 3573
rect -8370 3539 -8336 3561
rect -8370 3493 -8336 3501
rect -8370 3467 -8336 3493
rect -8146 4417 -8112 4443
rect -8146 4409 -8112 4417
rect -8146 4349 -8112 4371
rect -8146 4337 -8112 4349
rect -8146 4281 -8112 4299
rect -8146 4265 -8112 4281
rect -8146 4213 -8112 4227
rect -8146 4193 -8112 4213
rect -8146 4145 -8112 4155
rect -8146 4121 -8112 4145
rect -8146 4077 -8112 4083
rect -8146 4049 -8112 4077
rect -8146 4009 -8112 4011
rect -8146 3977 -8112 4009
rect -8146 3907 -8112 3939
rect -8146 3905 -8112 3907
rect -8146 3839 -8112 3867
rect -8146 3833 -8112 3839
rect -8146 3771 -8112 3795
rect -8146 3761 -8112 3771
rect -8146 3703 -8112 3723
rect -8146 3689 -8112 3703
rect -8146 3635 -8112 3651
rect -8146 3617 -8112 3635
rect -8146 3567 -8112 3579
rect -8146 3545 -8112 3567
rect -8146 3499 -8112 3507
rect -8146 3473 -8112 3499
rect -14884 3253 -14850 3287
rect -16144 3108 -16110 3142
rect -18158 2998 -18124 3032
rect -13220 3259 -13186 3293
rect -13941 3110 -13907 3144
rect -14886 2994 -14852 3028
rect -12016 3265 -11982 3299
rect -12288 3123 -12254 3157
rect -13218 2996 -13184 3030
rect -8050 4417 -8016 4443
rect -8050 4409 -8016 4417
rect -8050 4349 -8016 4371
rect -8050 4337 -8016 4349
rect -8050 4281 -8016 4299
rect -8050 4265 -8016 4281
rect -8050 4213 -8016 4227
rect -8050 4193 -8016 4213
rect -8050 4145 -8016 4155
rect -8050 4121 -8016 4145
rect -8050 4077 -8016 4083
rect -8050 4049 -8016 4077
rect -8050 4009 -8016 4011
rect -8050 3977 -8016 4009
rect -8050 3907 -8016 3939
rect -8050 3905 -8016 3907
rect -8050 3839 -8016 3867
rect -8050 3833 -8016 3839
rect -8050 3771 -8016 3795
rect -8050 3761 -8016 3771
rect -8050 3703 -8016 3723
rect -8050 3689 -8016 3703
rect -8050 3635 -8016 3651
rect -8050 3617 -8016 3635
rect -8050 3567 -8016 3579
rect -8050 3545 -8016 3567
rect -8050 3499 -8016 3507
rect -8050 3473 -8016 3499
rect -7954 4417 -7920 4443
rect -7954 4409 -7920 4417
rect -7954 4349 -7920 4371
rect -7954 4337 -7920 4349
rect -7954 4281 -7920 4299
rect -7954 4265 -7920 4281
rect -7954 4213 -7920 4227
rect -7954 4193 -7920 4213
rect -7954 4145 -7920 4155
rect -7954 4121 -7920 4145
rect -7954 4077 -7920 4083
rect -7954 4049 -7920 4077
rect -7954 4009 -7920 4011
rect -7954 3977 -7920 4009
rect -7954 3907 -7920 3939
rect -7954 3905 -7920 3907
rect -7954 3839 -7920 3867
rect -7954 3833 -7920 3839
rect -7954 3771 -7920 3795
rect -7954 3761 -7920 3771
rect -7954 3703 -7920 3723
rect -7954 3689 -7920 3703
rect -7954 3635 -7920 3651
rect -7954 3617 -7920 3635
rect -7954 3567 -7920 3579
rect -7954 3545 -7920 3567
rect -7954 3499 -7920 3507
rect -7954 3473 -7920 3499
rect -7858 4417 -7824 4443
rect -7858 4409 -7824 4417
rect -7858 4349 -7824 4371
rect -7858 4337 -7824 4349
rect -7858 4281 -7824 4299
rect -7858 4265 -7824 4281
rect -7858 4213 -7824 4227
rect -7858 4193 -7824 4213
rect -7858 4145 -7824 4155
rect -7858 4121 -7824 4145
rect -7858 4077 -7824 4083
rect -7858 4049 -7824 4077
rect -7858 4009 -7824 4011
rect -7858 3977 -7824 4009
rect -7858 3907 -7824 3939
rect -7858 3905 -7824 3907
rect -7858 3839 -7824 3867
rect -7858 3833 -7824 3839
rect -7858 3771 -7824 3795
rect -7858 3761 -7824 3771
rect -7858 3703 -7824 3723
rect -7858 3689 -7824 3703
rect -7858 3635 -7824 3651
rect -7858 3617 -7824 3635
rect -7858 3567 -7824 3579
rect -7858 3545 -7824 3567
rect -7858 3499 -7824 3507
rect -7858 3473 -7824 3499
rect -7762 4417 -7728 4443
rect -7762 4409 -7728 4417
rect -7762 4349 -7728 4371
rect -7762 4337 -7728 4349
rect -7762 4281 -7728 4299
rect -7762 4265 -7728 4281
rect -7762 4213 -7728 4227
rect -7762 4193 -7728 4213
rect -7762 4145 -7728 4155
rect -7762 4121 -7728 4145
rect -7762 4077 -7728 4083
rect -7762 4049 -7728 4077
rect -7762 4009 -7728 4011
rect -7762 3977 -7728 4009
rect -7762 3907 -7728 3939
rect -7762 3905 -7728 3907
rect -7762 3839 -7728 3867
rect -7762 3833 -7728 3839
rect -7762 3771 -7728 3795
rect -7762 3761 -7728 3771
rect -7762 3703 -7728 3723
rect -7762 3689 -7728 3703
rect -7762 3635 -7728 3651
rect -7762 3617 -7728 3635
rect -7762 3567 -7728 3579
rect -7762 3545 -7728 3567
rect -7762 3499 -7728 3507
rect -7762 3473 -7728 3499
rect -7666 4417 -7632 4443
rect -7666 4409 -7632 4417
rect -7666 4349 -7632 4371
rect -7666 4337 -7632 4349
rect -7666 4281 -7632 4299
rect -7666 4265 -7632 4281
rect -7666 4213 -7632 4227
rect -7666 4193 -7632 4213
rect -7666 4145 -7632 4155
rect -7666 4121 -7632 4145
rect -7666 4077 -7632 4083
rect -7666 4049 -7632 4077
rect -7666 4009 -7632 4011
rect -7666 3977 -7632 4009
rect -7666 3907 -7632 3939
rect -7666 3905 -7632 3907
rect -7666 3839 -7632 3867
rect -7666 3833 -7632 3839
rect -7666 3771 -7632 3795
rect -7666 3761 -7632 3771
rect -7666 3703 -7632 3723
rect -7666 3689 -7632 3703
rect -7666 3635 -7632 3651
rect -7666 3617 -7632 3635
rect -7666 3567 -7632 3579
rect -7666 3545 -7632 3567
rect -7666 3499 -7632 3507
rect -7666 3473 -7632 3499
rect -7570 4417 -7536 4443
rect -7570 4409 -7536 4417
rect -7570 4349 -7536 4371
rect -7570 4337 -7536 4349
rect -7570 4281 -7536 4299
rect -7570 4265 -7536 4281
rect -7570 4213 -7536 4227
rect -7570 4193 -7536 4213
rect -7570 4145 -7536 4155
rect -7570 4121 -7536 4145
rect -7570 4077 -7536 4083
rect -7570 4049 -7536 4077
rect -7570 4009 -7536 4011
rect -7570 3977 -7536 4009
rect -7570 3907 -7536 3939
rect -7570 3905 -7536 3907
rect -7570 3839 -7536 3867
rect -7570 3833 -7536 3839
rect -7570 3771 -7536 3795
rect -7570 3761 -7536 3771
rect -7570 3703 -7536 3723
rect -7570 3689 -7536 3703
rect -7570 3635 -7536 3651
rect -7570 3617 -7536 3635
rect -7570 3567 -7536 3579
rect -7570 3545 -7536 3567
rect -7570 3499 -7536 3507
rect -7570 3473 -7536 3499
rect -7474 4417 -7440 4443
rect -7474 4409 -7440 4417
rect -7474 4349 -7440 4371
rect -7474 4337 -7440 4349
rect -7474 4281 -7440 4299
rect -7474 4265 -7440 4281
rect -7474 4213 -7440 4227
rect -7474 4193 -7440 4213
rect -7474 4145 -7440 4155
rect -7474 4121 -7440 4145
rect -7474 4077 -7440 4083
rect -7474 4049 -7440 4077
rect -7474 4009 -7440 4011
rect -7474 3977 -7440 4009
rect -7474 3907 -7440 3939
rect -7474 3905 -7440 3907
rect -7474 3839 -7440 3867
rect -7474 3833 -7440 3839
rect -7474 3771 -7440 3795
rect -7474 3761 -7440 3771
rect -7474 3703 -7440 3723
rect -7474 3689 -7440 3703
rect -7474 3635 -7440 3651
rect -7474 3617 -7440 3635
rect -7474 3567 -7440 3579
rect -7474 3545 -7440 3567
rect -7474 3499 -7440 3507
rect -7474 3473 -7440 3499
rect -7378 4417 -7344 4443
rect -7378 4409 -7344 4417
rect -7378 4349 -7344 4371
rect -7378 4337 -7344 4349
rect -7378 4281 -7344 4299
rect -7378 4265 -7344 4281
rect -7378 4213 -7344 4227
rect -7378 4193 -7344 4213
rect -7378 4145 -7344 4155
rect -7378 4121 -7344 4145
rect -7378 4077 -7344 4083
rect -7378 4049 -7344 4077
rect -7378 4009 -7344 4011
rect -7378 3977 -7344 4009
rect -7378 3907 -7344 3939
rect -7378 3905 -7344 3907
rect -7378 3839 -7344 3867
rect -7378 3833 -7344 3839
rect -7378 3771 -7344 3795
rect -7378 3761 -7344 3771
rect -7378 3703 -7344 3723
rect -7378 3689 -7344 3703
rect -7378 3635 -7344 3651
rect -7378 3617 -7344 3635
rect -7378 3567 -7344 3579
rect -7378 3545 -7344 3567
rect -7378 3499 -7344 3507
rect -7378 3473 -7344 3499
rect -7282 4417 -7248 4443
rect -7282 4409 -7248 4417
rect -7282 4349 -7248 4371
rect -7282 4337 -7248 4349
rect -7282 4281 -7248 4299
rect -7282 4265 -7248 4281
rect -7282 4213 -7248 4227
rect -7282 4193 -7248 4213
rect -7282 4145 -7248 4155
rect -7282 4121 -7248 4145
rect -7282 4077 -7248 4083
rect -7282 4049 -7248 4077
rect -7282 4009 -7248 4011
rect -7282 3977 -7248 4009
rect -7282 3907 -7248 3939
rect -7282 3905 -7248 3907
rect -7282 3839 -7248 3867
rect -7282 3833 -7248 3839
rect -7282 3771 -7248 3795
rect -7282 3761 -7248 3771
rect -7282 3703 -7248 3723
rect -7282 3689 -7248 3703
rect -7282 3635 -7248 3651
rect -7282 3617 -7248 3635
rect -7282 3567 -7248 3579
rect -7282 3545 -7248 3567
rect -7282 3499 -7248 3507
rect -7282 3473 -7248 3499
rect -7186 4417 -7152 4443
rect -7186 4409 -7152 4417
rect -7186 4349 -7152 4371
rect -7186 4337 -7152 4349
rect -7186 4281 -7152 4299
rect -7186 4265 -7152 4281
rect -7186 4213 -7152 4227
rect -7186 4193 -7152 4213
rect -7186 4145 -7152 4155
rect -7186 4121 -7152 4145
rect -7186 4077 -7152 4083
rect -7186 4049 -7152 4077
rect -7186 4009 -7152 4011
rect -7186 3977 -7152 4009
rect -7186 3907 -7152 3939
rect -7186 3905 -7152 3907
rect -7186 3839 -7152 3867
rect -7186 3833 -7152 3839
rect -7186 3771 -7152 3795
rect -7186 3761 -7152 3771
rect -7186 3703 -7152 3723
rect -7186 3689 -7152 3703
rect -7186 3635 -7152 3651
rect -7186 3617 -7152 3635
rect -7186 3567 -7152 3579
rect -7186 3545 -7152 3567
rect -7186 3499 -7152 3507
rect -7186 3473 -7152 3499
rect -7090 4417 -7056 4443
rect -7090 4409 -7056 4417
rect -7090 4349 -7056 4371
rect -7090 4337 -7056 4349
rect -7090 4281 -7056 4299
rect -7090 4265 -7056 4281
rect -7090 4213 -7056 4227
rect -7090 4193 -7056 4213
rect -7090 4145 -7056 4155
rect -7090 4121 -7056 4145
rect -7090 4077 -7056 4083
rect -7090 4049 -7056 4077
rect -7090 4009 -7056 4011
rect -7090 3977 -7056 4009
rect -7090 3907 -7056 3939
rect -7090 3905 -7056 3907
rect -7090 3839 -7056 3867
rect -7090 3833 -7056 3839
rect -7090 3771 -7056 3795
rect -7090 3761 -7056 3771
rect -7090 3703 -7056 3723
rect -7090 3689 -7056 3703
rect -7090 3635 -7056 3651
rect -7090 3617 -7056 3635
rect -7090 3567 -7056 3579
rect -7090 3545 -7056 3567
rect -7090 3499 -7056 3507
rect -7090 3473 -7056 3499
rect -6994 4417 -6960 4443
rect -6994 4409 -6960 4417
rect -6994 4349 -6960 4371
rect -6994 4337 -6960 4349
rect -6994 4281 -6960 4299
rect -6994 4265 -6960 4281
rect -6994 4213 -6960 4227
rect -6994 4193 -6960 4213
rect -6994 4145 -6960 4155
rect -6994 4121 -6960 4145
rect -6994 4077 -6960 4083
rect -6994 4049 -6960 4077
rect -6994 4009 -6960 4011
rect -6994 3977 -6960 4009
rect -6994 3907 -6960 3939
rect -6994 3905 -6960 3907
rect -6994 3839 -6960 3867
rect -6994 3833 -6960 3839
rect -6994 3771 -6960 3795
rect -6994 3761 -6960 3771
rect -6994 3703 -6960 3723
rect -6994 3689 -6960 3703
rect -6994 3635 -6960 3651
rect -6994 3617 -6960 3635
rect -6994 3567 -6960 3579
rect -6994 3545 -6960 3567
rect -6994 3499 -6960 3507
rect -6994 3473 -6960 3499
rect -6898 4417 -6864 4443
rect -6898 4409 -6864 4417
rect -6898 4349 -6864 4371
rect -6898 4337 -6864 4349
rect -6898 4281 -6864 4299
rect -6898 4265 -6864 4281
rect -6898 4213 -6864 4227
rect -6898 4193 -6864 4213
rect -6898 4145 -6864 4155
rect -6898 4121 -6864 4145
rect -6898 4077 -6864 4083
rect -6898 4049 -6864 4077
rect -6898 4009 -6864 4011
rect -6898 3977 -6864 4009
rect -6898 3907 -6864 3939
rect -6898 3905 -6864 3907
rect -6898 3839 -6864 3867
rect -6898 3833 -6864 3839
rect -6898 3771 -6864 3795
rect -6898 3761 -6864 3771
rect -6898 3703 -6864 3723
rect -6898 3689 -6864 3703
rect -6898 3635 -6864 3651
rect -6898 3617 -6864 3635
rect -6898 3567 -6864 3579
rect -6898 3545 -6864 3567
rect -6898 3499 -6864 3507
rect -6898 3473 -6864 3499
rect -6802 4417 -6768 4443
rect -6802 4409 -6768 4417
rect -6802 4349 -6768 4371
rect -6802 4337 -6768 4349
rect -6802 4281 -6768 4299
rect -6802 4265 -6768 4281
rect -6802 4213 -6768 4227
rect -6802 4193 -6768 4213
rect -6802 4145 -6768 4155
rect -6802 4121 -6768 4145
rect -6802 4077 -6768 4083
rect -6802 4049 -6768 4077
rect -6802 4009 -6768 4011
rect -6802 3977 -6768 4009
rect -6802 3907 -6768 3939
rect -6802 3905 -6768 3907
rect -6802 3839 -6768 3867
rect -6802 3833 -6768 3839
rect -6802 3771 -6768 3795
rect -6802 3761 -6768 3771
rect -6802 3703 -6768 3723
rect -6802 3689 -6768 3703
rect -6802 3635 -6768 3651
rect -6802 3617 -6768 3635
rect -6802 3567 -6768 3579
rect -6802 3545 -6768 3567
rect -6802 3499 -6768 3507
rect -6802 3473 -6768 3499
rect -6706 4417 -6672 4443
rect -6706 4409 -6672 4417
rect -6706 4349 -6672 4371
rect -6706 4337 -6672 4349
rect -6706 4281 -6672 4299
rect -6706 4265 -6672 4281
rect -6706 4213 -6672 4227
rect -6706 4193 -6672 4213
rect -6706 4145 -6672 4155
rect -6706 4121 -6672 4145
rect -6706 4077 -6672 4083
rect -6706 4049 -6672 4077
rect -6706 4009 -6672 4011
rect -6706 3977 -6672 4009
rect -6706 3907 -6672 3939
rect -6706 3905 -6672 3907
rect -6706 3839 -6672 3867
rect -6706 3833 -6672 3839
rect -6706 3771 -6672 3795
rect -6706 3761 -6672 3771
rect -6706 3703 -6672 3723
rect -6706 3689 -6672 3703
rect -6706 3635 -6672 3651
rect -6706 3617 -6672 3635
rect -6706 3567 -6672 3579
rect -6706 3545 -6672 3567
rect -6706 3499 -6672 3507
rect -6706 3473 -6672 3499
rect -6462 4423 -6428 4449
rect -6462 4415 -6428 4423
rect -6462 4355 -6428 4377
rect -6462 4343 -6428 4355
rect -6462 4287 -6428 4305
rect -6462 4271 -6428 4287
rect -6462 4219 -6428 4233
rect -6462 4199 -6428 4219
rect -6462 4151 -6428 4161
rect -6462 4127 -6428 4151
rect -6462 4083 -6428 4089
rect -6462 4055 -6428 4083
rect -6462 4015 -6428 4017
rect -6462 3983 -6428 4015
rect -6462 3913 -6428 3945
rect -6462 3911 -6428 3913
rect -6462 3845 -6428 3873
rect -6462 3839 -6428 3845
rect -6462 3777 -6428 3801
rect -6462 3767 -6428 3777
rect -6462 3709 -6428 3729
rect -6462 3695 -6428 3709
rect -6462 3641 -6428 3657
rect -6462 3623 -6428 3641
rect -6462 3573 -6428 3585
rect -6462 3551 -6428 3573
rect -6462 3505 -6428 3513
rect -6462 3479 -6428 3505
rect -6366 4423 -6332 4449
rect -6366 4415 -6332 4423
rect -6366 4355 -6332 4377
rect -6366 4343 -6332 4355
rect -6366 4287 -6332 4305
rect -6366 4271 -6332 4287
rect -6366 4219 -6332 4233
rect -6366 4199 -6332 4219
rect -6366 4151 -6332 4161
rect -6366 4127 -6332 4151
rect -6366 4083 -6332 4089
rect -6366 4055 -6332 4083
rect -6366 4015 -6332 4017
rect -6366 3983 -6332 4015
rect -6366 3913 -6332 3945
rect -6366 3911 -6332 3913
rect -6366 3845 -6332 3873
rect -6366 3839 -6332 3845
rect -6366 3777 -6332 3801
rect -6366 3767 -6332 3777
rect -6366 3709 -6332 3729
rect -6366 3695 -6332 3709
rect -6366 3641 -6332 3657
rect -6366 3623 -6332 3641
rect -6366 3573 -6332 3585
rect -6366 3551 -6332 3573
rect -6366 3505 -6332 3513
rect -6366 3479 -6332 3505
rect -11328 3247 -11294 3281
rect -11472 3125 -11438 3159
rect -12020 3040 -11986 3074
rect -20000 2805 -19966 2831
rect -20000 2797 -19966 2805
rect -20000 2737 -19966 2759
rect -20000 2725 -19966 2737
rect -20000 2669 -19966 2687
rect -20000 2653 -19966 2669
rect -20000 2601 -19966 2615
rect -20000 2581 -19966 2601
rect -20000 2533 -19966 2543
rect -20000 2509 -19966 2533
rect -20000 2465 -19966 2471
rect -20000 2437 -19966 2465
rect -20000 2397 -19966 2399
rect -20000 2365 -19966 2397
rect -20000 2295 -19966 2327
rect -20000 2293 -19966 2295
rect -20000 2227 -19966 2255
rect -20000 2221 -19966 2227
rect -20000 2159 -19966 2183
rect -20000 2149 -19966 2159
rect -20000 2091 -19966 2111
rect -20000 2077 -19966 2091
rect -20000 2023 -19966 2039
rect -20000 2005 -19966 2023
rect -20000 1955 -19966 1967
rect -20000 1933 -19966 1955
rect -20000 1887 -19966 1895
rect -20000 1861 -19966 1887
rect -19904 2805 -19870 2831
rect -19904 2797 -19870 2805
rect -19904 2737 -19870 2759
rect -19904 2725 -19870 2737
rect -19904 2669 -19870 2687
rect -19904 2653 -19870 2669
rect -19904 2601 -19870 2615
rect -19904 2581 -19870 2601
rect -19904 2533 -19870 2543
rect -19904 2509 -19870 2533
rect -19904 2465 -19870 2471
rect -19904 2437 -19870 2465
rect -19904 2397 -19870 2399
rect -19904 2365 -19870 2397
rect -19904 2295 -19870 2327
rect -19904 2293 -19870 2295
rect -19904 2227 -19870 2255
rect -19904 2221 -19870 2227
rect -19904 2159 -19870 2183
rect -19904 2149 -19870 2159
rect -19904 2091 -19870 2111
rect -19904 2077 -19870 2091
rect -19904 2023 -19870 2039
rect -19904 2005 -19870 2023
rect -19904 1955 -19870 1967
rect -19904 1933 -19870 1955
rect -19904 1887 -19870 1895
rect -19904 1861 -19870 1887
rect -19666 2809 -19632 2835
rect -19666 2801 -19632 2809
rect -19666 2741 -19632 2763
rect -19666 2729 -19632 2741
rect -19666 2673 -19632 2691
rect -19666 2657 -19632 2673
rect -19666 2605 -19632 2619
rect -19666 2585 -19632 2605
rect -19666 2537 -19632 2547
rect -19666 2513 -19632 2537
rect -19666 2469 -19632 2475
rect -19666 2441 -19632 2469
rect -19666 2401 -19632 2403
rect -19666 2369 -19632 2401
rect -19666 2299 -19632 2331
rect -19666 2297 -19632 2299
rect -19666 2231 -19632 2259
rect -19666 2225 -19632 2231
rect -19666 2163 -19632 2187
rect -19666 2153 -19632 2163
rect -19666 2095 -19632 2115
rect -19666 2081 -19632 2095
rect -19666 2027 -19632 2043
rect -19666 2009 -19632 2027
rect -19666 1959 -19632 1971
rect -19666 1937 -19632 1959
rect -19666 1891 -19632 1899
rect -19666 1865 -19632 1891
rect -19570 2809 -19536 2835
rect -19570 2801 -19536 2809
rect -19570 2741 -19536 2763
rect -19570 2729 -19536 2741
rect -19570 2673 -19536 2691
rect -19570 2657 -19536 2673
rect -19570 2605 -19536 2619
rect -19570 2585 -19536 2605
rect -19570 2537 -19536 2547
rect -19570 2513 -19536 2537
rect -19570 2469 -19536 2475
rect -19570 2441 -19536 2469
rect -19570 2401 -19536 2403
rect -19570 2369 -19536 2401
rect -19570 2299 -19536 2331
rect -19570 2297 -19536 2299
rect -19570 2231 -19536 2259
rect -19570 2225 -19536 2231
rect -19570 2163 -19536 2187
rect -19570 2153 -19536 2163
rect -19570 2095 -19536 2115
rect -19570 2081 -19536 2095
rect -19570 2027 -19536 2043
rect -19570 2009 -19536 2027
rect -19570 1959 -19536 1971
rect -19570 1937 -19536 1959
rect -19570 1891 -19536 1899
rect -19570 1865 -19536 1891
rect -19474 2809 -19440 2835
rect -19474 2801 -19440 2809
rect -19474 2741 -19440 2763
rect -19474 2729 -19440 2741
rect -19474 2673 -19440 2691
rect -19474 2657 -19440 2673
rect -19474 2605 -19440 2619
rect -19474 2585 -19440 2605
rect -19474 2537 -19440 2547
rect -19474 2513 -19440 2537
rect -19474 2469 -19440 2475
rect -19474 2441 -19440 2469
rect -19474 2401 -19440 2403
rect -19474 2369 -19440 2401
rect -19474 2299 -19440 2331
rect -19474 2297 -19440 2299
rect -19474 2231 -19440 2259
rect -19474 2225 -19440 2231
rect -19474 2163 -19440 2187
rect -19474 2153 -19440 2163
rect -19474 2095 -19440 2115
rect -19474 2081 -19440 2095
rect -19474 2027 -19440 2043
rect -19474 2009 -19440 2027
rect -19474 1959 -19440 1971
rect -19474 1937 -19440 1959
rect -19474 1891 -19440 1899
rect -19474 1865 -19440 1891
rect -19378 2809 -19344 2835
rect -19378 2801 -19344 2809
rect -19378 2741 -19344 2763
rect -19378 2729 -19344 2741
rect -19378 2673 -19344 2691
rect -19378 2657 -19344 2673
rect -19378 2605 -19344 2619
rect -19378 2585 -19344 2605
rect -19378 2537 -19344 2547
rect -19378 2513 -19344 2537
rect -19378 2469 -19344 2475
rect -19378 2441 -19344 2469
rect -19378 2401 -19344 2403
rect -19378 2369 -19344 2401
rect -19378 2299 -19344 2331
rect -19378 2297 -19344 2299
rect -19378 2231 -19344 2259
rect -19378 2225 -19344 2231
rect -19378 2163 -19344 2187
rect -19378 2153 -19344 2163
rect -19378 2095 -19344 2115
rect -19378 2081 -19344 2095
rect -19378 2027 -19344 2043
rect -19378 2009 -19344 2027
rect -19378 1959 -19344 1971
rect -19378 1937 -19344 1959
rect -19378 1891 -19344 1899
rect -19378 1865 -19344 1891
rect -19282 2809 -19248 2835
rect -19282 2801 -19248 2809
rect -19282 2741 -19248 2763
rect -19282 2729 -19248 2741
rect -19282 2673 -19248 2691
rect -19282 2657 -19248 2673
rect -19282 2605 -19248 2619
rect -19282 2585 -19248 2605
rect -19282 2537 -19248 2547
rect -19282 2513 -19248 2537
rect -19282 2469 -19248 2475
rect -19282 2441 -19248 2469
rect -19282 2401 -19248 2403
rect -19282 2369 -19248 2401
rect -19282 2299 -19248 2331
rect -19282 2297 -19248 2299
rect -19282 2231 -19248 2259
rect -19282 2225 -19248 2231
rect -19282 2163 -19248 2187
rect -19282 2153 -19248 2163
rect -19282 2095 -19248 2115
rect -19282 2081 -19248 2095
rect -19282 2027 -19248 2043
rect -19282 2009 -19248 2027
rect -19282 1959 -19248 1971
rect -19282 1937 -19248 1959
rect -19282 1891 -19248 1899
rect -19282 1865 -19248 1891
rect -19186 2809 -19152 2835
rect -19186 2801 -19152 2809
rect -19186 2741 -19152 2763
rect -19186 2729 -19152 2741
rect -19186 2673 -19152 2691
rect -19186 2657 -19152 2673
rect -19186 2605 -19152 2619
rect -19186 2585 -19152 2605
rect -19186 2537 -19152 2547
rect -19186 2513 -19152 2537
rect -19186 2469 -19152 2475
rect -19186 2441 -19152 2469
rect -19186 2401 -19152 2403
rect -19186 2369 -19152 2401
rect -19186 2299 -19152 2331
rect -19186 2297 -19152 2299
rect -19186 2231 -19152 2259
rect -19186 2225 -19152 2231
rect -19186 2163 -19152 2187
rect -19186 2153 -19152 2163
rect -19186 2095 -19152 2115
rect -19186 2081 -19152 2095
rect -19186 2027 -19152 2043
rect -19186 2009 -19152 2027
rect -19186 1959 -19152 1971
rect -19186 1937 -19152 1959
rect -19186 1891 -19152 1899
rect -19186 1865 -19152 1891
rect -19090 2809 -19056 2835
rect -19090 2801 -19056 2809
rect -19090 2741 -19056 2763
rect -19090 2729 -19056 2741
rect -19090 2673 -19056 2691
rect -19090 2657 -19056 2673
rect -19090 2605 -19056 2619
rect -19090 2585 -19056 2605
rect -19090 2537 -19056 2547
rect -19090 2513 -19056 2537
rect -19090 2469 -19056 2475
rect -19090 2441 -19056 2469
rect -19090 2401 -19056 2403
rect -19090 2369 -19056 2401
rect -19090 2299 -19056 2331
rect -19090 2297 -19056 2299
rect -19090 2231 -19056 2259
rect -19090 2225 -19056 2231
rect -19090 2163 -19056 2187
rect -19090 2153 -19056 2163
rect -19090 2095 -19056 2115
rect -19090 2081 -19056 2095
rect -19090 2027 -19056 2043
rect -19090 2009 -19056 2027
rect -19090 1959 -19056 1971
rect -19090 1937 -19056 1959
rect -19090 1891 -19056 1899
rect -19090 1865 -19056 1891
rect -18994 2809 -18960 2835
rect -18994 2801 -18960 2809
rect -18994 2741 -18960 2763
rect -18994 2729 -18960 2741
rect -18994 2673 -18960 2691
rect -18994 2657 -18960 2673
rect -18994 2605 -18960 2619
rect -18994 2585 -18960 2605
rect -18994 2537 -18960 2547
rect -18994 2513 -18960 2537
rect -18994 2469 -18960 2475
rect -18994 2441 -18960 2469
rect -18994 2401 -18960 2403
rect -18994 2369 -18960 2401
rect -18994 2299 -18960 2331
rect -18994 2297 -18960 2299
rect -18994 2231 -18960 2259
rect -18994 2225 -18960 2231
rect -18994 2163 -18960 2187
rect -18994 2153 -18960 2163
rect -18994 2095 -18960 2115
rect -18994 2081 -18960 2095
rect -18994 2027 -18960 2043
rect -18994 2009 -18960 2027
rect -18994 1959 -18960 1971
rect -18994 1937 -18960 1959
rect -18994 1891 -18960 1899
rect -18994 1865 -18960 1891
rect -18898 2809 -18864 2835
rect -18898 2801 -18864 2809
rect -18898 2741 -18864 2763
rect -18898 2729 -18864 2741
rect -18898 2673 -18864 2691
rect -18898 2657 -18864 2673
rect -18898 2605 -18864 2619
rect -18898 2585 -18864 2605
rect -18898 2537 -18864 2547
rect -18898 2513 -18864 2537
rect -18898 2469 -18864 2475
rect -18898 2441 -18864 2469
rect -18898 2401 -18864 2403
rect -18898 2369 -18864 2401
rect -18898 2299 -18864 2331
rect -18898 2297 -18864 2299
rect -18898 2231 -18864 2259
rect -18898 2225 -18864 2231
rect -18898 2163 -18864 2187
rect -18898 2153 -18864 2163
rect -18898 2095 -18864 2115
rect -18898 2081 -18864 2095
rect -18898 2027 -18864 2043
rect -18898 2009 -18864 2027
rect -18898 1959 -18864 1971
rect -18898 1937 -18864 1959
rect -18898 1891 -18864 1899
rect -18898 1865 -18864 1891
rect -18802 2809 -18768 2835
rect -18802 2801 -18768 2809
rect -18802 2741 -18768 2763
rect -18802 2729 -18768 2741
rect -18802 2673 -18768 2691
rect -18802 2657 -18768 2673
rect -18802 2605 -18768 2619
rect -18802 2585 -18768 2605
rect -18802 2537 -18768 2547
rect -18802 2513 -18768 2537
rect -18802 2469 -18768 2475
rect -18802 2441 -18768 2469
rect -18802 2401 -18768 2403
rect -18802 2369 -18768 2401
rect -18802 2299 -18768 2331
rect -18802 2297 -18768 2299
rect -18802 2231 -18768 2259
rect -18802 2225 -18768 2231
rect -18802 2163 -18768 2187
rect -18802 2153 -18768 2163
rect -18802 2095 -18768 2115
rect -18802 2081 -18768 2095
rect -18802 2027 -18768 2043
rect -18802 2009 -18768 2027
rect -18802 1959 -18768 1971
rect -18802 1937 -18768 1959
rect -18802 1891 -18768 1899
rect -18802 1865 -18768 1891
rect -18706 2809 -18672 2835
rect -18706 2801 -18672 2809
rect -18706 2741 -18672 2763
rect -18706 2729 -18672 2741
rect -18706 2673 -18672 2691
rect -18706 2657 -18672 2673
rect -18706 2605 -18672 2619
rect -18706 2585 -18672 2605
rect -18706 2537 -18672 2547
rect -18706 2513 -18672 2537
rect -18706 2469 -18672 2475
rect -18706 2441 -18672 2469
rect -18706 2401 -18672 2403
rect -18706 2369 -18672 2401
rect -18706 2299 -18672 2331
rect -18706 2297 -18672 2299
rect -18706 2231 -18672 2259
rect -18706 2225 -18672 2231
rect -18706 2163 -18672 2187
rect -18706 2153 -18672 2163
rect -18706 2095 -18672 2115
rect -18706 2081 -18672 2095
rect -18706 2027 -18672 2043
rect -18706 2009 -18672 2027
rect -18706 1959 -18672 1971
rect -18706 1937 -18672 1959
rect -18706 1891 -18672 1899
rect -18706 1865 -18672 1891
rect -18494 2819 -18460 2845
rect -18494 2811 -18460 2819
rect -18494 2751 -18460 2773
rect -18494 2739 -18460 2751
rect -18494 2683 -18460 2701
rect -18494 2667 -18460 2683
rect -18494 2615 -18460 2629
rect -18494 2595 -18460 2615
rect -18494 2547 -18460 2557
rect -18494 2523 -18460 2547
rect -18494 2479 -18460 2485
rect -18494 2451 -18460 2479
rect -18494 2411 -18460 2413
rect -18494 2379 -18460 2411
rect -18494 2309 -18460 2341
rect -18494 2307 -18460 2309
rect -18494 2241 -18460 2269
rect -18494 2235 -18460 2241
rect -18494 2173 -18460 2197
rect -18494 2163 -18460 2173
rect -18494 2105 -18460 2125
rect -18494 2091 -18460 2105
rect -18494 2037 -18460 2053
rect -18494 2019 -18460 2037
rect -18494 1969 -18460 1981
rect -18494 1947 -18460 1969
rect -18494 1901 -18460 1909
rect -18494 1875 -18460 1901
rect -18398 2819 -18364 2845
rect -18398 2811 -18364 2819
rect -18398 2751 -18364 2773
rect -18398 2739 -18364 2751
rect -18398 2683 -18364 2701
rect -18398 2667 -18364 2683
rect -18398 2615 -18364 2629
rect -18398 2595 -18364 2615
rect -18398 2547 -18364 2557
rect -18398 2523 -18364 2547
rect -18398 2479 -18364 2485
rect -18398 2451 -18364 2479
rect -18398 2411 -18364 2413
rect -18398 2379 -18364 2411
rect -18398 2309 -18364 2341
rect -18398 2307 -18364 2309
rect -18398 2241 -18364 2269
rect -18398 2235 -18364 2241
rect -18398 2173 -18364 2197
rect -18398 2163 -18364 2173
rect -18398 2105 -18364 2125
rect -18398 2091 -18364 2105
rect -18398 2037 -18364 2053
rect -18398 2019 -18364 2037
rect -18398 1969 -18364 1981
rect -18398 1947 -18364 1969
rect -18398 1901 -18364 1909
rect -18398 1875 -18364 1901
rect -18302 2819 -18268 2845
rect -18302 2811 -18268 2819
rect -18302 2751 -18268 2773
rect -18302 2739 -18268 2751
rect -18302 2683 -18268 2701
rect -18302 2667 -18268 2683
rect -18302 2615 -18268 2629
rect -18302 2595 -18268 2615
rect -18302 2547 -18268 2557
rect -18302 2523 -18268 2547
rect -18302 2479 -18268 2485
rect -18302 2451 -18268 2479
rect -18302 2411 -18268 2413
rect -18302 2379 -18268 2411
rect -18302 2309 -18268 2341
rect -18302 2307 -18268 2309
rect -18302 2241 -18268 2269
rect -18302 2235 -18268 2241
rect -18302 2173 -18268 2197
rect -18302 2163 -18268 2173
rect -18302 2105 -18268 2125
rect -18302 2091 -18268 2105
rect -18302 2037 -18268 2053
rect -18302 2019 -18268 2037
rect -18302 1969 -18268 1981
rect -18302 1947 -18268 1969
rect -18302 1901 -18268 1909
rect -18302 1875 -18268 1901
rect -18206 2819 -18172 2845
rect -18206 2811 -18172 2819
rect -18206 2751 -18172 2773
rect -18206 2739 -18172 2751
rect -18206 2683 -18172 2701
rect -18206 2667 -18172 2683
rect -18206 2615 -18172 2629
rect -18206 2595 -18172 2615
rect -18206 2547 -18172 2557
rect -18206 2523 -18172 2547
rect -18206 2479 -18172 2485
rect -18206 2451 -18172 2479
rect -18206 2411 -18172 2413
rect -18206 2379 -18172 2411
rect -18206 2309 -18172 2341
rect -18206 2307 -18172 2309
rect -18206 2241 -18172 2269
rect -18206 2235 -18172 2241
rect -18206 2173 -18172 2197
rect -18206 2163 -18172 2173
rect -18206 2105 -18172 2125
rect -18206 2091 -18172 2105
rect -18206 2037 -18172 2053
rect -18206 2019 -18172 2037
rect -18206 1969 -18172 1981
rect -18206 1947 -18172 1969
rect -18206 1901 -18172 1909
rect -18206 1875 -18172 1901
rect -18110 2819 -18076 2845
rect -18110 2811 -18076 2819
rect -18110 2751 -18076 2773
rect -18110 2739 -18076 2751
rect -18110 2683 -18076 2701
rect -18110 2667 -18076 2683
rect -18110 2615 -18076 2629
rect -18110 2595 -18076 2615
rect -18110 2547 -18076 2557
rect -18110 2523 -18076 2547
rect -18110 2479 -18076 2485
rect -18110 2451 -18076 2479
rect -18110 2411 -18076 2413
rect -18110 2379 -18076 2411
rect -18110 2309 -18076 2341
rect -18110 2307 -18076 2309
rect -18110 2241 -18076 2269
rect -18110 2235 -18076 2241
rect -18110 2173 -18076 2197
rect -18110 2163 -18076 2173
rect -18110 2105 -18076 2125
rect -18110 2091 -18076 2105
rect -18110 2037 -18076 2053
rect -18110 2019 -18076 2037
rect -18110 1969 -18076 1981
rect -18110 1947 -18076 1969
rect -18110 1901 -18076 1909
rect -18110 1875 -18076 1901
rect -18014 2819 -17980 2845
rect -18014 2811 -17980 2819
rect -18014 2751 -17980 2773
rect -18014 2739 -17980 2751
rect -18014 2683 -17980 2701
rect -18014 2667 -17980 2683
rect -18014 2615 -17980 2629
rect -18014 2595 -17980 2615
rect -18014 2547 -17980 2557
rect -18014 2523 -17980 2547
rect -18014 2479 -17980 2485
rect -18014 2451 -17980 2479
rect -18014 2411 -17980 2413
rect -18014 2379 -17980 2411
rect -18014 2309 -17980 2341
rect -18014 2307 -17980 2309
rect -18014 2241 -17980 2269
rect -18014 2235 -17980 2241
rect -18014 2173 -17980 2197
rect -18014 2163 -17980 2173
rect -18014 2105 -17980 2125
rect -18014 2091 -17980 2105
rect -18014 2037 -17980 2053
rect -18014 2019 -17980 2037
rect -18014 1969 -17980 1981
rect -18014 1947 -17980 1969
rect -18014 1901 -17980 1909
rect -18014 1875 -17980 1901
rect -16662 2825 -16628 2851
rect -16662 2817 -16628 2825
rect -16662 2757 -16628 2779
rect -16662 2745 -16628 2757
rect -16662 2689 -16628 2707
rect -16662 2673 -16628 2689
rect -16662 2621 -16628 2635
rect -16662 2601 -16628 2621
rect -16662 2553 -16628 2563
rect -16662 2529 -16628 2553
rect -16662 2485 -16628 2491
rect -16662 2457 -16628 2485
rect -16662 2417 -16628 2419
rect -16662 2385 -16628 2417
rect -16662 2315 -16628 2347
rect -16662 2313 -16628 2315
rect -16662 2247 -16628 2275
rect -16662 2241 -16628 2247
rect -16662 2179 -16628 2203
rect -16662 2169 -16628 2179
rect -16662 2111 -16628 2131
rect -16662 2097 -16628 2111
rect -16662 2043 -16628 2059
rect -16662 2025 -16628 2043
rect -16662 1975 -16628 1987
rect -16662 1953 -16628 1975
rect -16662 1907 -16628 1915
rect -16662 1881 -16628 1907
rect -16566 2825 -16532 2851
rect -16566 2817 -16532 2825
rect -16566 2757 -16532 2779
rect -16566 2745 -16532 2757
rect -16566 2689 -16532 2707
rect -16566 2673 -16532 2689
rect -16566 2621 -16532 2635
rect -16566 2601 -16532 2621
rect -16566 2553 -16532 2563
rect -16566 2529 -16532 2553
rect -16566 2485 -16532 2491
rect -16566 2457 -16532 2485
rect -16566 2417 -16532 2419
rect -16566 2385 -16532 2417
rect -16566 2315 -16532 2347
rect -16566 2313 -16532 2315
rect -16566 2247 -16532 2275
rect -16566 2241 -16532 2247
rect -16566 2179 -16532 2203
rect -16566 2169 -16532 2179
rect -16566 2111 -16532 2131
rect -16566 2097 -16532 2111
rect -16566 2043 -16532 2059
rect -16566 2025 -16532 2043
rect -16566 1975 -16532 1987
rect -16566 1953 -16532 1975
rect -16566 1907 -16532 1915
rect -16566 1881 -16532 1907
rect -16470 2825 -16436 2851
rect -16470 2817 -16436 2825
rect -16470 2757 -16436 2779
rect -16470 2745 -16436 2757
rect -16470 2689 -16436 2707
rect -16470 2673 -16436 2689
rect -16470 2621 -16436 2635
rect -16470 2601 -16436 2621
rect -16470 2553 -16436 2563
rect -16470 2529 -16436 2553
rect -16470 2485 -16436 2491
rect -16470 2457 -16436 2485
rect -16470 2417 -16436 2419
rect -16470 2385 -16436 2417
rect -16470 2315 -16436 2347
rect -16470 2313 -16436 2315
rect -16470 2247 -16436 2275
rect -16470 2241 -16436 2247
rect -16470 2179 -16436 2203
rect -16470 2169 -16436 2179
rect -16470 2111 -16436 2131
rect -16470 2097 -16436 2111
rect -16470 2043 -16436 2059
rect -16470 2025 -16436 2043
rect -16470 1975 -16436 1987
rect -16470 1953 -16436 1975
rect -16470 1907 -16436 1915
rect -16470 1881 -16436 1907
rect -16374 2825 -16340 2851
rect -16374 2817 -16340 2825
rect -16374 2757 -16340 2779
rect -16374 2745 -16340 2757
rect -16374 2689 -16340 2707
rect -16374 2673 -16340 2689
rect -16374 2621 -16340 2635
rect -16374 2601 -16340 2621
rect -16374 2553 -16340 2563
rect -16374 2529 -16340 2553
rect -16374 2485 -16340 2491
rect -16374 2457 -16340 2485
rect -16374 2417 -16340 2419
rect -16374 2385 -16340 2417
rect -16374 2315 -16340 2347
rect -16374 2313 -16340 2315
rect -16374 2247 -16340 2275
rect -16374 2241 -16340 2247
rect -16374 2179 -16340 2203
rect -16374 2169 -16340 2179
rect -16374 2111 -16340 2131
rect -16374 2097 -16340 2111
rect -16374 2043 -16340 2059
rect -16374 2025 -16340 2043
rect -16374 1975 -16340 1987
rect -16374 1953 -16340 1975
rect -16374 1907 -16340 1915
rect -16374 1881 -16340 1907
rect -16278 2825 -16244 2851
rect -16278 2817 -16244 2825
rect -16278 2757 -16244 2779
rect -16278 2745 -16244 2757
rect -16278 2689 -16244 2707
rect -16278 2673 -16244 2689
rect -16278 2621 -16244 2635
rect -16278 2601 -16244 2621
rect -16278 2553 -16244 2563
rect -16278 2529 -16244 2553
rect -16278 2485 -16244 2491
rect -16278 2457 -16244 2485
rect -16278 2417 -16244 2419
rect -16278 2385 -16244 2417
rect -16278 2315 -16244 2347
rect -16278 2313 -16244 2315
rect -16278 2247 -16244 2275
rect -16278 2241 -16244 2247
rect -16278 2179 -16244 2203
rect -16278 2169 -16244 2179
rect -16278 2111 -16244 2131
rect -16278 2097 -16244 2111
rect -16278 2043 -16244 2059
rect -16278 2025 -16244 2043
rect -16278 1975 -16244 1987
rect -16278 1953 -16244 1975
rect -16278 1907 -16244 1915
rect -16278 1881 -16244 1907
rect -16182 2825 -16148 2851
rect -16182 2817 -16148 2825
rect -16182 2757 -16148 2779
rect -16182 2745 -16148 2757
rect -16182 2689 -16148 2707
rect -16182 2673 -16148 2689
rect -16182 2621 -16148 2635
rect -16182 2601 -16148 2621
rect -16182 2553 -16148 2563
rect -16182 2529 -16148 2553
rect -16182 2485 -16148 2491
rect -16182 2457 -16148 2485
rect -16182 2417 -16148 2419
rect -16182 2385 -16148 2417
rect -16182 2315 -16148 2347
rect -16182 2313 -16148 2315
rect -16182 2247 -16148 2275
rect -16182 2241 -16148 2247
rect -16182 2179 -16148 2203
rect -16182 2169 -16148 2179
rect -16182 2111 -16148 2131
rect -16182 2097 -16148 2111
rect -16182 2043 -16148 2059
rect -16182 2025 -16148 2043
rect -16182 1975 -16148 1987
rect -16182 1953 -16148 1975
rect -16182 1907 -16148 1915
rect -16182 1881 -16148 1907
rect -16086 2825 -16052 2851
rect -16086 2817 -16052 2825
rect -16086 2757 -16052 2779
rect -16086 2745 -16052 2757
rect -16086 2689 -16052 2707
rect -16086 2673 -16052 2689
rect -16086 2621 -16052 2635
rect -16086 2601 -16052 2621
rect -16086 2553 -16052 2563
rect -16086 2529 -16052 2553
rect -16086 2485 -16052 2491
rect -16086 2457 -16052 2485
rect -16086 2417 -16052 2419
rect -16086 2385 -16052 2417
rect -16086 2315 -16052 2347
rect -16086 2313 -16052 2315
rect -16086 2247 -16052 2275
rect -16086 2241 -16052 2247
rect -16086 2179 -16052 2203
rect -16086 2169 -16052 2179
rect -16086 2111 -16052 2131
rect -16086 2097 -16052 2111
rect -16086 2043 -16052 2059
rect -16086 2025 -16052 2043
rect -16086 1975 -16052 1987
rect -16086 1953 -16052 1975
rect -16086 1907 -16052 1915
rect -16086 1881 -16052 1907
rect -15990 2825 -15956 2851
rect -15990 2817 -15956 2825
rect -15990 2757 -15956 2779
rect -15990 2745 -15956 2757
rect -15990 2689 -15956 2707
rect -15990 2673 -15956 2689
rect -15990 2621 -15956 2635
rect -15990 2601 -15956 2621
rect -15990 2553 -15956 2563
rect -15990 2529 -15956 2553
rect -15990 2485 -15956 2491
rect -15990 2457 -15956 2485
rect -15990 2417 -15956 2419
rect -15990 2385 -15956 2417
rect -15990 2315 -15956 2347
rect -15990 2313 -15956 2315
rect -15990 2247 -15956 2275
rect -15990 2241 -15956 2247
rect -15990 2179 -15956 2203
rect -15990 2169 -15956 2179
rect -15990 2111 -15956 2131
rect -15990 2097 -15956 2111
rect -15990 2043 -15956 2059
rect -15990 2025 -15956 2043
rect -15990 1975 -15956 1987
rect -15990 1953 -15956 1975
rect -15990 1907 -15956 1915
rect -15990 1881 -15956 1907
rect -15894 2825 -15860 2851
rect -15894 2817 -15860 2825
rect -15894 2757 -15860 2779
rect -15894 2745 -15860 2757
rect -15894 2689 -15860 2707
rect -15894 2673 -15860 2689
rect -15894 2621 -15860 2635
rect -15894 2601 -15860 2621
rect -15894 2553 -15860 2563
rect -15894 2529 -15860 2553
rect -15894 2485 -15860 2491
rect -15894 2457 -15860 2485
rect -15894 2417 -15860 2419
rect -15894 2385 -15860 2417
rect -15894 2315 -15860 2347
rect -15894 2313 -15860 2315
rect -15894 2247 -15860 2275
rect -15894 2241 -15860 2247
rect -15894 2179 -15860 2203
rect -15894 2169 -15860 2179
rect -15894 2111 -15860 2131
rect -15894 2097 -15860 2111
rect -15894 2043 -15860 2059
rect -15894 2025 -15860 2043
rect -15894 1975 -15860 1987
rect -15894 1953 -15860 1975
rect -15894 1907 -15860 1915
rect -15894 1881 -15860 1907
rect -15798 2825 -15764 2851
rect -15798 2817 -15764 2825
rect -15798 2757 -15764 2779
rect -15798 2745 -15764 2757
rect -15798 2689 -15764 2707
rect -15798 2673 -15764 2689
rect -15798 2621 -15764 2635
rect -15798 2601 -15764 2621
rect -15798 2553 -15764 2563
rect -15798 2529 -15764 2553
rect -15798 2485 -15764 2491
rect -15798 2457 -15764 2485
rect -15798 2417 -15764 2419
rect -15798 2385 -15764 2417
rect -15798 2315 -15764 2347
rect -15798 2313 -15764 2315
rect -15798 2247 -15764 2275
rect -15798 2241 -15764 2247
rect -15798 2179 -15764 2203
rect -15798 2169 -15764 2179
rect -15798 2111 -15764 2131
rect -15798 2097 -15764 2111
rect -15798 2043 -15764 2059
rect -15798 2025 -15764 2043
rect -15798 1975 -15764 1987
rect -15798 1953 -15764 1975
rect -15798 1907 -15764 1915
rect -15798 1881 -15764 1907
rect -15702 2825 -15668 2851
rect -15702 2817 -15668 2825
rect -15702 2757 -15668 2779
rect -15702 2745 -15668 2757
rect -15702 2689 -15668 2707
rect -15702 2673 -15668 2689
rect -15702 2621 -15668 2635
rect -15702 2601 -15668 2621
rect -15702 2553 -15668 2563
rect -15702 2529 -15668 2553
rect -15702 2485 -15668 2491
rect -15702 2457 -15668 2485
rect -15702 2417 -15668 2419
rect -15702 2385 -15668 2417
rect -15702 2315 -15668 2347
rect -15702 2313 -15668 2315
rect -15702 2247 -15668 2275
rect -15702 2241 -15668 2247
rect -15702 2179 -15668 2203
rect -15702 2169 -15668 2179
rect -15702 2111 -15668 2131
rect -15702 2097 -15668 2111
rect -15702 2043 -15668 2059
rect -15702 2025 -15668 2043
rect -15702 1975 -15668 1987
rect -15702 1953 -15668 1975
rect -15702 1907 -15668 1915
rect -15702 1881 -15668 1907
rect -15606 2825 -15572 2851
rect -15606 2817 -15572 2825
rect -15606 2757 -15572 2779
rect -15606 2745 -15572 2757
rect -15606 2689 -15572 2707
rect -15606 2673 -15572 2689
rect -15606 2621 -15572 2635
rect -15606 2601 -15572 2621
rect -15606 2553 -15572 2563
rect -15606 2529 -15572 2553
rect -15606 2485 -15572 2491
rect -15606 2457 -15572 2485
rect -15606 2417 -15572 2419
rect -15606 2385 -15572 2417
rect -15606 2315 -15572 2347
rect -15606 2313 -15572 2315
rect -15606 2247 -15572 2275
rect -15606 2241 -15572 2247
rect -15606 2179 -15572 2203
rect -15606 2169 -15572 2179
rect -15606 2111 -15572 2131
rect -15606 2097 -15572 2111
rect -15606 2043 -15572 2059
rect -15606 2025 -15572 2043
rect -15606 1975 -15572 1987
rect -15606 1953 -15572 1975
rect -15606 1907 -15572 1915
rect -15606 1881 -15572 1907
rect -15510 2825 -15476 2851
rect -15510 2817 -15476 2825
rect -15510 2757 -15476 2779
rect -15510 2745 -15476 2757
rect -15510 2689 -15476 2707
rect -15510 2673 -15476 2689
rect -15510 2621 -15476 2635
rect -15510 2601 -15476 2621
rect -15510 2553 -15476 2563
rect -15510 2529 -15476 2553
rect -15510 2485 -15476 2491
rect -15510 2457 -15476 2485
rect -15510 2417 -15476 2419
rect -15510 2385 -15476 2417
rect -15510 2315 -15476 2347
rect -15510 2313 -15476 2315
rect -15510 2247 -15476 2275
rect -15510 2241 -15476 2247
rect -15510 2179 -15476 2203
rect -15510 2169 -15476 2179
rect -15510 2111 -15476 2131
rect -15510 2097 -15476 2111
rect -15510 2043 -15476 2059
rect -15510 2025 -15476 2043
rect -15510 1975 -15476 1987
rect -15510 1953 -15476 1975
rect -15510 1907 -15476 1915
rect -15510 1881 -15476 1907
rect -15414 2825 -15380 2851
rect -15414 2817 -15380 2825
rect -15414 2757 -15380 2779
rect -15414 2745 -15380 2757
rect -15414 2689 -15380 2707
rect -15414 2673 -15380 2689
rect -15414 2621 -15380 2635
rect -15414 2601 -15380 2621
rect -15414 2553 -15380 2563
rect -15414 2529 -15380 2553
rect -15414 2485 -15380 2491
rect -15414 2457 -15380 2485
rect -15414 2417 -15380 2419
rect -15414 2385 -15380 2417
rect -15414 2315 -15380 2347
rect -15414 2313 -15380 2315
rect -15414 2247 -15380 2275
rect -15414 2241 -15380 2247
rect -15414 2179 -15380 2203
rect -15414 2169 -15380 2179
rect -15414 2111 -15380 2131
rect -15414 2097 -15380 2111
rect -15414 2043 -15380 2059
rect -15414 2025 -15380 2043
rect -15414 1975 -15380 1987
rect -15414 1953 -15380 1975
rect -15414 1907 -15380 1915
rect -15414 1881 -15380 1907
rect -15318 2825 -15284 2851
rect -15318 2817 -15284 2825
rect -15318 2757 -15284 2779
rect -15318 2745 -15284 2757
rect -15318 2689 -15284 2707
rect -15318 2673 -15284 2689
rect -15318 2621 -15284 2635
rect -15318 2601 -15284 2621
rect -15318 2553 -15284 2563
rect -15318 2529 -15284 2553
rect -15318 2485 -15284 2491
rect -15318 2457 -15284 2485
rect -15318 2417 -15284 2419
rect -15318 2385 -15284 2417
rect -15318 2315 -15284 2347
rect -15318 2313 -15284 2315
rect -15318 2247 -15284 2275
rect -15318 2241 -15284 2247
rect -15318 2179 -15284 2203
rect -15318 2169 -15284 2179
rect -15318 2111 -15284 2131
rect -15318 2097 -15284 2111
rect -15318 2043 -15284 2059
rect -15318 2025 -15284 2043
rect -15318 1975 -15284 1987
rect -15318 1953 -15284 1975
rect -15318 1907 -15284 1915
rect -15318 1881 -15284 1907
rect -15222 2825 -15188 2851
rect -15222 2817 -15188 2825
rect -15222 2757 -15188 2779
rect -15222 2745 -15188 2757
rect -15222 2689 -15188 2707
rect -15222 2673 -15188 2689
rect -15222 2621 -15188 2635
rect -15222 2601 -15188 2621
rect -15222 2553 -15188 2563
rect -15222 2529 -15188 2553
rect -15222 2485 -15188 2491
rect -15222 2457 -15188 2485
rect -15222 2417 -15188 2419
rect -15222 2385 -15188 2417
rect -15222 2315 -15188 2347
rect -15222 2313 -15188 2315
rect -15222 2247 -15188 2275
rect -15222 2241 -15188 2247
rect -15222 2179 -15188 2203
rect -15222 2169 -15188 2179
rect -15222 2111 -15188 2131
rect -15222 2097 -15188 2111
rect -15222 2043 -15188 2059
rect -15222 2025 -15188 2043
rect -15222 1975 -15188 1987
rect -15222 1953 -15188 1975
rect -15222 1907 -15188 1915
rect -15222 1881 -15188 1907
rect -15126 2825 -15092 2851
rect -15126 2817 -15092 2825
rect -15126 2757 -15092 2779
rect -15126 2745 -15092 2757
rect -15126 2689 -15092 2707
rect -15126 2673 -15092 2689
rect -15126 2621 -15092 2635
rect -15126 2601 -15092 2621
rect -15126 2553 -15092 2563
rect -15126 2529 -15092 2553
rect -15126 2485 -15092 2491
rect -15126 2457 -15092 2485
rect -15126 2417 -15092 2419
rect -15126 2385 -15092 2417
rect -15126 2315 -15092 2347
rect -15126 2313 -15092 2315
rect -15126 2247 -15092 2275
rect -15126 2241 -15092 2247
rect -15126 2179 -15092 2203
rect -15126 2169 -15092 2179
rect -15126 2111 -15092 2131
rect -15126 2097 -15092 2111
rect -15126 2043 -15092 2059
rect -15126 2025 -15092 2043
rect -15126 1975 -15092 1987
rect -15126 1953 -15092 1975
rect -15126 1907 -15092 1915
rect -15126 1881 -15092 1907
rect -15030 2825 -14996 2851
rect -15030 2817 -14996 2825
rect -15030 2757 -14996 2779
rect -15030 2745 -14996 2757
rect -15030 2689 -14996 2707
rect -15030 2673 -14996 2689
rect -15030 2621 -14996 2635
rect -15030 2601 -14996 2621
rect -15030 2553 -14996 2563
rect -15030 2529 -14996 2553
rect -15030 2485 -14996 2491
rect -15030 2457 -14996 2485
rect -15030 2417 -14996 2419
rect -15030 2385 -14996 2417
rect -15030 2315 -14996 2347
rect -15030 2313 -14996 2315
rect -15030 2247 -14996 2275
rect -15030 2241 -14996 2247
rect -15030 2179 -14996 2203
rect -15030 2169 -14996 2179
rect -15030 2111 -14996 2131
rect -15030 2097 -14996 2111
rect -15030 2043 -14996 2059
rect -15030 2025 -14996 2043
rect -15030 1975 -14996 1987
rect -15030 1953 -14996 1975
rect -15030 1907 -14996 1915
rect -15030 1881 -14996 1907
rect -14934 2825 -14900 2851
rect -14934 2817 -14900 2825
rect -14934 2757 -14900 2779
rect -14934 2745 -14900 2757
rect -14934 2689 -14900 2707
rect -14934 2673 -14900 2689
rect -14934 2621 -14900 2635
rect -14934 2601 -14900 2621
rect -14934 2553 -14900 2563
rect -14934 2529 -14900 2553
rect -14934 2485 -14900 2491
rect -14934 2457 -14900 2485
rect -14934 2417 -14900 2419
rect -14934 2385 -14900 2417
rect -14934 2315 -14900 2347
rect -14934 2313 -14900 2315
rect -14934 2247 -14900 2275
rect -14934 2241 -14900 2247
rect -14934 2179 -14900 2203
rect -14934 2169 -14900 2179
rect -14934 2111 -14900 2131
rect -14934 2097 -14900 2111
rect -14934 2043 -14900 2059
rect -14934 2025 -14900 2043
rect -14934 1975 -14900 1987
rect -14934 1953 -14900 1975
rect -14934 1907 -14900 1915
rect -14934 1881 -14900 1907
rect -14838 2825 -14804 2851
rect -14838 2817 -14804 2825
rect -14838 2757 -14804 2779
rect -14838 2745 -14804 2757
rect -14838 2689 -14804 2707
rect -14838 2673 -14804 2689
rect -14838 2621 -14804 2635
rect -14838 2601 -14804 2621
rect -14838 2553 -14804 2563
rect -14838 2529 -14804 2553
rect -14838 2485 -14804 2491
rect -14838 2457 -14804 2485
rect -14838 2417 -14804 2419
rect -14838 2385 -14804 2417
rect -14838 2315 -14804 2347
rect -14838 2313 -14804 2315
rect -14838 2247 -14804 2275
rect -14838 2241 -14804 2247
rect -14838 2179 -14804 2203
rect -14838 2169 -14804 2179
rect -14838 2111 -14804 2131
rect -14838 2097 -14804 2111
rect -14838 2043 -14804 2059
rect -14838 2025 -14804 2043
rect -14838 1975 -14804 1987
rect -14838 1953 -14804 1975
rect -14838 1907 -14804 1915
rect -14838 1881 -14804 1907
rect -14742 2825 -14708 2851
rect -14742 2817 -14708 2825
rect -14742 2757 -14708 2779
rect -14742 2745 -14708 2757
rect -14742 2689 -14708 2707
rect -14742 2673 -14708 2689
rect -14742 2621 -14708 2635
rect -14742 2601 -14708 2621
rect -14742 2553 -14708 2563
rect -14742 2529 -14708 2553
rect -14742 2485 -14708 2491
rect -14742 2457 -14708 2485
rect -14742 2417 -14708 2419
rect -14742 2385 -14708 2417
rect -14742 2315 -14708 2347
rect -14742 2313 -14708 2315
rect -14742 2247 -14708 2275
rect -14742 2241 -14708 2247
rect -14742 2179 -14708 2203
rect -14742 2169 -14708 2179
rect -14742 2111 -14708 2131
rect -14742 2097 -14708 2111
rect -14742 2043 -14708 2059
rect -14742 2025 -14708 2043
rect -14742 1975 -14708 1987
rect -14742 1953 -14708 1975
rect -14742 1907 -14708 1915
rect -14742 1881 -14708 1907
rect -14514 2817 -14480 2843
rect -14514 2809 -14480 2817
rect -14514 2749 -14480 2771
rect -14514 2737 -14480 2749
rect -14514 2681 -14480 2699
rect -14514 2665 -14480 2681
rect -14514 2613 -14480 2627
rect -14514 2593 -14480 2613
rect -14514 2545 -14480 2555
rect -14514 2521 -14480 2545
rect -14514 2477 -14480 2483
rect -14514 2449 -14480 2477
rect -14514 2409 -14480 2411
rect -14514 2377 -14480 2409
rect -14514 2307 -14480 2339
rect -14514 2305 -14480 2307
rect -14514 2239 -14480 2267
rect -14514 2233 -14480 2239
rect -14514 2171 -14480 2195
rect -14514 2161 -14480 2171
rect -14514 2103 -14480 2123
rect -14514 2089 -14480 2103
rect -14514 2035 -14480 2051
rect -14514 2017 -14480 2035
rect -14514 1967 -14480 1979
rect -14514 1945 -14480 1967
rect -14514 1899 -14480 1907
rect -14514 1873 -14480 1899
rect -14418 2817 -14384 2843
rect -14418 2809 -14384 2817
rect -14418 2749 -14384 2771
rect -14418 2737 -14384 2749
rect -14418 2681 -14384 2699
rect -14418 2665 -14384 2681
rect -14418 2613 -14384 2627
rect -14418 2593 -14384 2613
rect -14418 2545 -14384 2555
rect -14418 2521 -14384 2545
rect -14418 2477 -14384 2483
rect -14418 2449 -14384 2477
rect -14418 2409 -14384 2411
rect -14418 2377 -14384 2409
rect -14418 2307 -14384 2339
rect -14418 2305 -14384 2307
rect -14418 2239 -14384 2267
rect -14418 2233 -14384 2239
rect -14418 2171 -14384 2195
rect -14418 2161 -14384 2171
rect -14418 2103 -14384 2123
rect -14418 2089 -14384 2103
rect -14418 2035 -14384 2051
rect -14418 2017 -14384 2035
rect -14418 1967 -14384 1979
rect -14418 1945 -14384 1967
rect -14418 1899 -14384 1907
rect -14418 1873 -14384 1899
rect -14322 2817 -14288 2843
rect -14322 2809 -14288 2817
rect -14322 2749 -14288 2771
rect -14322 2737 -14288 2749
rect -14322 2681 -14288 2699
rect -14322 2665 -14288 2681
rect -14322 2613 -14288 2627
rect -14322 2593 -14288 2613
rect -14322 2545 -14288 2555
rect -14322 2521 -14288 2545
rect -14322 2477 -14288 2483
rect -14322 2449 -14288 2477
rect -14322 2409 -14288 2411
rect -14322 2377 -14288 2409
rect -14322 2307 -14288 2339
rect -14322 2305 -14288 2307
rect -14322 2239 -14288 2267
rect -14322 2233 -14288 2239
rect -14322 2171 -14288 2195
rect -14322 2161 -14288 2171
rect -14322 2103 -14288 2123
rect -14322 2089 -14288 2103
rect -14322 2035 -14288 2051
rect -14322 2017 -14288 2035
rect -14322 1967 -14288 1979
rect -14322 1945 -14288 1967
rect -14322 1899 -14288 1907
rect -14322 1873 -14288 1899
rect -14226 2817 -14192 2843
rect -14226 2809 -14192 2817
rect -14226 2749 -14192 2771
rect -14226 2737 -14192 2749
rect -14226 2681 -14192 2699
rect -14226 2665 -14192 2681
rect -14226 2613 -14192 2627
rect -14226 2593 -14192 2613
rect -14226 2545 -14192 2555
rect -14226 2521 -14192 2545
rect -14226 2477 -14192 2483
rect -14226 2449 -14192 2477
rect -14226 2409 -14192 2411
rect -14226 2377 -14192 2409
rect -14226 2307 -14192 2339
rect -14226 2305 -14192 2307
rect -14226 2239 -14192 2267
rect -14226 2233 -14192 2239
rect -14226 2171 -14192 2195
rect -14226 2161 -14192 2171
rect -14226 2103 -14192 2123
rect -14226 2089 -14192 2103
rect -14226 2035 -14192 2051
rect -14226 2017 -14192 2035
rect -14226 1967 -14192 1979
rect -14226 1945 -14192 1967
rect -14226 1899 -14192 1907
rect -14226 1873 -14192 1899
rect -14130 2817 -14096 2843
rect -14130 2809 -14096 2817
rect -14130 2749 -14096 2771
rect -14130 2737 -14096 2749
rect -14130 2681 -14096 2699
rect -14130 2665 -14096 2681
rect -14130 2613 -14096 2627
rect -14130 2593 -14096 2613
rect -14130 2545 -14096 2555
rect -14130 2521 -14096 2545
rect -14130 2477 -14096 2483
rect -14130 2449 -14096 2477
rect -14130 2409 -14096 2411
rect -14130 2377 -14096 2409
rect -14130 2307 -14096 2339
rect -14130 2305 -14096 2307
rect -14130 2239 -14096 2267
rect -14130 2233 -14096 2239
rect -14130 2171 -14096 2195
rect -14130 2161 -14096 2171
rect -14130 2103 -14096 2123
rect -14130 2089 -14096 2103
rect -14130 2035 -14096 2051
rect -14130 2017 -14096 2035
rect -14130 1967 -14096 1979
rect -14130 1945 -14096 1967
rect -14130 1899 -14096 1907
rect -14130 1873 -14096 1899
rect -14034 2817 -14000 2843
rect -14034 2809 -14000 2817
rect -14034 2749 -14000 2771
rect -14034 2737 -14000 2749
rect -14034 2681 -14000 2699
rect -14034 2665 -14000 2681
rect -14034 2613 -14000 2627
rect -14034 2593 -14000 2613
rect -14034 2545 -14000 2555
rect -14034 2521 -14000 2545
rect -14034 2477 -14000 2483
rect -14034 2449 -14000 2477
rect -14034 2409 -14000 2411
rect -14034 2377 -14000 2409
rect -14034 2307 -14000 2339
rect -14034 2305 -14000 2307
rect -14034 2239 -14000 2267
rect -14034 2233 -14000 2239
rect -14034 2171 -14000 2195
rect -14034 2161 -14000 2171
rect -14034 2103 -14000 2123
rect -14034 2089 -14000 2103
rect -14034 2035 -14000 2051
rect -14034 2017 -14000 2035
rect -14034 1967 -14000 1979
rect -14034 1945 -14000 1967
rect -14034 1899 -14000 1907
rect -14034 1873 -14000 1899
rect -13938 2817 -13904 2843
rect -13938 2809 -13904 2817
rect -13938 2749 -13904 2771
rect -13938 2737 -13904 2749
rect -13938 2681 -13904 2699
rect -13938 2665 -13904 2681
rect -13938 2613 -13904 2627
rect -13938 2593 -13904 2613
rect -13938 2545 -13904 2555
rect -13938 2521 -13904 2545
rect -13938 2477 -13904 2483
rect -13938 2449 -13904 2477
rect -13938 2409 -13904 2411
rect -13938 2377 -13904 2409
rect -13938 2307 -13904 2339
rect -13938 2305 -13904 2307
rect -13938 2239 -13904 2267
rect -13938 2233 -13904 2239
rect -13938 2171 -13904 2195
rect -13938 2161 -13904 2171
rect -13938 2103 -13904 2123
rect -13938 2089 -13904 2103
rect -13938 2035 -13904 2051
rect -13938 2017 -13904 2035
rect -13938 1967 -13904 1979
rect -13938 1945 -13904 1967
rect -13938 1899 -13904 1907
rect -13938 1873 -13904 1899
rect -13842 2817 -13808 2843
rect -13842 2809 -13808 2817
rect -13842 2749 -13808 2771
rect -13842 2737 -13808 2749
rect -13842 2681 -13808 2699
rect -13842 2665 -13808 2681
rect -13842 2613 -13808 2627
rect -13842 2593 -13808 2613
rect -13842 2545 -13808 2555
rect -13842 2521 -13808 2545
rect -13842 2477 -13808 2483
rect -13842 2449 -13808 2477
rect -13842 2409 -13808 2411
rect -13842 2377 -13808 2409
rect -13842 2307 -13808 2339
rect -13842 2305 -13808 2307
rect -13842 2239 -13808 2267
rect -13842 2233 -13808 2239
rect -13842 2171 -13808 2195
rect -13842 2161 -13808 2171
rect -13842 2103 -13808 2123
rect -13842 2089 -13808 2103
rect -13842 2035 -13808 2051
rect -13842 2017 -13808 2035
rect -13842 1967 -13808 1979
rect -13842 1945 -13808 1967
rect -13842 1899 -13808 1907
rect -13842 1873 -13808 1899
rect -13746 2817 -13712 2843
rect -13746 2809 -13712 2817
rect -13746 2749 -13712 2771
rect -13746 2737 -13712 2749
rect -13746 2681 -13712 2699
rect -13746 2665 -13712 2681
rect -13746 2613 -13712 2627
rect -13746 2593 -13712 2613
rect -13746 2545 -13712 2555
rect -13746 2521 -13712 2545
rect -13746 2477 -13712 2483
rect -13746 2449 -13712 2477
rect -13746 2409 -13712 2411
rect -13746 2377 -13712 2409
rect -13746 2307 -13712 2339
rect -13746 2305 -13712 2307
rect -13746 2239 -13712 2267
rect -13746 2233 -13712 2239
rect -13746 2171 -13712 2195
rect -13746 2161 -13712 2171
rect -13746 2103 -13712 2123
rect -13746 2089 -13712 2103
rect -13746 2035 -13712 2051
rect -13746 2017 -13712 2035
rect -13746 1967 -13712 1979
rect -13746 1945 -13712 1967
rect -13746 1899 -13712 1907
rect -13746 1873 -13712 1899
rect -13650 2817 -13616 2843
rect -13650 2809 -13616 2817
rect -13650 2749 -13616 2771
rect -13650 2737 -13616 2749
rect -13650 2681 -13616 2699
rect -13650 2665 -13616 2681
rect -13650 2613 -13616 2627
rect -13650 2593 -13616 2613
rect -13650 2545 -13616 2555
rect -13650 2521 -13616 2545
rect -13650 2477 -13616 2483
rect -13650 2449 -13616 2477
rect -13650 2409 -13616 2411
rect -13650 2377 -13616 2409
rect -13650 2307 -13616 2339
rect -13650 2305 -13616 2307
rect -13650 2239 -13616 2267
rect -13650 2233 -13616 2239
rect -13650 2171 -13616 2195
rect -13650 2161 -13616 2171
rect -13650 2103 -13616 2123
rect -13650 2089 -13616 2103
rect -13650 2035 -13616 2051
rect -13650 2017 -13616 2035
rect -13650 1967 -13616 1979
rect -13650 1945 -13616 1967
rect -13650 1899 -13616 1907
rect -13650 1873 -13616 1899
rect -13554 2817 -13520 2843
rect -13554 2809 -13520 2817
rect -13554 2749 -13520 2771
rect -13554 2737 -13520 2749
rect -13554 2681 -13520 2699
rect -13554 2665 -13520 2681
rect -13554 2613 -13520 2627
rect -13554 2593 -13520 2613
rect -13554 2545 -13520 2555
rect -13554 2521 -13520 2545
rect -13554 2477 -13520 2483
rect -13554 2449 -13520 2477
rect -13554 2409 -13520 2411
rect -13554 2377 -13520 2409
rect -13554 2307 -13520 2339
rect -13554 2305 -13520 2307
rect -13554 2239 -13520 2267
rect -13554 2233 -13520 2239
rect -13554 2171 -13520 2195
rect -13554 2161 -13520 2171
rect -13554 2103 -13520 2123
rect -13554 2089 -13520 2103
rect -13554 2035 -13520 2051
rect -13554 2017 -13520 2035
rect -13554 1967 -13520 1979
rect -13554 1945 -13520 1967
rect -13554 1899 -13520 1907
rect -13554 1873 -13520 1899
rect -13458 2817 -13424 2843
rect -13458 2809 -13424 2817
rect -13458 2749 -13424 2771
rect -13458 2737 -13424 2749
rect -13458 2681 -13424 2699
rect -13458 2665 -13424 2681
rect -13458 2613 -13424 2627
rect -13458 2593 -13424 2613
rect -13458 2545 -13424 2555
rect -13458 2521 -13424 2545
rect -13458 2477 -13424 2483
rect -13458 2449 -13424 2477
rect -13458 2409 -13424 2411
rect -13458 2377 -13424 2409
rect -13458 2307 -13424 2339
rect -13458 2305 -13424 2307
rect -13458 2239 -13424 2267
rect -13458 2233 -13424 2239
rect -13458 2171 -13424 2195
rect -13458 2161 -13424 2171
rect -13458 2103 -13424 2123
rect -13458 2089 -13424 2103
rect -13458 2035 -13424 2051
rect -13458 2017 -13424 2035
rect -13458 1967 -13424 1979
rect -13458 1945 -13424 1967
rect -13458 1899 -13424 1907
rect -13458 1873 -13424 1899
rect -13362 2817 -13328 2843
rect -13362 2809 -13328 2817
rect -13362 2749 -13328 2771
rect -13362 2737 -13328 2749
rect -13362 2681 -13328 2699
rect -13362 2665 -13328 2681
rect -13362 2613 -13328 2627
rect -13362 2593 -13328 2613
rect -13362 2545 -13328 2555
rect -13362 2521 -13328 2545
rect -13362 2477 -13328 2483
rect -13362 2449 -13328 2477
rect -13362 2409 -13328 2411
rect -13362 2377 -13328 2409
rect -13362 2307 -13328 2339
rect -13362 2305 -13328 2307
rect -13362 2239 -13328 2267
rect -13362 2233 -13328 2239
rect -13362 2171 -13328 2195
rect -13362 2161 -13328 2171
rect -13362 2103 -13328 2123
rect -13362 2089 -13328 2103
rect -13362 2035 -13328 2051
rect -13362 2017 -13328 2035
rect -13362 1967 -13328 1979
rect -13362 1945 -13328 1967
rect -13362 1899 -13328 1907
rect -13362 1873 -13328 1899
rect -13266 2817 -13232 2843
rect -13266 2809 -13232 2817
rect -13266 2749 -13232 2771
rect -13266 2737 -13232 2749
rect -13266 2681 -13232 2699
rect -13266 2665 -13232 2681
rect -13266 2613 -13232 2627
rect -13266 2593 -13232 2613
rect -13266 2545 -13232 2555
rect -13266 2521 -13232 2545
rect -13266 2477 -13232 2483
rect -13266 2449 -13232 2477
rect -13266 2409 -13232 2411
rect -13266 2377 -13232 2409
rect -13266 2307 -13232 2339
rect -13266 2305 -13232 2307
rect -13266 2239 -13232 2267
rect -13266 2233 -13232 2239
rect -13266 2171 -13232 2195
rect -13266 2161 -13232 2171
rect -13266 2103 -13232 2123
rect -13266 2089 -13232 2103
rect -13266 2035 -13232 2051
rect -13266 2017 -13232 2035
rect -13266 1967 -13232 1979
rect -13266 1945 -13232 1967
rect -13266 1899 -13232 1907
rect -13266 1873 -13232 1899
rect -6270 4423 -6236 4449
rect -6270 4415 -6236 4423
rect -6270 4355 -6236 4377
rect -6270 4343 -6236 4355
rect -6270 4287 -6236 4305
rect -6270 4271 -6236 4287
rect -6270 4219 -6236 4233
rect -6270 4199 -6236 4219
rect -6270 4151 -6236 4161
rect -6270 4127 -6236 4151
rect -6270 4083 -6236 4089
rect -6270 4055 -6236 4083
rect -6270 4015 -6236 4017
rect -6270 3983 -6236 4015
rect -6270 3913 -6236 3945
rect -6270 3911 -6236 3913
rect -6270 3845 -6236 3873
rect -6270 3839 -6236 3845
rect -6270 3777 -6236 3801
rect -6270 3767 -6236 3777
rect -6270 3709 -6236 3729
rect -6270 3695 -6236 3709
rect -6270 3641 -6236 3657
rect -6270 3623 -6236 3641
rect -6270 3573 -6236 3585
rect -6270 3551 -6236 3573
rect -6270 3505 -6236 3513
rect -6270 3479 -6236 3505
rect -6174 4423 -6140 4449
rect -6174 4415 -6140 4423
rect -6174 4355 -6140 4377
rect -6174 4343 -6140 4355
rect -6174 4287 -6140 4305
rect -6174 4271 -6140 4287
rect -6174 4219 -6140 4233
rect -6174 4199 -6140 4219
rect -6174 4151 -6140 4161
rect -6174 4127 -6140 4151
rect -6174 4083 -6140 4089
rect -6174 4055 -6140 4083
rect -6174 4015 -6140 4017
rect -6174 3983 -6140 4015
rect -6174 3913 -6140 3945
rect -6174 3911 -6140 3913
rect -6174 3845 -6140 3873
rect -6174 3839 -6140 3845
rect -6174 3777 -6140 3801
rect -6174 3767 -6140 3777
rect -6174 3709 -6140 3729
rect -6174 3695 -6140 3709
rect -6174 3641 -6140 3657
rect -6174 3623 -6140 3641
rect -6174 3573 -6140 3585
rect -6174 3551 -6140 3573
rect -6174 3505 -6140 3513
rect -6174 3479 -6140 3505
rect -6078 4423 -6044 4449
rect -6078 4415 -6044 4423
rect -6078 4355 -6044 4377
rect -6078 4343 -6044 4355
rect -6078 4287 -6044 4305
rect -6078 4271 -6044 4287
rect -6078 4219 -6044 4233
rect -6078 4199 -6044 4219
rect -6078 4151 -6044 4161
rect -6078 4127 -6044 4151
rect -6078 4083 -6044 4089
rect -6078 4055 -6044 4083
rect -6078 4015 -6044 4017
rect -6078 3983 -6044 4015
rect -6078 3913 -6044 3945
rect -6078 3911 -6044 3913
rect -6078 3845 -6044 3873
rect -6078 3839 -6044 3845
rect -6078 3777 -6044 3801
rect -6078 3767 -6044 3777
rect -6078 3709 -6044 3729
rect -6078 3695 -6044 3709
rect -6078 3641 -6044 3657
rect -6078 3623 -6044 3641
rect -6078 3573 -6044 3585
rect -6078 3551 -6044 3573
rect -6078 3505 -6044 3513
rect -6078 3479 -6044 3505
rect -5982 4423 -5948 4449
rect -5982 4415 -5948 4423
rect -5982 4355 -5948 4377
rect -5982 4343 -5948 4355
rect -5982 4287 -5948 4305
rect -5982 4271 -5948 4287
rect -5982 4219 -5948 4233
rect -5982 4199 -5948 4219
rect -5982 4151 -5948 4161
rect -5982 4127 -5948 4151
rect -5982 4083 -5948 4089
rect -5982 4055 -5948 4083
rect -5982 4015 -5948 4017
rect -5982 3983 -5948 4015
rect -5982 3913 -5948 3945
rect -5982 3911 -5948 3913
rect -5982 3845 -5948 3873
rect -5982 3839 -5948 3845
rect -5982 3777 -5948 3801
rect -5982 3767 -5948 3777
rect -5982 3709 -5948 3729
rect -5982 3695 -5948 3709
rect -5982 3641 -5948 3657
rect -5982 3623 -5948 3641
rect -5982 3573 -5948 3585
rect -5982 3551 -5948 3573
rect -5982 3505 -5948 3513
rect -5982 3479 -5948 3505
rect -5886 4423 -5852 4449
rect -5886 4415 -5852 4423
rect -5886 4355 -5852 4377
rect -5886 4343 -5852 4355
rect -5886 4287 -5852 4305
rect -5886 4271 -5852 4287
rect -5886 4219 -5852 4233
rect -5886 4199 -5852 4219
rect -5886 4151 -5852 4161
rect -5886 4127 -5852 4151
rect -5886 4083 -5852 4089
rect -5886 4055 -5852 4083
rect -5886 4015 -5852 4017
rect -5886 3983 -5852 4015
rect -5886 3913 -5852 3945
rect -5886 3911 -5852 3913
rect -5886 3845 -5852 3873
rect -5886 3839 -5852 3845
rect -5886 3777 -5852 3801
rect -5886 3767 -5852 3777
rect -5886 3709 -5852 3729
rect -5886 3695 -5852 3709
rect -5886 3641 -5852 3657
rect -5886 3623 -5852 3641
rect -5886 3573 -5852 3585
rect -5886 3551 -5852 3573
rect -5886 3505 -5852 3513
rect -5886 3479 -5852 3505
rect -5790 4423 -5756 4449
rect -5790 4415 -5756 4423
rect -5790 4355 -5756 4377
rect -5790 4343 -5756 4355
rect -5790 4287 -5756 4305
rect -5790 4271 -5756 4287
rect -5790 4219 -5756 4233
rect -5790 4199 -5756 4219
rect -5790 4151 -5756 4161
rect -5790 4127 -5756 4151
rect -5790 4083 -5756 4089
rect -5790 4055 -5756 4083
rect -5790 4015 -5756 4017
rect -5790 3983 -5756 4015
rect -5790 3913 -5756 3945
rect -5790 3911 -5756 3913
rect -5790 3845 -5756 3873
rect -5790 3839 -5756 3845
rect -5790 3777 -5756 3801
rect -5790 3767 -5756 3777
rect -5790 3709 -5756 3729
rect -5790 3695 -5756 3709
rect -5790 3641 -5756 3657
rect -5790 3623 -5756 3641
rect -5790 3573 -5756 3585
rect -5790 3551 -5756 3573
rect -5790 3505 -5756 3513
rect -5790 3479 -5756 3505
rect -5694 4423 -5660 4449
rect -5694 4415 -5660 4423
rect -5694 4355 -5660 4377
rect -5694 4343 -5660 4355
rect -5694 4287 -5660 4305
rect -5694 4271 -5660 4287
rect -5694 4219 -5660 4233
rect -5694 4199 -5660 4219
rect -5694 4151 -5660 4161
rect -5694 4127 -5660 4151
rect -5694 4083 -5660 4089
rect -5694 4055 -5660 4083
rect -5694 4015 -5660 4017
rect -5694 3983 -5660 4015
rect -5694 3913 -5660 3945
rect -5694 3911 -5660 3913
rect -5694 3845 -5660 3873
rect -5694 3839 -5660 3845
rect -5694 3777 -5660 3801
rect -5694 3767 -5660 3777
rect -5694 3709 -5660 3729
rect -5694 3695 -5660 3709
rect -5694 3641 -5660 3657
rect -5694 3623 -5660 3641
rect -5694 3573 -5660 3585
rect -5694 3551 -5660 3573
rect -5694 3505 -5660 3513
rect -5694 3479 -5660 3505
rect -5598 4423 -5564 4449
rect -5598 4415 -5564 4423
rect -5598 4355 -5564 4377
rect -5598 4343 -5564 4355
rect -5598 4287 -5564 4305
rect -5598 4271 -5564 4287
rect -5598 4219 -5564 4233
rect -5598 4199 -5564 4219
rect -5598 4151 -5564 4161
rect -5598 4127 -5564 4151
rect -5598 4083 -5564 4089
rect -5598 4055 -5564 4083
rect -5598 4015 -5564 4017
rect -5598 3983 -5564 4015
rect -5598 3913 -5564 3945
rect -5598 3911 -5564 3913
rect -5598 3845 -5564 3873
rect -5598 3839 -5564 3845
rect -5598 3777 -5564 3801
rect -5598 3767 -5564 3777
rect -5598 3709 -5564 3729
rect -5598 3695 -5564 3709
rect -5598 3641 -5564 3657
rect -5598 3623 -5564 3641
rect -5598 3573 -5564 3585
rect -5598 3551 -5564 3573
rect -5598 3505 -5564 3513
rect -5598 3479 -5564 3505
rect -5502 4423 -5468 4449
rect -5502 4415 -5468 4423
rect -5502 4355 -5468 4377
rect -5502 4343 -5468 4355
rect -5502 4287 -5468 4305
rect -5502 4271 -5468 4287
rect -5502 4219 -5468 4233
rect -5502 4199 -5468 4219
rect -5502 4151 -5468 4161
rect -5502 4127 -5468 4151
rect -5502 4083 -5468 4089
rect -5502 4055 -5468 4083
rect -5502 4015 -5468 4017
rect -5502 3983 -5468 4015
rect -5502 3913 -5468 3945
rect -5502 3911 -5468 3913
rect -5502 3845 -5468 3873
rect -5502 3839 -5468 3845
rect -5502 3777 -5468 3801
rect -5502 3767 -5468 3777
rect -5502 3709 -5468 3729
rect -5502 3695 -5468 3709
rect -5502 3641 -5468 3657
rect -5502 3623 -5468 3641
rect -5502 3573 -5468 3585
rect -5502 3551 -5468 3573
rect -5502 3505 -5468 3513
rect -5502 3479 -5468 3505
rect -5294 4425 -5260 4451
rect -5294 4417 -5260 4425
rect -5294 4357 -5260 4379
rect -5294 4345 -5260 4357
rect -5294 4289 -5260 4307
rect -5294 4273 -5260 4289
rect -5294 4221 -5260 4235
rect -5294 4201 -5260 4221
rect -5294 4153 -5260 4163
rect -5294 4129 -5260 4153
rect -5294 4085 -5260 4091
rect -5294 4057 -5260 4085
rect -5294 4017 -5260 4019
rect -5294 3985 -5260 4017
rect -5294 3915 -5260 3947
rect -5294 3913 -5260 3915
rect -5294 3847 -5260 3875
rect -5294 3841 -5260 3847
rect -5294 3779 -5260 3803
rect -5294 3769 -5260 3779
rect -5294 3711 -5260 3731
rect -5294 3697 -5260 3711
rect -5294 3643 -5260 3659
rect -5294 3625 -5260 3643
rect -5294 3575 -5260 3587
rect -5294 3553 -5260 3575
rect -5294 3507 -5260 3515
rect -5294 3481 -5260 3507
rect -5198 4425 -5164 4451
rect -5198 4417 -5164 4425
rect -5198 4357 -5164 4379
rect -5198 4345 -5164 4357
rect -5198 4289 -5164 4307
rect -5198 4273 -5164 4289
rect -5198 4221 -5164 4235
rect -5198 4201 -5164 4221
rect -5198 4153 -5164 4163
rect -5198 4129 -5164 4153
rect -5198 4085 -5164 4091
rect -5198 4057 -5164 4085
rect -5198 4017 -5164 4019
rect -5198 3985 -5164 4017
rect -5198 3915 -5164 3947
rect -5198 3913 -5164 3915
rect -5198 3847 -5164 3875
rect -5198 3841 -5164 3847
rect -5198 3779 -5164 3803
rect -5198 3769 -5164 3779
rect -5198 3711 -5164 3731
rect -5198 3697 -5164 3711
rect -5198 3643 -5164 3659
rect -5198 3625 -5164 3643
rect -5198 3575 -5164 3587
rect -5198 3553 -5164 3575
rect -5198 3507 -5164 3515
rect -5198 3481 -5164 3507
rect -5102 4425 -5068 4451
rect -5102 4417 -5068 4425
rect -5102 4357 -5068 4379
rect -5102 4345 -5068 4357
rect -5102 4289 -5068 4307
rect -5102 4273 -5068 4289
rect -5102 4221 -5068 4235
rect -5102 4201 -5068 4221
rect -5102 4153 -5068 4163
rect -5102 4129 -5068 4153
rect -5102 4085 -5068 4091
rect -5102 4057 -5068 4085
rect -5102 4017 -5068 4019
rect -5102 3985 -5068 4017
rect -5102 3915 -5068 3947
rect -5102 3913 -5068 3915
rect -5102 3847 -5068 3875
rect -5102 3841 -5068 3847
rect -5102 3779 -5068 3803
rect -5102 3769 -5068 3779
rect -5102 3711 -5068 3731
rect -5102 3697 -5068 3711
rect -5102 3643 -5068 3659
rect -5102 3625 -5068 3643
rect -5102 3575 -5068 3587
rect -5102 3553 -5068 3575
rect -5102 3507 -5068 3515
rect -5102 3481 -5068 3507
rect -5006 4425 -4972 4451
rect -5006 4417 -4972 4425
rect -5006 4357 -4972 4379
rect -5006 4345 -4972 4357
rect -5006 4289 -4972 4307
rect -5006 4273 -4972 4289
rect -5006 4221 -4972 4235
rect -5006 4201 -4972 4221
rect -5006 4153 -4972 4163
rect -5006 4129 -4972 4153
rect -5006 4085 -4972 4091
rect -5006 4057 -4972 4085
rect -5006 4017 -4972 4019
rect -5006 3985 -4972 4017
rect -5006 3915 -4972 3947
rect -5006 3913 -4972 3915
rect -5006 3847 -4972 3875
rect -5006 3841 -4972 3847
rect -5006 3779 -4972 3803
rect -5006 3769 -4972 3779
rect -5006 3711 -4972 3731
rect -5006 3697 -4972 3711
rect -5006 3643 -4972 3659
rect -5006 3625 -4972 3643
rect -5006 3575 -4972 3587
rect -5006 3553 -4972 3575
rect -5006 3507 -4972 3515
rect -5006 3481 -4972 3507
rect -4910 4425 -4876 4451
rect -4910 4417 -4876 4425
rect -4910 4357 -4876 4379
rect -4910 4345 -4876 4357
rect -4910 4289 -4876 4307
rect -4910 4273 -4876 4289
rect -4910 4221 -4876 4235
rect -4910 4201 -4876 4221
rect -4910 4153 -4876 4163
rect -4910 4129 -4876 4153
rect -4910 4085 -4876 4091
rect -4910 4057 -4876 4085
rect -4910 4017 -4876 4019
rect -4910 3985 -4876 4017
rect -4910 3915 -4876 3947
rect -4910 3913 -4876 3915
rect -4910 3847 -4876 3875
rect -4910 3841 -4876 3847
rect -4910 3779 -4876 3803
rect -4910 3769 -4876 3779
rect -4910 3711 -4876 3731
rect -4910 3697 -4876 3711
rect -4910 3643 -4876 3659
rect -4910 3625 -4876 3643
rect -4910 3575 -4876 3587
rect -4910 3553 -4876 3575
rect -4910 3507 -4876 3515
rect -4910 3481 -4876 3507
rect -4814 4425 -4780 4451
rect -4814 4417 -4780 4425
rect -4814 4357 -4780 4379
rect -4814 4345 -4780 4357
rect -4814 4289 -4780 4307
rect -4814 4273 -4780 4289
rect -4814 4221 -4780 4235
rect -4814 4201 -4780 4221
rect -4814 4153 -4780 4163
rect -4814 4129 -4780 4153
rect -4814 4085 -4780 4091
rect -4814 4057 -4780 4085
rect -4814 4017 -4780 4019
rect -4814 3985 -4780 4017
rect -4814 3915 -4780 3947
rect 1484 4535 1518 4563
rect 1484 4495 1518 4497
rect 1484 4463 1518 4495
rect 1484 4393 1518 4425
rect 1484 4391 1518 4393
rect 1484 4325 1518 4353
rect 1484 4319 1518 4325
rect 1484 4257 1518 4281
rect 1484 4247 1518 4257
rect 1484 4189 1518 4209
rect 1484 4175 1518 4189
rect 1484 4121 1518 4137
rect 1484 4103 1518 4121
rect 1484 4053 1518 4065
rect 1484 4031 1518 4053
rect 1484 3985 1518 3993
rect 1484 3959 1518 3985
rect 1580 4903 1614 4929
rect 1580 4895 1614 4903
rect 1580 4835 1614 4857
rect 1580 4823 1614 4835
rect 1580 4767 1614 4785
rect 1580 4751 1614 4767
rect 1580 4699 1614 4713
rect 1580 4679 1614 4699
rect 1580 4631 1614 4641
rect 1580 4607 1614 4631
rect 1580 4563 1614 4569
rect 1580 4535 1614 4563
rect 1580 4495 1614 4497
rect 1580 4463 1614 4495
rect 1580 4393 1614 4425
rect 1580 4391 1614 4393
rect 1580 4325 1614 4353
rect 1580 4319 1614 4325
rect 1580 4257 1614 4281
rect 1580 4247 1614 4257
rect 1580 4189 1614 4209
rect 1580 4175 1614 4189
rect 1580 4121 1614 4137
rect 1580 4103 1614 4121
rect 1580 4053 1614 4065
rect 1580 4031 1614 4053
rect 1580 3985 1614 3993
rect 1580 3959 1614 3985
rect -4814 3913 -4780 3915
rect -4814 3847 -4780 3875
rect 1676 4903 1710 4929
rect 1676 4895 1710 4903
rect 1676 4835 1710 4857
rect 1676 4823 1710 4835
rect 1676 4767 1710 4785
rect 1676 4751 1710 4767
rect 1676 4699 1710 4713
rect 1676 4679 1710 4699
rect 1676 4631 1710 4641
rect 1676 4607 1710 4631
rect 1676 4563 1710 4569
rect 1676 4535 1710 4563
rect 1676 4495 1710 4497
rect 1676 4463 1710 4495
rect 1676 4393 1710 4425
rect 1676 4391 1710 4393
rect 1676 4325 1710 4353
rect 1676 4319 1710 4325
rect 1676 4257 1710 4281
rect 1676 4247 1710 4257
rect 1676 4189 1710 4209
rect 1676 4175 1710 4189
rect 1676 4121 1710 4137
rect 1676 4103 1710 4121
rect 1676 4053 1710 4065
rect 1676 4031 1710 4053
rect 1676 3985 1710 3993
rect 1676 3959 1710 3985
rect 1772 4903 1806 4929
rect 1772 4895 1806 4903
rect 1772 4835 1806 4857
rect 1772 4823 1806 4835
rect 1772 4767 1806 4785
rect 1772 4751 1806 4767
rect 1772 4699 1806 4713
rect 1772 4679 1806 4699
rect 1772 4631 1806 4641
rect 1772 4607 1806 4631
rect 1772 4563 1806 4569
rect 1772 4535 1806 4563
rect 1772 4495 1806 4497
rect 1772 4463 1806 4495
rect 1772 4393 1806 4425
rect 1772 4391 1806 4393
rect 1772 4325 1806 4353
rect 1772 4319 1806 4325
rect 1772 4257 1806 4281
rect 1772 4247 1806 4257
rect 1772 4189 1806 4209
rect 1772 4175 1806 4189
rect 1772 4121 1806 4137
rect 1772 4103 1806 4121
rect 1772 4053 1806 4065
rect 1772 4031 1806 4053
rect 1772 3985 1806 3993
rect 1772 3959 1806 3985
rect 13810 5046 13844 5080
rect 1868 4903 1902 4929
rect 1868 4895 1902 4903
rect 1868 4835 1902 4857
rect 1868 4823 1902 4835
rect 1868 4767 1902 4785
rect 1868 4751 1902 4767
rect 1868 4699 1902 4713
rect 1868 4679 1902 4699
rect 1868 4631 1902 4641
rect 1868 4607 1902 4631
rect 1868 4563 1902 4569
rect 1868 4535 1902 4563
rect 1868 4495 1902 4497
rect 1868 4463 1902 4495
rect 1868 4393 1902 4425
rect 1868 4391 1902 4393
rect 1868 4325 1902 4353
rect 1868 4319 1902 4325
rect 1868 4257 1902 4281
rect 1868 4247 1902 4257
rect 1868 4189 1902 4209
rect 1868 4175 1902 4189
rect 1868 4121 1902 4137
rect 1868 4103 1902 4121
rect 1868 4053 1902 4065
rect 1868 4031 1902 4053
rect 1868 3985 1902 3993
rect 1868 3959 1902 3985
rect 4440 4887 4474 4913
rect 4440 4879 4474 4887
rect 4440 4819 4474 4841
rect 4440 4807 4474 4819
rect 4440 4751 4474 4769
rect 4440 4735 4474 4751
rect 4440 4683 4474 4697
rect 4440 4663 4474 4683
rect 4440 4615 4474 4625
rect 4440 4591 4474 4615
rect 4440 4547 4474 4553
rect 4440 4519 4474 4547
rect 4440 4479 4474 4481
rect 4440 4447 4474 4479
rect 4440 4377 4474 4409
rect 4440 4375 4474 4377
rect 4440 4309 4474 4337
rect 4440 4303 4474 4309
rect 4440 4241 4474 4265
rect 4440 4231 4474 4241
rect 4440 4173 4474 4193
rect 4440 4159 4474 4173
rect 4440 4105 4474 4121
rect 4440 4087 4474 4105
rect 4440 4037 4474 4049
rect 4440 4015 4474 4037
rect 4440 3969 4474 3977
rect 4440 3943 4474 3969
rect 4536 4887 4570 4913
rect 4536 4879 4570 4887
rect 4536 4819 4570 4841
rect 4536 4807 4570 4819
rect 4536 4751 4570 4769
rect 4536 4735 4570 4751
rect 4536 4683 4570 4697
rect 4536 4663 4570 4683
rect 4536 4615 4570 4625
rect 4536 4591 4570 4615
rect 4536 4547 4570 4553
rect 4536 4519 4570 4547
rect 4536 4479 4570 4481
rect 4536 4447 4570 4479
rect 4536 4377 4570 4409
rect 4536 4375 4570 4377
rect 4536 4309 4570 4337
rect 4536 4303 4570 4309
rect 4536 4241 4570 4265
rect 4536 4231 4570 4241
rect 4536 4173 4570 4193
rect 4536 4159 4570 4173
rect 4536 4105 4570 4121
rect 4536 4087 4570 4105
rect 4536 4037 4570 4049
rect 4536 4015 4570 4037
rect 4536 3969 4570 3977
rect 4536 3943 4570 3969
rect 4632 4887 4666 4913
rect 4632 4879 4666 4887
rect 4632 4819 4666 4841
rect 4632 4807 4666 4819
rect 4632 4751 4666 4769
rect 4632 4735 4666 4751
rect 4632 4683 4666 4697
rect 4632 4663 4666 4683
rect 4632 4615 4666 4625
rect 4632 4591 4666 4615
rect 4632 4547 4666 4553
rect 4632 4519 4666 4547
rect 4632 4479 4666 4481
rect 4632 4447 4666 4479
rect 4632 4377 4666 4409
rect 4632 4375 4666 4377
rect 4632 4309 4666 4337
rect 4632 4303 4666 4309
rect 4632 4241 4666 4265
rect 4632 4231 4666 4241
rect 4632 4173 4666 4193
rect 4632 4159 4666 4173
rect 4632 4105 4666 4121
rect 4632 4087 4666 4105
rect 4632 4037 4666 4049
rect 4632 4015 4666 4037
rect 4632 3969 4666 3977
rect 4632 3943 4666 3969
rect 4728 4887 4762 4913
rect 4728 4879 4762 4887
rect 4728 4819 4762 4841
rect 4728 4807 4762 4819
rect 4728 4751 4762 4769
rect 4728 4735 4762 4751
rect 4728 4683 4762 4697
rect 4728 4663 4762 4683
rect 4728 4615 4762 4625
rect 4728 4591 4762 4615
rect 4728 4547 4762 4553
rect 4728 4519 4762 4547
rect 4728 4479 4762 4481
rect 4728 4447 4762 4479
rect 4728 4377 4762 4409
rect 4728 4375 4762 4377
rect 4728 4309 4762 4337
rect 4728 4303 4762 4309
rect 4728 4241 4762 4265
rect 4728 4231 4762 4241
rect 4728 4173 4762 4193
rect 4728 4159 4762 4173
rect 4728 4105 4762 4121
rect 4728 4087 4762 4105
rect 4728 4037 4762 4049
rect 4728 4015 4762 4037
rect 4728 3969 4762 3977
rect 4728 3943 4762 3969
rect 4824 4887 4858 4913
rect 4824 4879 4858 4887
rect 4824 4819 4858 4841
rect 4824 4807 4858 4819
rect 4824 4751 4858 4769
rect 4824 4735 4858 4751
rect 4824 4683 4858 4697
rect 4824 4663 4858 4683
rect 4824 4615 4858 4625
rect 4824 4591 4858 4615
rect 4824 4547 4858 4553
rect 4824 4519 4858 4547
rect 4824 4479 4858 4481
rect 4824 4447 4858 4479
rect 4824 4377 4858 4409
rect 4824 4375 4858 4377
rect 4824 4309 4858 4337
rect 4824 4303 4858 4309
rect 4824 4241 4858 4265
rect 4824 4231 4858 4241
rect 4824 4173 4858 4193
rect 4824 4159 4858 4173
rect 4824 4105 4858 4121
rect 4824 4087 4858 4105
rect 4824 4037 4858 4049
rect 4824 4015 4858 4037
rect 4824 3969 4858 3977
rect 4824 3943 4858 3969
rect 7470 4887 7504 4913
rect 7470 4879 7504 4887
rect 7470 4819 7504 4841
rect 7470 4807 7504 4819
rect 7470 4751 7504 4769
rect 7470 4735 7504 4751
rect 7470 4683 7504 4697
rect 7470 4663 7504 4683
rect 7470 4615 7504 4625
rect 7470 4591 7504 4615
rect 7470 4547 7504 4553
rect 7470 4519 7504 4547
rect 7470 4479 7504 4481
rect 7470 4447 7504 4479
rect 7470 4377 7504 4409
rect 7470 4375 7504 4377
rect 7470 4309 7504 4337
rect 7470 4303 7504 4309
rect 7470 4241 7504 4265
rect 7470 4231 7504 4241
rect 7470 4173 7504 4193
rect 7470 4159 7504 4173
rect 7470 4105 7504 4121
rect 7470 4087 7504 4105
rect 7470 4037 7504 4049
rect 7470 4015 7504 4037
rect 7470 3969 7504 3977
rect 7470 3943 7504 3969
rect 7566 4887 7600 4913
rect 7566 4879 7600 4887
rect 7566 4819 7600 4841
rect 7566 4807 7600 4819
rect 7566 4751 7600 4769
rect 7566 4735 7600 4751
rect 7566 4683 7600 4697
rect 7566 4663 7600 4683
rect 7566 4615 7600 4625
rect 7566 4591 7600 4615
rect 7566 4547 7600 4553
rect 7566 4519 7600 4547
rect 7566 4479 7600 4481
rect 7566 4447 7600 4479
rect 7566 4377 7600 4409
rect 7566 4375 7600 4377
rect 7566 4309 7600 4337
rect 7566 4303 7600 4309
rect 7566 4241 7600 4265
rect 7566 4231 7600 4241
rect 7566 4173 7600 4193
rect 7566 4159 7600 4173
rect 7566 4105 7600 4121
rect 7566 4087 7600 4105
rect 7566 4037 7600 4049
rect 7566 4015 7600 4037
rect 7566 3969 7600 3977
rect 7566 3943 7600 3969
rect -4814 3841 -4780 3847
rect -4814 3779 -4780 3803
rect -4814 3769 -4780 3779
rect 1580 3743 1614 3777
rect 7662 4887 7696 4913
rect 7662 4879 7696 4887
rect 7662 4819 7696 4841
rect 7662 4807 7696 4819
rect 7662 4751 7696 4769
rect 7662 4735 7696 4751
rect 7662 4683 7696 4697
rect 7662 4663 7696 4683
rect 7662 4615 7696 4625
rect 7662 4591 7696 4615
rect 7662 4547 7696 4553
rect 7662 4519 7696 4547
rect 7662 4479 7696 4481
rect 7662 4447 7696 4479
rect 7662 4377 7696 4409
rect 7662 4375 7696 4377
rect 7662 4309 7696 4337
rect 7662 4303 7696 4309
rect 7662 4241 7696 4265
rect 7662 4231 7696 4241
rect 7662 4173 7696 4193
rect 7662 4159 7696 4173
rect 7662 4105 7696 4121
rect 7662 4087 7696 4105
rect 7662 4037 7696 4049
rect 7662 4015 7696 4037
rect 7662 3969 7696 3977
rect 7662 3943 7696 3969
rect 7758 4887 7792 4913
rect 7758 4879 7792 4887
rect 7758 4819 7792 4841
rect 7758 4807 7792 4819
rect 7758 4751 7792 4769
rect 7758 4735 7792 4751
rect 7758 4683 7792 4697
rect 7758 4663 7792 4683
rect 7758 4615 7792 4625
rect 7758 4591 7792 4615
rect 7758 4547 7792 4553
rect 7758 4519 7792 4547
rect 7758 4479 7792 4481
rect 7758 4447 7792 4479
rect 7758 4377 7792 4409
rect 7758 4375 7792 4377
rect 7758 4309 7792 4337
rect 7758 4303 7792 4309
rect 7758 4241 7792 4265
rect 7758 4231 7792 4241
rect 7758 4173 7792 4193
rect 7758 4159 7792 4173
rect 7758 4105 7792 4121
rect 7758 4087 7792 4105
rect 7758 4037 7792 4049
rect 7758 4015 7792 4037
rect 7758 3969 7792 3977
rect 7758 3943 7792 3969
rect 15518 5079 15552 5087
rect 15518 5053 15552 5079
rect 15518 5011 15552 5015
rect 7854 4887 7888 4913
rect 7854 4879 7888 4887
rect 7854 4819 7888 4841
rect 7854 4807 7888 4819
rect 7854 4751 7888 4769
rect 7854 4735 7888 4751
rect 7854 4683 7888 4697
rect 7854 4663 7888 4683
rect 7854 4615 7888 4625
rect 7854 4591 7888 4615
rect 7854 4547 7888 4553
rect 7854 4519 7888 4547
rect 7854 4479 7888 4481
rect 7854 4447 7888 4479
rect 7854 4377 7888 4409
rect 7854 4375 7888 4377
rect 7854 4309 7888 4337
rect 7854 4303 7888 4309
rect 7854 4241 7888 4265
rect 7854 4231 7888 4241
rect 7854 4173 7888 4193
rect 7854 4159 7888 4173
rect 7854 4105 7888 4121
rect 7854 4087 7888 4105
rect 7854 4037 7888 4049
rect 7854 4015 7888 4037
rect 7854 3969 7888 3977
rect 7854 3943 7888 3969
rect 10558 4885 10592 4911
rect 10558 4877 10592 4885
rect 10558 4817 10592 4839
rect 10558 4805 10592 4817
rect 10558 4749 10592 4767
rect 10558 4733 10592 4749
rect 10558 4681 10592 4695
rect 10558 4661 10592 4681
rect 10558 4613 10592 4623
rect 10558 4589 10592 4613
rect 10558 4545 10592 4551
rect 10558 4517 10592 4545
rect 10558 4477 10592 4479
rect 10558 4445 10592 4477
rect 10558 4375 10592 4407
rect 10558 4373 10592 4375
rect 10558 4307 10592 4335
rect 10558 4301 10592 4307
rect 10558 4239 10592 4263
rect 10558 4229 10592 4239
rect 10558 4171 10592 4191
rect 10558 4157 10592 4171
rect 10558 4103 10592 4119
rect 10558 4085 10592 4103
rect 10558 4035 10592 4047
rect 10558 4013 10592 4035
rect 10558 3967 10592 3975
rect 10558 3941 10592 3967
rect 10654 4885 10688 4911
rect 10654 4877 10688 4885
rect 10654 4817 10688 4839
rect 10654 4805 10688 4817
rect 10654 4749 10688 4767
rect 10654 4733 10688 4749
rect 10654 4681 10688 4695
rect 10654 4661 10688 4681
rect 10654 4613 10688 4623
rect 10654 4589 10688 4613
rect 10654 4545 10688 4551
rect 10654 4517 10688 4545
rect 10654 4477 10688 4479
rect 10654 4445 10688 4477
rect 10654 4375 10688 4407
rect 10654 4373 10688 4375
rect 10654 4307 10688 4335
rect 10654 4301 10688 4307
rect 10654 4239 10688 4263
rect 10654 4229 10688 4239
rect 10654 4171 10688 4191
rect 10654 4157 10688 4171
rect 10654 4103 10688 4119
rect 10654 4085 10688 4103
rect 10654 4035 10688 4047
rect 10654 4013 10688 4035
rect 10654 3967 10688 3975
rect 10654 3941 10688 3967
rect 10750 4885 10784 4911
rect 10750 4877 10784 4885
rect 10750 4817 10784 4839
rect 10750 4805 10784 4817
rect 10750 4749 10784 4767
rect 10750 4733 10784 4749
rect 10750 4681 10784 4695
rect 10750 4661 10784 4681
rect 10750 4613 10784 4623
rect 10750 4589 10784 4613
rect 10750 4545 10784 4551
rect 10750 4517 10784 4545
rect 10750 4477 10784 4479
rect 10750 4445 10784 4477
rect 10750 4375 10784 4407
rect 10750 4373 10784 4375
rect 10750 4307 10784 4335
rect 10750 4301 10784 4307
rect 10750 4239 10784 4263
rect 10750 4229 10784 4239
rect 10750 4171 10784 4191
rect 10750 4157 10784 4171
rect 10750 4103 10784 4119
rect 10750 4085 10784 4103
rect 10750 4035 10784 4047
rect 10750 4013 10784 4035
rect 10750 3967 10784 3975
rect 10750 3941 10784 3967
rect 10846 4885 10880 4911
rect 10846 4877 10880 4885
rect 10846 4817 10880 4839
rect 10846 4805 10880 4817
rect 10846 4749 10880 4767
rect 10846 4733 10880 4749
rect 10846 4681 10880 4695
rect 10846 4661 10880 4681
rect 10846 4613 10880 4623
rect 10846 4589 10880 4613
rect 10846 4545 10880 4551
rect 10846 4517 10880 4545
rect 10846 4477 10880 4479
rect 10846 4445 10880 4477
rect 10846 4375 10880 4407
rect 10846 4373 10880 4375
rect 10846 4307 10880 4335
rect 10846 4301 10880 4307
rect 10846 4239 10880 4263
rect 10846 4229 10880 4239
rect 10846 4171 10880 4191
rect 10846 4157 10880 4171
rect 10846 4103 10880 4119
rect 10846 4085 10880 4103
rect 10846 4035 10880 4047
rect 10846 4013 10880 4035
rect 10846 3967 10880 3975
rect 10846 3941 10880 3967
rect 15518 4981 15552 5011
rect 10942 4885 10976 4911
rect 10942 4877 10976 4885
rect 10942 4817 10976 4839
rect 10942 4805 10976 4817
rect 10942 4749 10976 4767
rect 10942 4733 10976 4749
rect 10942 4681 10976 4695
rect 10942 4661 10976 4681
rect 10942 4613 10976 4623
rect 10942 4589 10976 4613
rect 10942 4545 10976 4551
rect 10942 4517 10976 4545
rect 10942 4477 10976 4479
rect 10942 4445 10976 4477
rect 10942 4375 10976 4407
rect 10942 4373 10976 4375
rect 10942 4307 10976 4335
rect 10942 4301 10976 4307
rect 10942 4239 10976 4263
rect 10942 4229 10976 4239
rect 10942 4171 10976 4191
rect 10942 4157 10976 4171
rect 10942 4103 10976 4119
rect 10942 4085 10976 4103
rect 10942 4035 10976 4047
rect 10942 4013 10976 4035
rect 10942 3967 10976 3975
rect 10942 3941 10976 3967
rect 13714 4859 13748 4885
rect 13714 4851 13748 4859
rect 13714 4791 13748 4813
rect 13714 4779 13748 4791
rect 13714 4723 13748 4741
rect 13714 4707 13748 4723
rect 13714 4655 13748 4669
rect 13714 4635 13748 4655
rect 13714 4587 13748 4597
rect 13714 4563 13748 4587
rect 13714 4519 13748 4525
rect 13714 4491 13748 4519
rect 13714 4451 13748 4453
rect 13714 4419 13748 4451
rect 13714 4349 13748 4381
rect 13714 4347 13748 4349
rect 13714 4281 13748 4309
rect 13714 4275 13748 4281
rect 13714 4213 13748 4237
rect 13714 4203 13748 4213
rect 13714 4145 13748 4165
rect 13714 4131 13748 4145
rect 13714 4077 13748 4093
rect 13714 4059 13748 4077
rect 13714 4009 13748 4021
rect 13714 3987 13748 4009
rect 13714 3941 13748 3949
rect 13714 3915 13748 3941
rect 13810 4859 13844 4885
rect 13810 4851 13844 4859
rect 13810 4791 13844 4813
rect 13810 4779 13844 4791
rect 13810 4723 13844 4741
rect 13810 4707 13844 4723
rect 13810 4655 13844 4669
rect 13810 4635 13844 4655
rect 13810 4587 13844 4597
rect 13810 4563 13844 4587
rect 13810 4519 13844 4525
rect 13810 4491 13844 4519
rect 13810 4451 13844 4453
rect 13810 4419 13844 4451
rect 13810 4349 13844 4381
rect 13810 4347 13844 4349
rect 13810 4281 13844 4309
rect 13810 4275 13844 4281
rect 13810 4213 13844 4237
rect 13810 4203 13844 4213
rect 13810 4145 13844 4165
rect 13810 4131 13844 4145
rect 13810 4077 13844 4093
rect 13810 4059 13844 4077
rect 13810 4009 13844 4021
rect 13810 3987 13844 4009
rect 13810 3941 13844 3949
rect 13810 3915 13844 3941
rect -4814 3711 -4780 3731
rect 1676 3720 1710 3754
rect 1772 3743 1806 3777
rect 4536 3727 4570 3761
rect -4814 3697 -4780 3711
rect 4632 3704 4666 3738
rect 4728 3727 4762 3761
rect 7566 3727 7600 3761
rect 13906 4859 13940 4885
rect 13906 4851 13940 4859
rect 13906 4791 13940 4813
rect 13906 4779 13940 4791
rect 13906 4723 13940 4741
rect 13906 4707 13940 4723
rect 13906 4655 13940 4669
rect 13906 4635 13940 4655
rect 13906 4587 13940 4597
rect 13906 4563 13940 4587
rect 13906 4519 13940 4525
rect 13906 4491 13940 4519
rect 13906 4451 13940 4453
rect 13906 4419 13940 4451
rect 13906 4349 13940 4381
rect 13906 4347 13940 4349
rect 13906 4281 13940 4309
rect 13906 4275 13940 4281
rect 13906 4213 13940 4237
rect 13906 4203 13940 4213
rect 13906 4145 13940 4165
rect 13906 4131 13940 4145
rect 13906 4077 13940 4093
rect 13906 4059 13940 4077
rect 13906 4009 13940 4021
rect 13906 3987 13940 4009
rect 13906 3941 13940 3949
rect 13906 3915 13940 3941
rect 14002 4859 14036 4885
rect 14002 4851 14036 4859
rect 14002 4791 14036 4813
rect 14002 4779 14036 4791
rect 14002 4723 14036 4741
rect 14002 4707 14036 4723
rect 14002 4655 14036 4669
rect 14002 4635 14036 4655
rect 14002 4587 14036 4597
rect 14002 4563 14036 4587
rect 14002 4519 14036 4525
rect 14002 4491 14036 4519
rect 14002 4451 14036 4453
rect 14002 4419 14036 4451
rect 14002 4349 14036 4381
rect 14002 4347 14036 4349
rect 14002 4281 14036 4309
rect 14002 4275 14036 4281
rect 14002 4213 14036 4237
rect 14002 4203 14036 4213
rect 14002 4145 14036 4165
rect 14002 4131 14036 4145
rect 14002 4077 14036 4093
rect 14002 4059 14036 4077
rect 14002 4009 14036 4021
rect 14002 3987 14036 4009
rect 14002 3941 14036 3949
rect 14002 3915 14036 3941
rect 14098 4859 14132 4885
rect 14098 4851 14132 4859
rect 14098 4791 14132 4813
rect 14098 4779 14132 4791
rect 14098 4723 14132 4741
rect 14098 4707 14132 4723
rect 14098 4655 14132 4669
rect 14098 4635 14132 4655
rect 14098 4587 14132 4597
rect 14098 4563 14132 4587
rect 14098 4519 14132 4525
rect 14098 4491 14132 4519
rect 14098 4451 14132 4453
rect 14098 4419 14132 4451
rect 14098 4349 14132 4381
rect 14098 4347 14132 4349
rect 14098 4281 14132 4309
rect 14098 4275 14132 4281
rect 14098 4213 14132 4237
rect 14098 4203 14132 4213
rect 14098 4145 14132 4165
rect 14098 4131 14132 4145
rect 14098 4077 14132 4093
rect 14098 4059 14132 4077
rect 14098 4009 14132 4021
rect 14098 3987 14132 4009
rect 14098 3941 14132 3949
rect 14098 3915 14132 3941
rect 15518 4909 15552 4943
rect 15518 4841 15552 4871
rect 15518 4837 15552 4841
rect 15518 4773 15552 4799
rect 15518 4765 15552 4773
rect 15518 4705 15552 4727
rect 15518 4693 15552 4705
rect 15518 4637 15552 4655
rect 15518 4621 15552 4637
rect 15518 4569 15552 4583
rect 15518 4549 15552 4569
rect 15518 4501 15552 4511
rect 15518 4477 15552 4501
rect 15518 4433 15552 4439
rect 15518 4405 15552 4433
rect 15518 4365 15552 4367
rect 15518 4333 15552 4365
rect 15518 4263 15552 4295
rect 15518 4261 15552 4263
rect 15518 4195 15552 4223
rect 15518 4189 15552 4195
rect 15518 4127 15552 4151
rect 15518 4117 15552 4127
rect 15518 4059 15552 4079
rect 15518 4045 15552 4059
rect 15518 3991 15552 4007
rect 15518 3973 15552 3991
rect 15614 5861 15648 5879
rect 15614 5845 15648 5861
rect 15614 5793 15648 5807
rect 15614 5773 15648 5793
rect 15614 5725 15648 5735
rect 15614 5701 15648 5725
rect 15614 5657 15648 5663
rect 15614 5629 15648 5657
rect 15614 5589 15648 5591
rect 15614 5557 15648 5589
rect 15614 5487 15648 5519
rect 15614 5485 15648 5487
rect 15614 5419 15648 5447
rect 15614 5413 15648 5419
rect 15614 5351 15648 5375
rect 15614 5341 15648 5351
rect 15614 5283 15648 5303
rect 15614 5269 15648 5283
rect 15614 5215 15648 5231
rect 15614 5197 15648 5215
rect 15614 5147 15648 5159
rect 15614 5125 15648 5147
rect 15614 5079 15648 5087
rect 15614 5053 15648 5079
rect 15614 5011 15648 5015
rect 15614 4981 15648 5011
rect 15614 4909 15648 4943
rect 15614 4841 15648 4871
rect 15614 4837 15648 4841
rect 15614 4773 15648 4799
rect 15614 4765 15648 4773
rect 15614 4705 15648 4727
rect 15614 4693 15648 4705
rect 15614 4637 15648 4655
rect 15614 4621 15648 4637
rect 15614 4569 15648 4583
rect 15614 4549 15648 4569
rect 15614 4501 15648 4511
rect 15614 4477 15648 4501
rect 15614 4433 15648 4439
rect 15614 4405 15648 4433
rect 15614 4365 15648 4367
rect 15614 4333 15648 4365
rect 15614 4263 15648 4295
rect 15614 4261 15648 4263
rect 15614 4195 15648 4223
rect 15614 4189 15648 4195
rect 15614 4127 15648 4151
rect 15614 4117 15648 4127
rect 15614 4059 15648 4079
rect 15614 4045 15648 4059
rect 15614 3991 15648 4007
rect 15614 3973 15648 3991
rect 15710 5861 15744 5879
rect 15710 5845 15744 5861
rect 15710 5793 15744 5807
rect 15710 5773 15744 5793
rect 15710 5725 15744 5735
rect 15710 5701 15744 5725
rect 15710 5657 15744 5663
rect 15710 5629 15744 5657
rect 15710 5589 15744 5591
rect 15710 5557 15744 5589
rect 15710 5487 15744 5519
rect 15710 5485 15744 5487
rect 15710 5419 15744 5447
rect 15710 5413 15744 5419
rect 15710 5351 15744 5375
rect 15710 5341 15744 5351
rect 15710 5283 15744 5303
rect 17019 5344 17197 5450
rect 19014 5336 19192 5442
rect 21017 5338 21195 5444
rect 23566 5341 23744 5447
rect 25603 5340 25709 5446
rect 27563 5335 27741 5441
rect 15710 5269 15744 5283
rect 15710 5215 15744 5231
rect 15710 5197 15744 5215
rect 15710 5147 15744 5159
rect 15710 5125 15744 5147
rect 15710 5079 15744 5087
rect 15710 5053 15744 5079
rect 15710 5011 15744 5015
rect 15710 4981 15744 5011
rect 15710 4909 15744 4943
rect 15710 4841 15744 4871
rect 15710 4837 15744 4841
rect 15710 4773 15744 4799
rect 15710 4765 15744 4773
rect 15710 4705 15744 4727
rect 15710 4693 15744 4705
rect 15710 4637 15744 4655
rect 15710 4621 15744 4637
rect 15710 4569 15744 4583
rect 15710 4549 15744 4569
rect 15710 4501 15744 4511
rect 15710 4477 15744 4501
rect 15710 4433 15744 4439
rect 15710 4405 15744 4433
rect 15710 4365 15744 4367
rect 15710 4333 15744 4365
rect 15710 4263 15744 4295
rect 15710 4261 15744 4263
rect 15710 4195 15744 4223
rect 15710 4189 15744 4195
rect 15710 4127 15744 4151
rect 15710 4117 15744 4127
rect 16782 5089 16816 5115
rect 16782 5081 16816 5089
rect 16782 5021 16816 5043
rect 16782 5009 16816 5021
rect 16782 4953 16816 4971
rect 16782 4937 16816 4953
rect 16782 4885 16816 4899
rect 16782 4865 16816 4885
rect 16782 4817 16816 4827
rect 16782 4793 16816 4817
rect 16782 4749 16816 4755
rect 16782 4721 16816 4749
rect 16782 4681 16816 4683
rect 16782 4649 16816 4681
rect 16782 4579 16816 4611
rect 16782 4577 16816 4579
rect 16782 4511 16816 4539
rect 16782 4505 16816 4511
rect 16782 4443 16816 4467
rect 16782 4433 16816 4443
rect 16782 4375 16816 4395
rect 16782 4361 16816 4375
rect 16782 4307 16816 4323
rect 16782 4289 16816 4307
rect 16782 4239 16816 4251
rect 16782 4217 16816 4239
rect 16782 4171 16816 4179
rect 16782 4145 16816 4171
rect 16878 5089 16912 5115
rect 16878 5081 16912 5089
rect 16878 5021 16912 5043
rect 16878 5009 16912 5021
rect 16878 4953 16912 4971
rect 16878 4937 16912 4953
rect 16878 4885 16912 4899
rect 16878 4865 16912 4885
rect 16878 4817 16912 4827
rect 16878 4793 16912 4817
rect 16878 4749 16912 4755
rect 16878 4721 16912 4749
rect 16878 4681 16912 4683
rect 16878 4649 16912 4681
rect 16878 4579 16912 4611
rect 16878 4577 16912 4579
rect 16878 4511 16912 4539
rect 16878 4505 16912 4511
rect 16878 4443 16912 4467
rect 16878 4433 16912 4443
rect 16878 4375 16912 4395
rect 16878 4361 16912 4375
rect 16878 4307 16912 4323
rect 16878 4289 16912 4307
rect 16878 4239 16912 4251
rect 16878 4217 16912 4239
rect 16878 4171 16912 4179
rect 16878 4145 16912 4171
rect 15710 4059 15744 4079
rect 16974 5089 17008 5115
rect 16974 5081 17008 5089
rect 16974 5021 17008 5043
rect 16974 5009 17008 5021
rect 16974 4953 17008 4971
rect 16974 4937 17008 4953
rect 16974 4885 17008 4899
rect 16974 4865 17008 4885
rect 16974 4817 17008 4827
rect 16974 4793 17008 4817
rect 16974 4749 17008 4755
rect 16974 4721 17008 4749
rect 16974 4681 17008 4683
rect 16974 4649 17008 4681
rect 16974 4579 17008 4611
rect 16974 4577 17008 4579
rect 16974 4511 17008 4539
rect 16974 4505 17008 4511
rect 16974 4443 17008 4467
rect 16974 4433 17008 4443
rect 16974 4375 17008 4395
rect 16974 4361 17008 4375
rect 16974 4307 17008 4323
rect 16974 4289 17008 4307
rect 16974 4239 17008 4251
rect 16974 4217 17008 4239
rect 16974 4171 17008 4179
rect 16974 4145 17008 4171
rect 17070 5089 17104 5115
rect 17070 5081 17104 5089
rect 17070 5021 17104 5043
rect 17070 5009 17104 5021
rect 17070 4953 17104 4971
rect 17070 4937 17104 4953
rect 17070 4885 17104 4899
rect 17070 4865 17104 4885
rect 17070 4817 17104 4827
rect 17070 4793 17104 4817
rect 17070 4749 17104 4755
rect 17070 4721 17104 4749
rect 17070 4681 17104 4683
rect 17070 4649 17104 4681
rect 17070 4579 17104 4611
rect 17070 4577 17104 4579
rect 17070 4511 17104 4539
rect 17070 4505 17104 4511
rect 17070 4443 17104 4467
rect 17070 4433 17104 4443
rect 17070 4375 17104 4395
rect 17070 4361 17104 4375
rect 17070 4307 17104 4323
rect 17070 4289 17104 4307
rect 17070 4239 17104 4251
rect 17070 4217 17104 4239
rect 17070 4171 17104 4179
rect 17070 4145 17104 4171
rect 17166 5089 17200 5115
rect 17166 5081 17200 5089
rect 17166 5021 17200 5043
rect 17166 5009 17200 5021
rect 17166 4953 17200 4971
rect 17166 4937 17200 4953
rect 17166 4885 17200 4899
rect 17166 4865 17200 4885
rect 17166 4817 17200 4827
rect 17166 4793 17200 4817
rect 17166 4749 17200 4755
rect 17166 4721 17200 4749
rect 17166 4681 17200 4683
rect 17166 4649 17200 4681
rect 17166 4579 17200 4611
rect 17166 4577 17200 4579
rect 17166 4511 17200 4539
rect 17166 4505 17200 4511
rect 17166 4443 17200 4467
rect 17166 4433 17200 4443
rect 17166 4375 17200 4395
rect 17166 4361 17200 4375
rect 17166 4307 17200 4323
rect 17166 4289 17200 4307
rect 17166 4239 17200 4251
rect 17166 4217 17200 4239
rect 17166 4171 17200 4179
rect 17166 4145 17200 4171
rect 17262 5089 17296 5115
rect 17262 5081 17296 5089
rect 17262 5021 17296 5043
rect 17262 5009 17296 5021
rect 17262 4953 17296 4971
rect 17262 4937 17296 4953
rect 17262 4885 17296 4899
rect 17262 4865 17296 4885
rect 17262 4817 17296 4827
rect 17262 4793 17296 4817
rect 17262 4749 17296 4755
rect 17262 4721 17296 4749
rect 17262 4681 17296 4683
rect 17262 4649 17296 4681
rect 17262 4579 17296 4611
rect 17262 4577 17296 4579
rect 17262 4511 17296 4539
rect 17262 4505 17296 4511
rect 17262 4443 17296 4467
rect 17262 4433 17296 4443
rect 17262 4375 17296 4395
rect 17262 4361 17296 4375
rect 17262 4307 17296 4323
rect 17262 4289 17296 4307
rect 17262 4239 17296 4251
rect 17262 4217 17296 4239
rect 17262 4171 17296 4179
rect 17262 4145 17296 4171
rect 17470 5087 17504 5113
rect 17470 5079 17504 5087
rect 17470 5019 17504 5041
rect 17470 5007 17504 5019
rect 17470 4951 17504 4969
rect 17470 4935 17504 4951
rect 17470 4883 17504 4897
rect 17470 4863 17504 4883
rect 17470 4815 17504 4825
rect 17470 4791 17504 4815
rect 17470 4747 17504 4753
rect 17470 4719 17504 4747
rect 17470 4679 17504 4681
rect 17470 4647 17504 4679
rect 17470 4577 17504 4609
rect 17470 4575 17504 4577
rect 17470 4509 17504 4537
rect 17470 4503 17504 4509
rect 17470 4441 17504 4465
rect 17470 4431 17504 4441
rect 17470 4373 17504 4393
rect 17470 4359 17504 4373
rect 17470 4305 17504 4321
rect 17470 4287 17504 4305
rect 17470 4237 17504 4249
rect 17470 4215 17504 4237
rect 17470 4169 17504 4177
rect 17470 4143 17504 4169
rect 17566 5087 17600 5113
rect 17566 5079 17600 5087
rect 17566 5019 17600 5041
rect 17566 5007 17600 5019
rect 17566 4951 17600 4969
rect 17566 4935 17600 4951
rect 17566 4883 17600 4897
rect 17566 4863 17600 4883
rect 17566 4815 17600 4825
rect 17566 4791 17600 4815
rect 17566 4747 17600 4753
rect 17566 4719 17600 4747
rect 17566 4679 17600 4681
rect 17566 4647 17600 4679
rect 17566 4577 17600 4609
rect 17566 4575 17600 4577
rect 17566 4509 17600 4537
rect 17566 4503 17600 4509
rect 17566 4441 17600 4465
rect 17566 4431 17600 4441
rect 17566 4373 17600 4393
rect 17566 4359 17600 4373
rect 17566 4305 17600 4321
rect 17566 4287 17600 4305
rect 17566 4237 17600 4249
rect 17566 4215 17600 4237
rect 17566 4169 17600 4177
rect 17566 4143 17600 4169
rect 15710 4045 15744 4059
rect 17662 5087 17696 5113
rect 17662 5079 17696 5087
rect 17662 5019 17696 5041
rect 17662 5007 17696 5019
rect 17662 4951 17696 4969
rect 17662 4935 17696 4951
rect 17662 4883 17696 4897
rect 17662 4863 17696 4883
rect 17662 4815 17696 4825
rect 17662 4791 17696 4815
rect 17662 4747 17696 4753
rect 17662 4719 17696 4747
rect 17662 4679 17696 4681
rect 17662 4647 17696 4679
rect 17662 4577 17696 4609
rect 17662 4575 17696 4577
rect 17662 4509 17696 4537
rect 17662 4503 17696 4509
rect 17662 4441 17696 4465
rect 17662 4431 17696 4441
rect 17662 4373 17696 4393
rect 17662 4359 17696 4373
rect 17662 4305 17696 4321
rect 17662 4287 17696 4305
rect 17662 4237 17696 4249
rect 17662 4215 17696 4237
rect 17662 4169 17696 4177
rect 17662 4143 17696 4169
rect 17758 5087 17792 5113
rect 17758 5079 17792 5087
rect 17758 5019 17792 5041
rect 17758 5007 17792 5019
rect 17758 4951 17792 4969
rect 17758 4935 17792 4951
rect 17758 4883 17792 4897
rect 17758 4863 17792 4883
rect 17758 4815 17792 4825
rect 17758 4791 17792 4815
rect 17758 4747 17792 4753
rect 17758 4719 17792 4747
rect 17758 4679 17792 4681
rect 17758 4647 17792 4679
rect 17758 4577 17792 4609
rect 17758 4575 17792 4577
rect 17758 4509 17792 4537
rect 17758 4503 17792 4509
rect 17758 4441 17792 4465
rect 17758 4431 17792 4441
rect 17758 4373 17792 4393
rect 17758 4359 17792 4373
rect 17758 4305 17792 4321
rect 17758 4287 17792 4305
rect 17758 4237 17792 4249
rect 17758 4215 17792 4237
rect 17758 4169 17792 4177
rect 17758 4143 17792 4169
rect 17854 5087 17888 5113
rect 17854 5079 17888 5087
rect 17854 5019 17888 5041
rect 17854 5007 17888 5019
rect 17854 4951 17888 4969
rect 17854 4935 17888 4951
rect 17854 4883 17888 4897
rect 17854 4863 17888 4883
rect 17854 4815 17888 4825
rect 17854 4791 17888 4815
rect 17854 4747 17888 4753
rect 17854 4719 17888 4747
rect 17854 4679 17888 4681
rect 17854 4647 17888 4679
rect 17854 4577 17888 4609
rect 17854 4575 17888 4577
rect 17854 4509 17888 4537
rect 17854 4503 17888 4509
rect 17854 4441 17888 4465
rect 17854 4431 17888 4441
rect 17854 4373 17888 4393
rect 17854 4359 17888 4373
rect 17854 4305 17888 4321
rect 17854 4287 17888 4305
rect 17854 4237 17888 4249
rect 17854 4215 17888 4237
rect 17854 4169 17888 4177
rect 17854 4143 17888 4169
rect 17950 5087 17984 5113
rect 17950 5079 17984 5087
rect 17950 5019 17984 5041
rect 17950 5007 17984 5019
rect 17950 4951 17984 4969
rect 17950 4935 17984 4951
rect 17950 4883 17984 4897
rect 17950 4863 17984 4883
rect 17950 4815 17984 4825
rect 17950 4791 17984 4815
rect 17950 4747 17984 4753
rect 17950 4719 17984 4747
rect 17950 4679 17984 4681
rect 17950 4647 17984 4679
rect 17950 4577 17984 4609
rect 17950 4575 17984 4577
rect 17950 4509 17984 4537
rect 17950 4503 17984 4509
rect 17950 4441 17984 4465
rect 17950 4431 17984 4441
rect 17950 4373 17984 4393
rect 17950 4359 17984 4373
rect 17950 4305 17984 4321
rect 17950 4287 17984 4305
rect 17950 4237 17984 4249
rect 17950 4215 17984 4237
rect 17950 4169 17984 4177
rect 17950 4143 17984 4169
rect 18046 5087 18080 5113
rect 18046 5079 18080 5087
rect 18046 5019 18080 5041
rect 18046 5007 18080 5019
rect 18046 4951 18080 4969
rect 18046 4935 18080 4951
rect 18046 4883 18080 4897
rect 18046 4863 18080 4883
rect 18046 4815 18080 4825
rect 18046 4791 18080 4815
rect 18046 4747 18080 4753
rect 18046 4719 18080 4747
rect 18046 4679 18080 4681
rect 18046 4647 18080 4679
rect 18046 4577 18080 4609
rect 18046 4575 18080 4577
rect 18046 4509 18080 4537
rect 18046 4503 18080 4509
rect 18046 4441 18080 4465
rect 18046 4431 18080 4441
rect 18046 4373 18080 4393
rect 18046 4359 18080 4373
rect 18046 4305 18080 4321
rect 18046 4287 18080 4305
rect 18046 4237 18080 4249
rect 18046 4215 18080 4237
rect 18046 4169 18080 4177
rect 18046 4143 18080 4169
rect 18142 5087 18176 5113
rect 18142 5079 18176 5087
rect 18142 5019 18176 5041
rect 18142 5007 18176 5019
rect 18142 4951 18176 4969
rect 18142 4935 18176 4951
rect 18142 4883 18176 4897
rect 18142 4863 18176 4883
rect 18142 4815 18176 4825
rect 18142 4791 18176 4815
rect 18142 4747 18176 4753
rect 18142 4719 18176 4747
rect 18142 4679 18176 4681
rect 18142 4647 18176 4679
rect 18142 4577 18176 4609
rect 18142 4575 18176 4577
rect 18142 4509 18176 4537
rect 18142 4503 18176 4509
rect 18142 4441 18176 4465
rect 18142 4431 18176 4441
rect 18142 4373 18176 4393
rect 18142 4359 18176 4373
rect 18142 4305 18176 4321
rect 18142 4287 18176 4305
rect 18142 4237 18176 4249
rect 18142 4215 18176 4237
rect 18142 4169 18176 4177
rect 18142 4143 18176 4169
rect 18238 5087 18272 5113
rect 18238 5079 18272 5087
rect 18238 5019 18272 5041
rect 18238 5007 18272 5019
rect 18238 4951 18272 4969
rect 18238 4935 18272 4951
rect 18238 4883 18272 4897
rect 18238 4863 18272 4883
rect 18238 4815 18272 4825
rect 18238 4791 18272 4815
rect 18238 4747 18272 4753
rect 18238 4719 18272 4747
rect 18238 4679 18272 4681
rect 18238 4647 18272 4679
rect 18238 4577 18272 4609
rect 18238 4575 18272 4577
rect 18238 4509 18272 4537
rect 18238 4503 18272 4509
rect 18238 4441 18272 4465
rect 18238 4431 18272 4441
rect 18238 4373 18272 4393
rect 18238 4359 18272 4373
rect 18238 4305 18272 4321
rect 18238 4287 18272 4305
rect 18238 4237 18272 4249
rect 18238 4215 18272 4237
rect 18238 4169 18272 4177
rect 18238 4143 18272 4169
rect 18334 5087 18368 5113
rect 18334 5079 18368 5087
rect 18334 5019 18368 5041
rect 18334 5007 18368 5019
rect 18334 4951 18368 4969
rect 18334 4935 18368 4951
rect 18334 4883 18368 4897
rect 18334 4863 18368 4883
rect 18334 4815 18368 4825
rect 18334 4791 18368 4815
rect 18334 4747 18368 4753
rect 18334 4719 18368 4747
rect 18334 4679 18368 4681
rect 18334 4647 18368 4679
rect 18334 4577 18368 4609
rect 18334 4575 18368 4577
rect 18334 4509 18368 4537
rect 18334 4503 18368 4509
rect 18334 4441 18368 4465
rect 18334 4431 18368 4441
rect 18334 4373 18368 4393
rect 18334 4359 18368 4373
rect 18334 4305 18368 4321
rect 18334 4287 18368 4305
rect 18334 4237 18368 4249
rect 18334 4215 18368 4237
rect 18334 4169 18368 4177
rect 18334 4143 18368 4169
rect 18430 5087 18464 5113
rect 18430 5079 18464 5087
rect 18430 5019 18464 5041
rect 18430 5007 18464 5019
rect 18430 4951 18464 4969
rect 18430 4935 18464 4951
rect 18430 4883 18464 4897
rect 18430 4863 18464 4883
rect 18430 4815 18464 4825
rect 18430 4791 18464 4815
rect 18430 4747 18464 4753
rect 18430 4719 18464 4747
rect 18430 4679 18464 4681
rect 18430 4647 18464 4679
rect 18430 4577 18464 4609
rect 18430 4575 18464 4577
rect 18430 4509 18464 4537
rect 18430 4503 18464 4509
rect 18430 4441 18464 4465
rect 18430 4431 18464 4441
rect 18430 4373 18464 4393
rect 18430 4359 18464 4373
rect 18430 4305 18464 4321
rect 18430 4287 18464 4305
rect 18430 4237 18464 4249
rect 18430 4215 18464 4237
rect 18430 4169 18464 4177
rect 18430 4143 18464 4169
rect 18674 5081 18708 5107
rect 18674 5073 18708 5081
rect 18674 5013 18708 5035
rect 18674 5001 18708 5013
rect 18674 4945 18708 4963
rect 18674 4929 18708 4945
rect 18674 4877 18708 4891
rect 18674 4857 18708 4877
rect 18674 4809 18708 4819
rect 18674 4785 18708 4809
rect 18674 4741 18708 4747
rect 18674 4713 18708 4741
rect 18674 4673 18708 4675
rect 18674 4641 18708 4673
rect 18674 4571 18708 4603
rect 18674 4569 18708 4571
rect 18674 4503 18708 4531
rect 18674 4497 18708 4503
rect 18674 4435 18708 4459
rect 18674 4425 18708 4435
rect 18674 4367 18708 4387
rect 18674 4353 18708 4367
rect 18674 4299 18708 4315
rect 18674 4281 18708 4299
rect 18674 4231 18708 4243
rect 18674 4209 18708 4231
rect 18674 4163 18708 4171
rect 18674 4137 18708 4163
rect 18770 5081 18804 5107
rect 18770 5073 18804 5081
rect 18770 5013 18804 5035
rect 18770 5001 18804 5013
rect 18770 4945 18804 4963
rect 18770 4929 18804 4945
rect 18770 4877 18804 4891
rect 18770 4857 18804 4877
rect 18770 4809 18804 4819
rect 18770 4785 18804 4809
rect 18770 4741 18804 4747
rect 18770 4713 18804 4741
rect 18770 4673 18804 4675
rect 18770 4641 18804 4673
rect 18770 4571 18804 4603
rect 18770 4569 18804 4571
rect 18770 4503 18804 4531
rect 18770 4497 18804 4503
rect 18770 4435 18804 4459
rect 18770 4425 18804 4435
rect 18770 4367 18804 4387
rect 18770 4353 18804 4367
rect 18770 4299 18804 4315
rect 18770 4281 18804 4299
rect 18770 4231 18804 4243
rect 18770 4209 18804 4231
rect 18770 4163 18804 4171
rect 18770 4137 18804 4163
rect 15710 3991 15744 4007
rect 15710 3973 15744 3991
rect 16830 3909 16864 3943
rect 7662 3704 7696 3738
rect 7758 3727 7792 3761
rect 10654 3725 10688 3759
rect 10750 3702 10784 3736
rect 10846 3725 10880 3759
rect 13810 3699 13844 3733
rect 15566 3745 15600 3779
rect 13906 3676 13940 3710
rect 14002 3699 14036 3733
rect 15710 3726 15744 3760
rect 18866 5081 18900 5107
rect 18866 5073 18900 5081
rect 18866 5013 18900 5035
rect 18866 5001 18900 5013
rect 18866 4945 18900 4963
rect 18866 4929 18900 4945
rect 18866 4877 18900 4891
rect 18866 4857 18900 4877
rect 18866 4809 18900 4819
rect 18866 4785 18900 4809
rect 18866 4741 18900 4747
rect 18866 4713 18900 4741
rect 18866 4673 18900 4675
rect 18866 4641 18900 4673
rect 18866 4571 18900 4603
rect 18866 4569 18900 4571
rect 18866 4503 18900 4531
rect 18866 4497 18900 4503
rect 18866 4435 18900 4459
rect 18866 4425 18900 4435
rect 18866 4367 18900 4387
rect 18866 4353 18900 4367
rect 18866 4299 18900 4315
rect 18866 4281 18900 4299
rect 18866 4231 18900 4243
rect 18866 4209 18900 4231
rect 18866 4163 18900 4171
rect 18866 4137 18900 4163
rect 18962 5081 18996 5107
rect 18962 5073 18996 5081
rect 18962 5013 18996 5035
rect 18962 5001 18996 5013
rect 18962 4945 18996 4963
rect 18962 4929 18996 4945
rect 18962 4877 18996 4891
rect 18962 4857 18996 4877
rect 18962 4809 18996 4819
rect 18962 4785 18996 4809
rect 18962 4741 18996 4747
rect 18962 4713 18996 4741
rect 18962 4673 18996 4675
rect 18962 4641 18996 4673
rect 18962 4571 18996 4603
rect 18962 4569 18996 4571
rect 18962 4503 18996 4531
rect 18962 4497 18996 4503
rect 18962 4435 18996 4459
rect 18962 4425 18996 4435
rect 18962 4367 18996 4387
rect 18962 4353 18996 4367
rect 18962 4299 18996 4315
rect 18962 4281 18996 4299
rect 18962 4231 18996 4243
rect 18962 4209 18996 4231
rect 18962 4163 18996 4171
rect 18962 4137 18996 4163
rect 19058 5081 19092 5107
rect 19058 5073 19092 5081
rect 19058 5013 19092 5035
rect 19058 5001 19092 5013
rect 19058 4945 19092 4963
rect 19058 4929 19092 4945
rect 19058 4877 19092 4891
rect 19058 4857 19092 4877
rect 19058 4809 19092 4819
rect 19058 4785 19092 4809
rect 19058 4741 19092 4747
rect 19058 4713 19092 4741
rect 19058 4673 19092 4675
rect 19058 4641 19092 4673
rect 19058 4571 19092 4603
rect 19058 4569 19092 4571
rect 19058 4503 19092 4531
rect 19058 4497 19092 4503
rect 19058 4435 19092 4459
rect 19058 4425 19092 4435
rect 19058 4367 19092 4387
rect 19058 4353 19092 4367
rect 19058 4299 19092 4315
rect 19058 4281 19092 4299
rect 19058 4231 19092 4243
rect 19058 4209 19092 4231
rect 19058 4163 19092 4171
rect 19058 4137 19092 4163
rect 19154 5081 19188 5107
rect 19154 5073 19188 5081
rect 19154 5013 19188 5035
rect 19154 5001 19188 5013
rect 19154 4945 19188 4963
rect 19154 4929 19188 4945
rect 19154 4877 19188 4891
rect 19154 4857 19188 4877
rect 19154 4809 19188 4819
rect 19154 4785 19188 4809
rect 19154 4741 19188 4747
rect 19154 4713 19188 4741
rect 19154 4673 19188 4675
rect 19154 4641 19188 4673
rect 19154 4571 19188 4603
rect 19154 4569 19188 4571
rect 19154 4503 19188 4531
rect 19154 4497 19188 4503
rect 19154 4435 19188 4459
rect 19154 4425 19188 4435
rect 19154 4367 19188 4387
rect 19154 4353 19188 4367
rect 19154 4299 19188 4315
rect 19154 4281 19188 4299
rect 19154 4231 19188 4243
rect 19154 4209 19188 4231
rect 19154 4163 19188 4171
rect 19154 4137 19188 4163
rect 19250 5081 19284 5107
rect 19250 5073 19284 5081
rect 19250 5013 19284 5035
rect 19250 5001 19284 5013
rect 19250 4945 19284 4963
rect 19250 4929 19284 4945
rect 19250 4877 19284 4891
rect 19250 4857 19284 4877
rect 19250 4809 19284 4819
rect 19250 4785 19284 4809
rect 19250 4741 19284 4747
rect 19250 4713 19284 4741
rect 19250 4673 19284 4675
rect 19250 4641 19284 4673
rect 19250 4571 19284 4603
rect 19250 4569 19284 4571
rect 19250 4503 19284 4531
rect 19250 4497 19284 4503
rect 19250 4435 19284 4459
rect 19250 4425 19284 4435
rect 19250 4367 19284 4387
rect 19250 4353 19284 4367
rect 19250 4299 19284 4315
rect 19250 4281 19284 4299
rect 19250 4231 19284 4243
rect 19250 4209 19284 4231
rect 19250 4163 19284 4171
rect 19250 4137 19284 4163
rect 19346 5081 19380 5107
rect 19346 5073 19380 5081
rect 19346 5013 19380 5035
rect 19346 5001 19380 5013
rect 19346 4945 19380 4963
rect 19346 4929 19380 4945
rect 19346 4877 19380 4891
rect 19346 4857 19380 4877
rect 19346 4809 19380 4819
rect 19346 4785 19380 4809
rect 19346 4741 19380 4747
rect 19346 4713 19380 4741
rect 19346 4673 19380 4675
rect 19346 4641 19380 4673
rect 19346 4571 19380 4603
rect 19346 4569 19380 4571
rect 19346 4503 19380 4531
rect 19346 4497 19380 4503
rect 19346 4435 19380 4459
rect 19346 4425 19380 4435
rect 19346 4367 19380 4387
rect 19346 4353 19380 4367
rect 19346 4299 19380 4315
rect 19346 4281 19380 4299
rect 19346 4231 19380 4243
rect 19346 4209 19380 4231
rect 19346 4163 19380 4171
rect 19346 4137 19380 4163
rect 19442 5081 19476 5107
rect 19442 5073 19476 5081
rect 19442 5013 19476 5035
rect 19442 5001 19476 5013
rect 19442 4945 19476 4963
rect 19442 4929 19476 4945
rect 19442 4877 19476 4891
rect 19442 4857 19476 4877
rect 19442 4809 19476 4819
rect 19442 4785 19476 4809
rect 19442 4741 19476 4747
rect 19442 4713 19476 4741
rect 19442 4673 19476 4675
rect 19442 4641 19476 4673
rect 19442 4571 19476 4603
rect 19442 4569 19476 4571
rect 19442 4503 19476 4531
rect 19442 4497 19476 4503
rect 19442 4435 19476 4459
rect 19442 4425 19476 4435
rect 19442 4367 19476 4387
rect 19442 4353 19476 4367
rect 19442 4299 19476 4315
rect 19442 4281 19476 4299
rect 19442 4231 19476 4243
rect 19442 4209 19476 4231
rect 19442 4163 19476 4171
rect 19442 4137 19476 4163
rect 19538 5081 19572 5107
rect 19538 5073 19572 5081
rect 19538 5013 19572 5035
rect 19538 5001 19572 5013
rect 19538 4945 19572 4963
rect 19538 4929 19572 4945
rect 19538 4877 19572 4891
rect 19538 4857 19572 4877
rect 19538 4809 19572 4819
rect 19538 4785 19572 4809
rect 19538 4741 19572 4747
rect 19538 4713 19572 4741
rect 19538 4673 19572 4675
rect 19538 4641 19572 4673
rect 19538 4571 19572 4603
rect 19538 4569 19572 4571
rect 19538 4503 19572 4531
rect 19538 4497 19572 4503
rect 19538 4435 19572 4459
rect 19538 4425 19572 4435
rect 19538 4367 19572 4387
rect 19538 4353 19572 4367
rect 19538 4299 19572 4315
rect 19538 4281 19572 4299
rect 19538 4231 19572 4243
rect 19538 4209 19572 4231
rect 19538 4163 19572 4171
rect 19538 4137 19572 4163
rect 19634 5081 19668 5107
rect 19634 5073 19668 5081
rect 19634 5013 19668 5035
rect 19634 5001 19668 5013
rect 19634 4945 19668 4963
rect 19634 4929 19668 4945
rect 19634 4877 19668 4891
rect 19634 4857 19668 4877
rect 19634 4809 19668 4819
rect 19634 4785 19668 4809
rect 19634 4741 19668 4747
rect 19634 4713 19668 4741
rect 19634 4673 19668 4675
rect 19634 4641 19668 4673
rect 19634 4571 19668 4603
rect 19634 4569 19668 4571
rect 19634 4503 19668 4531
rect 19634 4497 19668 4503
rect 19634 4435 19668 4459
rect 19634 4425 19668 4435
rect 19634 4367 19668 4387
rect 19634 4353 19668 4367
rect 19634 4299 19668 4315
rect 19634 4281 19668 4299
rect 19634 4231 19668 4243
rect 19634 4209 19668 4231
rect 19634 4163 19668 4171
rect 19634 4137 19668 4163
rect 19730 5081 19764 5107
rect 19730 5073 19764 5081
rect 19730 5013 19764 5035
rect 19730 5001 19764 5013
rect 19730 4945 19764 4963
rect 19730 4929 19764 4945
rect 19730 4877 19764 4891
rect 19730 4857 19764 4877
rect 19730 4809 19764 4819
rect 19730 4785 19764 4809
rect 19730 4741 19764 4747
rect 19730 4713 19764 4741
rect 19730 4673 19764 4675
rect 19730 4641 19764 4673
rect 19730 4571 19764 4603
rect 19730 4569 19764 4571
rect 19730 4503 19764 4531
rect 19730 4497 19764 4503
rect 19730 4435 19764 4459
rect 19730 4425 19764 4435
rect 19730 4367 19764 4387
rect 19730 4353 19764 4367
rect 19730 4299 19764 4315
rect 19730 4281 19764 4299
rect 19730 4231 19764 4243
rect 19730 4209 19764 4231
rect 19730 4163 19764 4171
rect 19730 4137 19764 4163
rect 19826 5081 19860 5107
rect 19826 5073 19860 5081
rect 19826 5013 19860 5035
rect 19826 5001 19860 5013
rect 19826 4945 19860 4963
rect 19826 4929 19860 4945
rect 19826 4877 19860 4891
rect 19826 4857 19860 4877
rect 19826 4809 19860 4819
rect 19826 4785 19860 4809
rect 19826 4741 19860 4747
rect 19826 4713 19860 4741
rect 19826 4673 19860 4675
rect 19826 4641 19860 4673
rect 19826 4571 19860 4603
rect 19826 4569 19860 4571
rect 19826 4503 19860 4531
rect 19826 4497 19860 4503
rect 19826 4435 19860 4459
rect 19826 4425 19860 4435
rect 19826 4367 19860 4387
rect 19826 4353 19860 4367
rect 19826 4299 19860 4315
rect 19826 4281 19860 4299
rect 19826 4231 19860 4243
rect 19826 4209 19860 4231
rect 19826 4163 19860 4171
rect 19826 4137 19860 4163
rect 19922 5081 19956 5107
rect 19922 5073 19956 5081
rect 19922 5013 19956 5035
rect 19922 5001 19956 5013
rect 19922 4945 19956 4963
rect 19922 4929 19956 4945
rect 19922 4877 19956 4891
rect 19922 4857 19956 4877
rect 19922 4809 19956 4819
rect 19922 4785 19956 4809
rect 19922 4741 19956 4747
rect 19922 4713 19956 4741
rect 19922 4673 19956 4675
rect 19922 4641 19956 4673
rect 19922 4571 19956 4603
rect 19922 4569 19956 4571
rect 19922 4503 19956 4531
rect 19922 4497 19956 4503
rect 19922 4435 19956 4459
rect 19922 4425 19956 4435
rect 19922 4367 19956 4387
rect 19922 4353 19956 4367
rect 19922 4299 19956 4315
rect 19922 4281 19956 4299
rect 19922 4231 19956 4243
rect 19922 4209 19956 4231
rect 19922 4163 19956 4171
rect 19922 4137 19956 4163
rect 20018 5081 20052 5107
rect 20018 5073 20052 5081
rect 20018 5013 20052 5035
rect 20018 5001 20052 5013
rect 20018 4945 20052 4963
rect 20018 4929 20052 4945
rect 20018 4877 20052 4891
rect 20018 4857 20052 4877
rect 20018 4809 20052 4819
rect 20018 4785 20052 4809
rect 20018 4741 20052 4747
rect 20018 4713 20052 4741
rect 20018 4673 20052 4675
rect 20018 4641 20052 4673
rect 20018 4571 20052 4603
rect 20018 4569 20052 4571
rect 20018 4503 20052 4531
rect 20018 4497 20052 4503
rect 20018 4435 20052 4459
rect 20018 4425 20052 4435
rect 20018 4367 20052 4387
rect 20018 4353 20052 4367
rect 20018 4299 20052 4315
rect 20018 4281 20052 4299
rect 20018 4231 20052 4243
rect 20018 4209 20052 4231
rect 20018 4163 20052 4171
rect 20018 4137 20052 4163
rect 20114 5081 20148 5107
rect 20114 5073 20148 5081
rect 20114 5013 20148 5035
rect 20114 5001 20148 5013
rect 20114 4945 20148 4963
rect 20114 4929 20148 4945
rect 20114 4877 20148 4891
rect 20114 4857 20148 4877
rect 20114 4809 20148 4819
rect 20114 4785 20148 4809
rect 20114 4741 20148 4747
rect 20114 4713 20148 4741
rect 20114 4673 20148 4675
rect 20114 4641 20148 4673
rect 20114 4571 20148 4603
rect 20114 4569 20148 4571
rect 20114 4503 20148 4531
rect 20114 4497 20148 4503
rect 20114 4435 20148 4459
rect 20114 4425 20148 4435
rect 20114 4367 20148 4387
rect 20114 4353 20148 4367
rect 20114 4299 20148 4315
rect 20114 4281 20148 4299
rect 20114 4231 20148 4243
rect 20114 4209 20148 4231
rect 20114 4163 20148 4171
rect 20114 4137 20148 4163
rect 20338 5075 20372 5101
rect 20338 5067 20372 5075
rect 20338 5007 20372 5029
rect 20338 4995 20372 5007
rect 20338 4939 20372 4957
rect 20338 4923 20372 4939
rect 20338 4871 20372 4885
rect 20338 4851 20372 4871
rect 20338 4803 20372 4813
rect 20338 4779 20372 4803
rect 20338 4735 20372 4741
rect 20338 4707 20372 4735
rect 20338 4667 20372 4669
rect 20338 4635 20372 4667
rect 20338 4565 20372 4597
rect 20338 4563 20372 4565
rect 20338 4497 20372 4525
rect 20338 4491 20372 4497
rect 20338 4429 20372 4453
rect 20338 4419 20372 4429
rect 20338 4361 20372 4381
rect 20338 4347 20372 4361
rect 20338 4293 20372 4309
rect 20338 4275 20372 4293
rect 20338 4225 20372 4237
rect 20338 4203 20372 4225
rect 20338 4157 20372 4165
rect 20338 4131 20372 4157
rect 20434 5075 20468 5101
rect 20434 5067 20468 5075
rect 20434 5007 20468 5029
rect 20434 4995 20468 5007
rect 20434 4939 20468 4957
rect 20434 4923 20468 4939
rect 20434 4871 20468 4885
rect 20434 4851 20468 4871
rect 20434 4803 20468 4813
rect 20434 4779 20468 4803
rect 20434 4735 20468 4741
rect 20434 4707 20468 4735
rect 20434 4667 20468 4669
rect 20434 4635 20468 4667
rect 20434 4565 20468 4597
rect 20434 4563 20468 4565
rect 20434 4497 20468 4525
rect 20434 4491 20468 4497
rect 20434 4429 20468 4453
rect 20434 4419 20468 4429
rect 20434 4361 20468 4381
rect 20434 4347 20468 4361
rect 20434 4293 20468 4309
rect 20434 4275 20468 4293
rect 20434 4225 20468 4237
rect 20434 4203 20468 4225
rect 20434 4157 20468 4165
rect 20434 4131 20468 4157
rect 17518 3927 17552 3961
rect 16974 3787 17008 3821
rect 16830 3672 16864 3706
rect -4814 3643 -4780 3659
rect -4814 3625 -4780 3643
rect 20530 5075 20564 5101
rect 20530 5067 20564 5075
rect 20530 5007 20564 5029
rect 20530 4995 20564 5007
rect 20530 4939 20564 4957
rect 20530 4923 20564 4939
rect 20530 4871 20564 4885
rect 20530 4851 20564 4871
rect 20530 4803 20564 4813
rect 20530 4779 20564 4803
rect 20530 4735 20564 4741
rect 20530 4707 20564 4735
rect 20530 4667 20564 4669
rect 20530 4635 20564 4667
rect 20530 4565 20564 4597
rect 20530 4563 20564 4565
rect 20530 4497 20564 4525
rect 20530 4491 20564 4497
rect 20530 4429 20564 4453
rect 20530 4419 20564 4429
rect 20530 4361 20564 4381
rect 20530 4347 20564 4361
rect 20530 4293 20564 4309
rect 20530 4275 20564 4293
rect 20530 4225 20564 4237
rect 20530 4203 20564 4225
rect 20530 4157 20564 4165
rect 20530 4131 20564 4157
rect 20626 5075 20660 5101
rect 20626 5067 20660 5075
rect 20626 5007 20660 5029
rect 20626 4995 20660 5007
rect 20626 4939 20660 4957
rect 20626 4923 20660 4939
rect 20626 4871 20660 4885
rect 20626 4851 20660 4871
rect 20626 4803 20660 4813
rect 20626 4779 20660 4803
rect 20626 4735 20660 4741
rect 20626 4707 20660 4735
rect 20626 4667 20660 4669
rect 20626 4635 20660 4667
rect 20626 4565 20660 4597
rect 20626 4563 20660 4565
rect 20626 4497 20660 4525
rect 20626 4491 20660 4497
rect 20626 4429 20660 4453
rect 20626 4419 20660 4429
rect 20626 4361 20660 4381
rect 20626 4347 20660 4361
rect 20626 4293 20660 4309
rect 20626 4275 20660 4293
rect 20626 4225 20660 4237
rect 20626 4203 20660 4225
rect 20626 4157 20660 4165
rect 20626 4131 20660 4157
rect 20722 5075 20756 5101
rect 20722 5067 20756 5075
rect 20722 5007 20756 5029
rect 20722 4995 20756 5007
rect 20722 4939 20756 4957
rect 20722 4923 20756 4939
rect 20722 4871 20756 4885
rect 20722 4851 20756 4871
rect 20722 4803 20756 4813
rect 20722 4779 20756 4803
rect 20722 4735 20756 4741
rect 20722 4707 20756 4735
rect 20722 4667 20756 4669
rect 20722 4635 20756 4667
rect 20722 4565 20756 4597
rect 20722 4563 20756 4565
rect 20722 4497 20756 4525
rect 20722 4491 20756 4497
rect 20722 4429 20756 4453
rect 20722 4419 20756 4429
rect 20722 4361 20756 4381
rect 20722 4347 20756 4361
rect 20722 4293 20756 4309
rect 20722 4275 20756 4293
rect 20722 4225 20756 4237
rect 20722 4203 20756 4225
rect 20722 4157 20756 4165
rect 20722 4131 20756 4157
rect 20818 5075 20852 5101
rect 20818 5067 20852 5075
rect 20818 5007 20852 5029
rect 20818 4995 20852 5007
rect 20818 4939 20852 4957
rect 20818 4923 20852 4939
rect 20818 4871 20852 4885
rect 20818 4851 20852 4871
rect 20818 4803 20852 4813
rect 20818 4779 20852 4803
rect 20818 4735 20852 4741
rect 20818 4707 20852 4735
rect 20818 4667 20852 4669
rect 20818 4635 20852 4667
rect 20818 4565 20852 4597
rect 20818 4563 20852 4565
rect 20818 4497 20852 4525
rect 20818 4491 20852 4497
rect 20818 4429 20852 4453
rect 20818 4419 20852 4429
rect 20818 4361 20852 4381
rect 20818 4347 20852 4361
rect 20818 4293 20852 4309
rect 20818 4275 20852 4293
rect 20818 4225 20852 4237
rect 20818 4203 20852 4225
rect 20818 4157 20852 4165
rect 20818 4131 20852 4157
rect 20914 5075 20948 5101
rect 20914 5067 20948 5075
rect 20914 5007 20948 5029
rect 20914 4995 20948 5007
rect 20914 4939 20948 4957
rect 20914 4923 20948 4939
rect 20914 4871 20948 4885
rect 20914 4851 20948 4871
rect 20914 4803 20948 4813
rect 20914 4779 20948 4803
rect 20914 4735 20948 4741
rect 20914 4707 20948 4735
rect 20914 4667 20948 4669
rect 20914 4635 20948 4667
rect 20914 4565 20948 4597
rect 20914 4563 20948 4565
rect 20914 4497 20948 4525
rect 20914 4491 20948 4497
rect 20914 4429 20948 4453
rect 20914 4419 20948 4429
rect 20914 4361 20948 4381
rect 20914 4347 20948 4361
rect 20914 4293 20948 4309
rect 20914 4275 20948 4293
rect 20914 4225 20948 4237
rect 20914 4203 20948 4225
rect 20914 4157 20948 4165
rect 20914 4131 20948 4157
rect 21010 5075 21044 5101
rect 21010 5067 21044 5075
rect 21010 5007 21044 5029
rect 21010 4995 21044 5007
rect 21010 4939 21044 4957
rect 21010 4923 21044 4939
rect 21010 4871 21044 4885
rect 21010 4851 21044 4871
rect 21010 4803 21044 4813
rect 21010 4779 21044 4803
rect 21010 4735 21044 4741
rect 21010 4707 21044 4735
rect 21010 4667 21044 4669
rect 21010 4635 21044 4667
rect 21010 4565 21044 4597
rect 21010 4563 21044 4565
rect 21010 4497 21044 4525
rect 21010 4491 21044 4497
rect 21010 4429 21044 4453
rect 21010 4419 21044 4429
rect 21010 4361 21044 4381
rect 21010 4347 21044 4361
rect 21010 4293 21044 4309
rect 21010 4275 21044 4293
rect 21010 4225 21044 4237
rect 21010 4203 21044 4225
rect 21010 4157 21044 4165
rect 21010 4131 21044 4157
rect 21106 5075 21140 5101
rect 21106 5067 21140 5075
rect 21106 5007 21140 5029
rect 21106 4995 21140 5007
rect 21106 4939 21140 4957
rect 21106 4923 21140 4939
rect 21106 4871 21140 4885
rect 21106 4851 21140 4871
rect 21106 4803 21140 4813
rect 21106 4779 21140 4803
rect 21106 4735 21140 4741
rect 21106 4707 21140 4735
rect 21106 4667 21140 4669
rect 21106 4635 21140 4667
rect 21106 4565 21140 4597
rect 21106 4563 21140 4565
rect 21106 4497 21140 4525
rect 21106 4491 21140 4497
rect 21106 4429 21140 4453
rect 21106 4419 21140 4429
rect 21106 4361 21140 4381
rect 21106 4347 21140 4361
rect 21106 4293 21140 4309
rect 21106 4275 21140 4293
rect 21106 4225 21140 4237
rect 21106 4203 21140 4225
rect 21106 4157 21140 4165
rect 21106 4131 21140 4157
rect 21202 5075 21236 5101
rect 21202 5067 21236 5075
rect 21202 5007 21236 5029
rect 21202 4995 21236 5007
rect 21202 4939 21236 4957
rect 21202 4923 21236 4939
rect 21202 4871 21236 4885
rect 21202 4851 21236 4871
rect 21202 4803 21236 4813
rect 21202 4779 21236 4803
rect 21202 4735 21236 4741
rect 21202 4707 21236 4735
rect 21202 4667 21236 4669
rect 21202 4635 21236 4667
rect 21202 4565 21236 4597
rect 21202 4563 21236 4565
rect 21202 4497 21236 4525
rect 21202 4491 21236 4497
rect 21202 4429 21236 4453
rect 21202 4419 21236 4429
rect 21202 4361 21236 4381
rect 21202 4347 21236 4361
rect 21202 4293 21236 4309
rect 21202 4275 21236 4293
rect 21202 4225 21236 4237
rect 21202 4203 21236 4225
rect 21202 4157 21236 4165
rect 21202 4131 21236 4157
rect 21298 5075 21332 5101
rect 21298 5067 21332 5075
rect 21298 5007 21332 5029
rect 21298 4995 21332 5007
rect 21298 4939 21332 4957
rect 21298 4923 21332 4939
rect 21298 4871 21332 4885
rect 21298 4851 21332 4871
rect 21298 4803 21332 4813
rect 21298 4779 21332 4803
rect 21298 4735 21332 4741
rect 21298 4707 21332 4735
rect 21298 4667 21332 4669
rect 21298 4635 21332 4667
rect 21298 4565 21332 4597
rect 21298 4563 21332 4565
rect 21298 4497 21332 4525
rect 21298 4491 21332 4497
rect 21298 4429 21332 4453
rect 21298 4419 21332 4429
rect 21298 4361 21332 4381
rect 21298 4347 21332 4361
rect 21298 4293 21332 4309
rect 21298 4275 21332 4293
rect 21298 4225 21332 4237
rect 21298 4203 21332 4225
rect 21298 4157 21332 4165
rect 21298 4131 21332 4157
rect 21394 5075 21428 5101
rect 21394 5067 21428 5075
rect 21394 5007 21428 5029
rect 21394 4995 21428 5007
rect 21394 4939 21428 4957
rect 21394 4923 21428 4939
rect 21394 4871 21428 4885
rect 21394 4851 21428 4871
rect 21394 4803 21428 4813
rect 21394 4779 21428 4803
rect 21394 4735 21428 4741
rect 21394 4707 21428 4735
rect 21394 4667 21428 4669
rect 21394 4635 21428 4667
rect 21394 4565 21428 4597
rect 21394 4563 21428 4565
rect 21394 4497 21428 4525
rect 21394 4491 21428 4497
rect 21394 4429 21428 4453
rect 21394 4419 21428 4429
rect 21394 4361 21428 4381
rect 21394 4347 21428 4361
rect 21394 4293 21428 4309
rect 21394 4275 21428 4293
rect 21394 4225 21428 4237
rect 21394 4203 21428 4225
rect 21394 4157 21428 4165
rect 21394 4131 21428 4157
rect 21490 5075 21524 5101
rect 21490 5067 21524 5075
rect 21490 5007 21524 5029
rect 21490 4995 21524 5007
rect 21490 4939 21524 4957
rect 21490 4923 21524 4939
rect 21490 4871 21524 4885
rect 21490 4851 21524 4871
rect 21490 4803 21524 4813
rect 21490 4779 21524 4803
rect 21490 4735 21524 4741
rect 21490 4707 21524 4735
rect 21490 4667 21524 4669
rect 21490 4635 21524 4667
rect 21490 4565 21524 4597
rect 21490 4563 21524 4565
rect 21490 4497 21524 4525
rect 21490 4491 21524 4497
rect 21490 4429 21524 4453
rect 21490 4419 21524 4429
rect 21490 4361 21524 4381
rect 21490 4347 21524 4361
rect 21490 4293 21524 4309
rect 21490 4275 21524 4293
rect 21490 4225 21524 4237
rect 21490 4203 21524 4225
rect 21490 4157 21524 4165
rect 21490 4131 21524 4157
rect 21586 5075 21620 5101
rect 21586 5067 21620 5075
rect 21586 5007 21620 5029
rect 21586 4995 21620 5007
rect 21586 4939 21620 4957
rect 21586 4923 21620 4939
rect 21586 4871 21620 4885
rect 21586 4851 21620 4871
rect 21586 4803 21620 4813
rect 21586 4779 21620 4803
rect 21586 4735 21620 4741
rect 21586 4707 21620 4735
rect 21586 4667 21620 4669
rect 21586 4635 21620 4667
rect 21586 4565 21620 4597
rect 21586 4563 21620 4565
rect 21586 4497 21620 4525
rect 21586 4491 21620 4497
rect 21586 4429 21620 4453
rect 21586 4419 21620 4429
rect 21586 4361 21620 4381
rect 21586 4347 21620 4361
rect 21586 4293 21620 4309
rect 21586 4275 21620 4293
rect 21586 4225 21620 4237
rect 21586 4203 21620 4225
rect 21586 4157 21620 4165
rect 21586 4131 21620 4157
rect 21682 5075 21716 5101
rect 21682 5067 21716 5075
rect 21682 5007 21716 5029
rect 21682 4995 21716 5007
rect 21682 4939 21716 4957
rect 21682 4923 21716 4939
rect 21682 4871 21716 4885
rect 21682 4851 21716 4871
rect 21682 4803 21716 4813
rect 21682 4779 21716 4803
rect 21682 4735 21716 4741
rect 21682 4707 21716 4735
rect 21682 4667 21716 4669
rect 21682 4635 21716 4667
rect 21682 4565 21716 4597
rect 21682 4563 21716 4565
rect 21682 4497 21716 4525
rect 21682 4491 21716 4497
rect 21682 4429 21716 4453
rect 21682 4419 21716 4429
rect 21682 4361 21716 4381
rect 21682 4347 21716 4361
rect 21682 4293 21716 4309
rect 21682 4275 21716 4293
rect 21682 4225 21716 4237
rect 21682 4203 21716 4225
rect 21682 4157 21716 4165
rect 21682 4131 21716 4157
rect 21778 5075 21812 5101
rect 21778 5067 21812 5075
rect 21778 5007 21812 5029
rect 21778 4995 21812 5007
rect 21778 4939 21812 4957
rect 21778 4923 21812 4939
rect 21778 4871 21812 4885
rect 21778 4851 21812 4871
rect 21778 4803 21812 4813
rect 21778 4779 21812 4803
rect 21778 4735 21812 4741
rect 21778 4707 21812 4735
rect 21778 4667 21812 4669
rect 21778 4635 21812 4667
rect 21778 4565 21812 4597
rect 21778 4563 21812 4565
rect 21778 4497 21812 4525
rect 21778 4491 21812 4497
rect 21778 4429 21812 4453
rect 21778 4419 21812 4429
rect 21778 4361 21812 4381
rect 21778 4347 21812 4361
rect 21778 4293 21812 4309
rect 21778 4275 21812 4293
rect 21778 4225 21812 4237
rect 21778 4203 21812 4225
rect 21778 4157 21812 4165
rect 21778 4131 21812 4157
rect 21874 5075 21908 5101
rect 21874 5067 21908 5075
rect 21874 5007 21908 5029
rect 21874 4995 21908 5007
rect 21874 4939 21908 4957
rect 21874 4923 21908 4939
rect 21874 4871 21908 4885
rect 21874 4851 21908 4871
rect 21874 4803 21908 4813
rect 21874 4779 21908 4803
rect 21874 4735 21908 4741
rect 21874 4707 21908 4735
rect 21874 4667 21908 4669
rect 21874 4635 21908 4667
rect 21874 4565 21908 4597
rect 21874 4563 21908 4565
rect 21874 4497 21908 4525
rect 21874 4491 21908 4497
rect 21874 4429 21908 4453
rect 21874 4419 21908 4429
rect 21874 4361 21908 4381
rect 21874 4347 21908 4361
rect 21874 4293 21908 4309
rect 21874 4275 21908 4293
rect 21874 4225 21908 4237
rect 21874 4203 21908 4225
rect 21874 4157 21908 4165
rect 21874 4131 21908 4157
rect 21970 5075 22004 5101
rect 21970 5067 22004 5075
rect 21970 5007 22004 5029
rect 21970 4995 22004 5007
rect 21970 4939 22004 4957
rect 21970 4923 22004 4939
rect 21970 4871 22004 4885
rect 21970 4851 22004 4871
rect 21970 4803 22004 4813
rect 21970 4779 22004 4803
rect 21970 4735 22004 4741
rect 21970 4707 22004 4735
rect 21970 4667 22004 4669
rect 21970 4635 22004 4667
rect 21970 4565 22004 4597
rect 21970 4563 22004 4565
rect 21970 4497 22004 4525
rect 21970 4491 22004 4497
rect 21970 4429 22004 4453
rect 21970 4419 22004 4429
rect 21970 4361 22004 4381
rect 21970 4347 22004 4361
rect 21970 4293 22004 4309
rect 21970 4275 22004 4293
rect 21970 4225 22004 4237
rect 21970 4203 22004 4225
rect 21970 4157 22004 4165
rect 21970 4131 22004 4157
rect 22066 5075 22100 5101
rect 22066 5067 22100 5075
rect 22066 5007 22100 5029
rect 22066 4995 22100 5007
rect 22066 4939 22100 4957
rect 22066 4923 22100 4939
rect 22066 4871 22100 4885
rect 22066 4851 22100 4871
rect 22066 4803 22100 4813
rect 22066 4779 22100 4803
rect 22066 4735 22100 4741
rect 22066 4707 22100 4735
rect 22066 4667 22100 4669
rect 22066 4635 22100 4667
rect 22066 4565 22100 4597
rect 22066 4563 22100 4565
rect 22066 4497 22100 4525
rect 22066 4491 22100 4497
rect 22066 4429 22100 4453
rect 22066 4419 22100 4429
rect 22066 4361 22100 4381
rect 22066 4347 22100 4361
rect 22066 4293 22100 4309
rect 22066 4275 22100 4293
rect 22066 4225 22100 4237
rect 22066 4203 22100 4225
rect 22066 4157 22100 4165
rect 22066 4131 22100 4157
rect 22162 5075 22196 5101
rect 22162 5067 22196 5075
rect 22162 5007 22196 5029
rect 22162 4995 22196 5007
rect 22162 4939 22196 4957
rect 22162 4923 22196 4939
rect 22162 4871 22196 4885
rect 22162 4851 22196 4871
rect 22162 4803 22196 4813
rect 22162 4779 22196 4803
rect 22162 4735 22196 4741
rect 22162 4707 22196 4735
rect 22162 4667 22196 4669
rect 22162 4635 22196 4667
rect 22162 4565 22196 4597
rect 22162 4563 22196 4565
rect 22162 4497 22196 4525
rect 22162 4491 22196 4497
rect 22162 4429 22196 4453
rect 22162 4419 22196 4429
rect 22162 4361 22196 4381
rect 22162 4347 22196 4361
rect 22162 4293 22196 4309
rect 22162 4275 22196 4293
rect 22162 4225 22196 4237
rect 22162 4203 22196 4225
rect 22162 4157 22196 4165
rect 22162 4131 22196 4157
rect 22258 5075 22292 5101
rect 22258 5067 22292 5075
rect 22258 5007 22292 5029
rect 22258 4995 22292 5007
rect 22258 4939 22292 4957
rect 22258 4923 22292 4939
rect 22258 4871 22292 4885
rect 22258 4851 22292 4871
rect 22258 4803 22292 4813
rect 22258 4779 22292 4803
rect 22258 4735 22292 4741
rect 22258 4707 22292 4735
rect 22258 4667 22292 4669
rect 22258 4635 22292 4667
rect 22258 4565 22292 4597
rect 22258 4563 22292 4565
rect 22258 4497 22292 4525
rect 22258 4491 22292 4497
rect 22258 4429 22292 4453
rect 22258 4419 22292 4429
rect 22258 4361 22292 4381
rect 22258 4347 22292 4361
rect 22258 4293 22292 4309
rect 22258 4275 22292 4293
rect 22258 4225 22292 4237
rect 22258 4203 22292 4225
rect 22258 4157 22292 4165
rect 22258 4131 22292 4157
rect 23270 5087 23304 5113
rect 23270 5079 23304 5087
rect 23270 5019 23304 5041
rect 23270 5007 23304 5019
rect 23270 4951 23304 4969
rect 23270 4935 23304 4951
rect 23270 4883 23304 4897
rect 23270 4863 23304 4883
rect 23270 4815 23304 4825
rect 23270 4791 23304 4815
rect 23270 4747 23304 4753
rect 23270 4719 23304 4747
rect 23270 4679 23304 4681
rect 23270 4647 23304 4679
rect 23270 4577 23304 4609
rect 23270 4575 23304 4577
rect 23270 4509 23304 4537
rect 23270 4503 23304 4509
rect 23270 4441 23304 4465
rect 23270 4431 23304 4441
rect 23270 4373 23304 4393
rect 23270 4359 23304 4373
rect 23270 4305 23304 4321
rect 23270 4287 23304 4305
rect 23270 4237 23304 4249
rect 23270 4215 23304 4237
rect 23270 4169 23304 4177
rect 23270 4143 23304 4169
rect 23366 5087 23400 5113
rect 23366 5079 23400 5087
rect 23366 5019 23400 5041
rect 23366 5007 23400 5019
rect 23366 4951 23400 4969
rect 23366 4935 23400 4951
rect 23366 4883 23400 4897
rect 23366 4863 23400 4883
rect 23366 4815 23400 4825
rect 23366 4791 23400 4815
rect 23366 4747 23400 4753
rect 23366 4719 23400 4747
rect 23366 4679 23400 4681
rect 23366 4647 23400 4679
rect 23366 4577 23400 4609
rect 23366 4575 23400 4577
rect 23366 4509 23400 4537
rect 23366 4503 23400 4509
rect 23366 4441 23400 4465
rect 23366 4431 23400 4441
rect 23366 4373 23400 4393
rect 23366 4359 23400 4373
rect 23366 4305 23400 4321
rect 23366 4287 23400 4305
rect 23366 4237 23400 4249
rect 23366 4215 23400 4237
rect 23366 4169 23400 4177
rect 23366 4143 23400 4169
rect 23462 5087 23496 5113
rect 23462 5079 23496 5087
rect 23462 5019 23496 5041
rect 23462 5007 23496 5019
rect 23462 4951 23496 4969
rect 23462 4935 23496 4951
rect 23462 4883 23496 4897
rect 23462 4863 23496 4883
rect 23462 4815 23496 4825
rect 23462 4791 23496 4815
rect 23462 4747 23496 4753
rect 23462 4719 23496 4747
rect 23462 4679 23496 4681
rect 23462 4647 23496 4679
rect 23462 4577 23496 4609
rect 23462 4575 23496 4577
rect 23462 4509 23496 4537
rect 23462 4503 23496 4509
rect 23462 4441 23496 4465
rect 23462 4431 23496 4441
rect 23462 4373 23496 4393
rect 23462 4359 23496 4373
rect 23462 4305 23496 4321
rect 23462 4287 23496 4305
rect 23462 4237 23496 4249
rect 23462 4215 23496 4237
rect 23462 4169 23496 4177
rect 23462 4143 23496 4169
rect 23558 5087 23592 5113
rect 23558 5079 23592 5087
rect 23558 5019 23592 5041
rect 23558 5007 23592 5019
rect 23558 4951 23592 4969
rect 23558 4935 23592 4951
rect 23558 4883 23592 4897
rect 23558 4863 23592 4883
rect 23558 4815 23592 4825
rect 23558 4791 23592 4815
rect 23558 4747 23592 4753
rect 23558 4719 23592 4747
rect 23558 4679 23592 4681
rect 23558 4647 23592 4679
rect 23558 4577 23592 4609
rect 23558 4575 23592 4577
rect 23558 4509 23592 4537
rect 23558 4503 23592 4509
rect 23558 4441 23592 4465
rect 23558 4431 23592 4441
rect 23558 4373 23592 4393
rect 23558 4359 23592 4373
rect 23558 4305 23592 4321
rect 23558 4287 23592 4305
rect 23558 4237 23592 4249
rect 23558 4215 23592 4237
rect 23558 4169 23592 4177
rect 23558 4143 23592 4169
rect 23654 5087 23688 5113
rect 23654 5079 23688 5087
rect 23654 5019 23688 5041
rect 23654 5007 23688 5019
rect 23654 4951 23688 4969
rect 23654 4935 23688 4951
rect 23654 4883 23688 4897
rect 23654 4863 23688 4883
rect 23654 4815 23688 4825
rect 23654 4791 23688 4815
rect 23654 4747 23688 4753
rect 23654 4719 23688 4747
rect 23654 4679 23688 4681
rect 23654 4647 23688 4679
rect 23654 4577 23688 4609
rect 23654 4575 23688 4577
rect 23654 4509 23688 4537
rect 23654 4503 23688 4509
rect 23654 4441 23688 4465
rect 23654 4431 23688 4441
rect 23654 4373 23688 4393
rect 23654 4359 23688 4373
rect 23654 4305 23688 4321
rect 23654 4287 23688 4305
rect 23654 4237 23688 4249
rect 23654 4215 23688 4237
rect 23654 4169 23688 4177
rect 23654 4143 23688 4169
rect 23750 5087 23784 5113
rect 23750 5079 23784 5087
rect 23750 5019 23784 5041
rect 23750 5007 23784 5019
rect 23750 4951 23784 4969
rect 23750 4935 23784 4951
rect 23750 4883 23784 4897
rect 23750 4863 23784 4883
rect 23750 4815 23784 4825
rect 23750 4791 23784 4815
rect 23750 4747 23784 4753
rect 23750 4719 23784 4747
rect 23750 4679 23784 4681
rect 23750 4647 23784 4679
rect 23750 4577 23784 4609
rect 23750 4575 23784 4577
rect 23750 4509 23784 4537
rect 23750 4503 23784 4509
rect 23750 4441 23784 4465
rect 23750 4431 23784 4441
rect 23750 4373 23784 4393
rect 23750 4359 23784 4373
rect 23750 4305 23784 4321
rect 23750 4287 23784 4305
rect 23750 4237 23784 4249
rect 23750 4215 23784 4237
rect 23750 4169 23784 4177
rect 23750 4143 23784 4169
rect 23958 5085 23992 5111
rect 23958 5077 23992 5085
rect 23958 5017 23992 5039
rect 23958 5005 23992 5017
rect 23958 4949 23992 4967
rect 23958 4933 23992 4949
rect 23958 4881 23992 4895
rect 23958 4861 23992 4881
rect 23958 4813 23992 4823
rect 23958 4789 23992 4813
rect 23958 4745 23992 4751
rect 23958 4717 23992 4745
rect 23958 4677 23992 4679
rect 23958 4645 23992 4677
rect 23958 4575 23992 4607
rect 23958 4573 23992 4575
rect 23958 4507 23992 4535
rect 23958 4501 23992 4507
rect 23958 4439 23992 4463
rect 23958 4429 23992 4439
rect 23958 4371 23992 4391
rect 23958 4357 23992 4371
rect 23958 4303 23992 4319
rect 23958 4285 23992 4303
rect 23958 4235 23992 4247
rect 23958 4213 23992 4235
rect 23958 4167 23992 4175
rect 23958 4141 23992 4167
rect 24054 5085 24088 5111
rect 24054 5077 24088 5085
rect 24054 5017 24088 5039
rect 24054 5005 24088 5017
rect 24054 4949 24088 4967
rect 24054 4933 24088 4949
rect 24054 4881 24088 4895
rect 24054 4861 24088 4881
rect 24054 4813 24088 4823
rect 24054 4789 24088 4813
rect 24054 4745 24088 4751
rect 24054 4717 24088 4745
rect 24054 4677 24088 4679
rect 24054 4645 24088 4677
rect 24054 4575 24088 4607
rect 24054 4573 24088 4575
rect 24054 4507 24088 4535
rect 24054 4501 24088 4507
rect 24054 4439 24088 4463
rect 24054 4429 24088 4439
rect 24054 4371 24088 4391
rect 24054 4357 24088 4371
rect 24054 4303 24088 4319
rect 24054 4285 24088 4303
rect 24054 4235 24088 4247
rect 24054 4213 24088 4235
rect 24054 4167 24088 4175
rect 24054 4141 24088 4167
rect 24150 5085 24184 5111
rect 24150 5077 24184 5085
rect 24150 5017 24184 5039
rect 24150 5005 24184 5017
rect 24150 4949 24184 4967
rect 24150 4933 24184 4949
rect 24150 4881 24184 4895
rect 24150 4861 24184 4881
rect 24150 4813 24184 4823
rect 24150 4789 24184 4813
rect 24150 4745 24184 4751
rect 24150 4717 24184 4745
rect 24150 4677 24184 4679
rect 24150 4645 24184 4677
rect 24150 4575 24184 4607
rect 24150 4573 24184 4575
rect 24150 4507 24184 4535
rect 24150 4501 24184 4507
rect 24150 4439 24184 4463
rect 24150 4429 24184 4439
rect 24150 4371 24184 4391
rect 24150 4357 24184 4371
rect 24150 4303 24184 4319
rect 24150 4285 24184 4303
rect 24150 4235 24184 4247
rect 24150 4213 24184 4235
rect 24150 4167 24184 4175
rect 24150 4141 24184 4167
rect 24246 5085 24280 5111
rect 24246 5077 24280 5085
rect 24246 5017 24280 5039
rect 24246 5005 24280 5017
rect 24246 4949 24280 4967
rect 24246 4933 24280 4949
rect 24246 4881 24280 4895
rect 24246 4861 24280 4881
rect 24246 4813 24280 4823
rect 24246 4789 24280 4813
rect 24246 4745 24280 4751
rect 24246 4717 24280 4745
rect 24246 4677 24280 4679
rect 24246 4645 24280 4677
rect 24246 4575 24280 4607
rect 24246 4573 24280 4575
rect 24246 4507 24280 4535
rect 24246 4501 24280 4507
rect 24246 4439 24280 4463
rect 24246 4429 24280 4439
rect 24246 4371 24280 4391
rect 24246 4357 24280 4371
rect 24246 4303 24280 4319
rect 24246 4285 24280 4303
rect 24246 4235 24280 4247
rect 24246 4213 24280 4235
rect 24246 4167 24280 4175
rect 24246 4141 24280 4167
rect 24342 5085 24376 5111
rect 24342 5077 24376 5085
rect 24342 5017 24376 5039
rect 24342 5005 24376 5017
rect 24342 4949 24376 4967
rect 24342 4933 24376 4949
rect 24342 4881 24376 4895
rect 24342 4861 24376 4881
rect 24342 4813 24376 4823
rect 24342 4789 24376 4813
rect 24342 4745 24376 4751
rect 24342 4717 24376 4745
rect 24342 4677 24376 4679
rect 24342 4645 24376 4677
rect 24342 4575 24376 4607
rect 24342 4573 24376 4575
rect 24342 4507 24376 4535
rect 24342 4501 24376 4507
rect 24342 4439 24376 4463
rect 24342 4429 24376 4439
rect 24342 4371 24376 4391
rect 24342 4357 24376 4371
rect 24342 4303 24376 4319
rect 24342 4285 24376 4303
rect 24342 4235 24376 4247
rect 24342 4213 24376 4235
rect 24342 4167 24376 4175
rect 24342 4141 24376 4167
rect 24438 5085 24472 5111
rect 24438 5077 24472 5085
rect 24438 5017 24472 5039
rect 24438 5005 24472 5017
rect 24438 4949 24472 4967
rect 24438 4933 24472 4949
rect 24438 4881 24472 4895
rect 24438 4861 24472 4881
rect 24438 4813 24472 4823
rect 24438 4789 24472 4813
rect 24438 4745 24472 4751
rect 24438 4717 24472 4745
rect 24438 4677 24472 4679
rect 24438 4645 24472 4677
rect 24438 4575 24472 4607
rect 24438 4573 24472 4575
rect 24438 4507 24472 4535
rect 24438 4501 24472 4507
rect 24438 4439 24472 4463
rect 24438 4429 24472 4439
rect 24438 4371 24472 4391
rect 24438 4357 24472 4371
rect 24438 4303 24472 4319
rect 24438 4285 24472 4303
rect 24438 4235 24472 4247
rect 24438 4213 24472 4235
rect 24438 4167 24472 4175
rect 24438 4141 24472 4167
rect 24534 5085 24568 5111
rect 24534 5077 24568 5085
rect 24534 5017 24568 5039
rect 24534 5005 24568 5017
rect 24534 4949 24568 4967
rect 24534 4933 24568 4949
rect 24534 4881 24568 4895
rect 24534 4861 24568 4881
rect 24534 4813 24568 4823
rect 24534 4789 24568 4813
rect 24534 4745 24568 4751
rect 24534 4717 24568 4745
rect 24534 4677 24568 4679
rect 24534 4645 24568 4677
rect 24534 4575 24568 4607
rect 24534 4573 24568 4575
rect 24534 4507 24568 4535
rect 24534 4501 24568 4507
rect 24534 4439 24568 4463
rect 24534 4429 24568 4439
rect 24534 4371 24568 4391
rect 24534 4357 24568 4371
rect 24534 4303 24568 4319
rect 24534 4285 24568 4303
rect 24534 4235 24568 4247
rect 24534 4213 24568 4235
rect 24534 4167 24568 4175
rect 24534 4141 24568 4167
rect 24630 5085 24664 5111
rect 24630 5077 24664 5085
rect 24630 5017 24664 5039
rect 24630 5005 24664 5017
rect 24630 4949 24664 4967
rect 24630 4933 24664 4949
rect 24630 4881 24664 4895
rect 24630 4861 24664 4881
rect 24630 4813 24664 4823
rect 24630 4789 24664 4813
rect 24630 4745 24664 4751
rect 24630 4717 24664 4745
rect 24630 4677 24664 4679
rect 24630 4645 24664 4677
rect 24630 4575 24664 4607
rect 24630 4573 24664 4575
rect 24630 4507 24664 4535
rect 24630 4501 24664 4507
rect 24630 4439 24664 4463
rect 24630 4429 24664 4439
rect 24630 4371 24664 4391
rect 24630 4357 24664 4371
rect 24630 4303 24664 4319
rect 24630 4285 24664 4303
rect 24630 4235 24664 4247
rect 24630 4213 24664 4235
rect 24630 4167 24664 4175
rect 24630 4141 24664 4167
rect 24726 5085 24760 5111
rect 24726 5077 24760 5085
rect 24726 5017 24760 5039
rect 24726 5005 24760 5017
rect 24726 4949 24760 4967
rect 24726 4933 24760 4949
rect 24726 4881 24760 4895
rect 24726 4861 24760 4881
rect 24726 4813 24760 4823
rect 24726 4789 24760 4813
rect 24726 4745 24760 4751
rect 24726 4717 24760 4745
rect 24726 4677 24760 4679
rect 24726 4645 24760 4677
rect 24726 4575 24760 4607
rect 24726 4573 24760 4575
rect 24726 4507 24760 4535
rect 24726 4501 24760 4507
rect 24726 4439 24760 4463
rect 24726 4429 24760 4439
rect 24726 4371 24760 4391
rect 24726 4357 24760 4371
rect 24726 4303 24760 4319
rect 24726 4285 24760 4303
rect 24726 4235 24760 4247
rect 24726 4213 24760 4235
rect 24726 4167 24760 4175
rect 24726 4141 24760 4167
rect 24822 5085 24856 5111
rect 24822 5077 24856 5085
rect 24822 5017 24856 5039
rect 24822 5005 24856 5017
rect 24822 4949 24856 4967
rect 24822 4933 24856 4949
rect 24822 4881 24856 4895
rect 24822 4861 24856 4881
rect 24822 4813 24856 4823
rect 24822 4789 24856 4813
rect 24822 4745 24856 4751
rect 24822 4717 24856 4745
rect 24822 4677 24856 4679
rect 24822 4645 24856 4677
rect 24822 4575 24856 4607
rect 24822 4573 24856 4575
rect 24822 4507 24856 4535
rect 24822 4501 24856 4507
rect 24822 4439 24856 4463
rect 24822 4429 24856 4439
rect 24822 4371 24856 4391
rect 24822 4357 24856 4371
rect 24822 4303 24856 4319
rect 24822 4285 24856 4303
rect 24822 4235 24856 4247
rect 24822 4213 24856 4235
rect 24822 4167 24856 4175
rect 24822 4141 24856 4167
rect 24918 5085 24952 5111
rect 24918 5077 24952 5085
rect 24918 5017 24952 5039
rect 24918 5005 24952 5017
rect 24918 4949 24952 4967
rect 24918 4933 24952 4949
rect 24918 4881 24952 4895
rect 24918 4861 24952 4881
rect 24918 4813 24952 4823
rect 24918 4789 24952 4813
rect 24918 4745 24952 4751
rect 24918 4717 24952 4745
rect 24918 4677 24952 4679
rect 24918 4645 24952 4677
rect 24918 4575 24952 4607
rect 24918 4573 24952 4575
rect 24918 4507 24952 4535
rect 24918 4501 24952 4507
rect 24918 4439 24952 4463
rect 24918 4429 24952 4439
rect 24918 4371 24952 4391
rect 24918 4357 24952 4371
rect 24918 4303 24952 4319
rect 24918 4285 24952 4303
rect 24918 4235 24952 4247
rect 24918 4213 24952 4235
rect 24918 4167 24952 4175
rect 24918 4141 24952 4167
rect 25162 5079 25196 5105
rect 25162 5071 25196 5079
rect 25162 5011 25196 5033
rect 25162 4999 25196 5011
rect 25162 4943 25196 4961
rect 25162 4927 25196 4943
rect 25162 4875 25196 4889
rect 25162 4855 25196 4875
rect 25162 4807 25196 4817
rect 25162 4783 25196 4807
rect 25162 4739 25196 4745
rect 25162 4711 25196 4739
rect 25162 4671 25196 4673
rect 25162 4639 25196 4671
rect 25162 4569 25196 4601
rect 25162 4567 25196 4569
rect 25162 4501 25196 4529
rect 25162 4495 25196 4501
rect 25162 4433 25196 4457
rect 25162 4423 25196 4433
rect 25162 4365 25196 4385
rect 25162 4351 25196 4365
rect 25162 4297 25196 4313
rect 25162 4279 25196 4297
rect 25162 4229 25196 4241
rect 25162 4207 25196 4229
rect 25162 4161 25196 4169
rect 25162 4135 25196 4161
rect 25258 5079 25292 5105
rect 25258 5071 25292 5079
rect 25258 5011 25292 5033
rect 25258 4999 25292 5011
rect 25258 4943 25292 4961
rect 25258 4927 25292 4943
rect 25258 4875 25292 4889
rect 25258 4855 25292 4875
rect 25258 4807 25292 4817
rect 25258 4783 25292 4807
rect 25258 4739 25292 4745
rect 25258 4711 25292 4739
rect 25258 4671 25292 4673
rect 25258 4639 25292 4671
rect 25258 4569 25292 4601
rect 25258 4567 25292 4569
rect 25258 4501 25292 4529
rect 25258 4495 25292 4501
rect 25258 4433 25292 4457
rect 25258 4423 25292 4433
rect 25258 4365 25292 4385
rect 25258 4351 25292 4365
rect 25258 4297 25292 4313
rect 25258 4279 25292 4297
rect 25258 4229 25292 4241
rect 25258 4207 25292 4229
rect 25258 4161 25292 4169
rect 25258 4135 25292 4161
rect 18722 3921 18756 3955
rect 17790 3785 17824 3819
rect 17522 3702 17556 3736
rect 20386 3915 20420 3949
rect 19443 3772 19477 3806
rect 18720 3658 18754 3692
rect -4814 3575 -4780 3587
rect -4814 3553 -4780 3575
rect -4814 3507 -4780 3515
rect -4814 3481 -4780 3507
rect 16686 3493 16720 3519
rect 16686 3485 16720 3493
rect -1590 3394 -1556 3428
rect 16686 3425 16720 3447
rect 16686 3413 16720 3425
rect -8418 3251 -8384 3285
rect -9678 3106 -9644 3140
rect -11328 3010 -11294 3044
rect -13170 2817 -13136 2843
rect -13170 2809 -13136 2817
rect -13170 2749 -13136 2771
rect -13170 2737 -13136 2749
rect -13170 2681 -13136 2699
rect -13170 2665 -13136 2681
rect -13170 2613 -13136 2627
rect -13170 2593 -13136 2613
rect -13170 2545 -13136 2555
rect -13170 2521 -13136 2545
rect -13170 2477 -13136 2483
rect -13170 2449 -13136 2477
rect -13170 2409 -13136 2411
rect -13170 2377 -13136 2409
rect -13170 2307 -13136 2339
rect -13170 2305 -13136 2307
rect -13170 2239 -13136 2267
rect -13170 2233 -13136 2239
rect -13170 2171 -13136 2195
rect -13170 2161 -13136 2171
rect -13170 2103 -13136 2123
rect -13170 2089 -13136 2103
rect -13170 2035 -13136 2051
rect -13170 2017 -13136 2035
rect -13170 1967 -13136 1979
rect -13170 1945 -13136 1967
rect -13170 1899 -13136 1907
rect -13170 1873 -13136 1899
rect -13074 2817 -13040 2843
rect -13074 2809 -13040 2817
rect -13074 2749 -13040 2771
rect -13074 2737 -13040 2749
rect -13074 2681 -13040 2699
rect -13074 2665 -13040 2681
rect -13074 2613 -13040 2627
rect -13074 2593 -13040 2613
rect -13074 2545 -13040 2555
rect -13074 2521 -13040 2545
rect -13074 2477 -13040 2483
rect -13074 2449 -13040 2477
rect -13074 2409 -13040 2411
rect -13074 2377 -13040 2409
rect -13074 2307 -13040 2339
rect -13074 2305 -13040 2307
rect -13074 2239 -13040 2267
rect -13074 2233 -13040 2239
rect -13074 2171 -13040 2195
rect -13074 2161 -13040 2171
rect -13074 2103 -13040 2123
rect -13074 2089 -13040 2103
rect -13074 2035 -13040 2051
rect -13074 2017 -13040 2035
rect -13074 1967 -13040 1979
rect -13074 1945 -13040 1967
rect -13074 1899 -13040 1907
rect -13074 1873 -13040 1899
rect -12836 2821 -12802 2847
rect -12836 2813 -12802 2821
rect -12836 2753 -12802 2775
rect -12836 2741 -12802 2753
rect -12836 2685 -12802 2703
rect -12836 2669 -12802 2685
rect -12836 2617 -12802 2631
rect -12836 2597 -12802 2617
rect -12836 2549 -12802 2559
rect -12836 2525 -12802 2549
rect -12836 2481 -12802 2487
rect -12836 2453 -12802 2481
rect -12836 2413 -12802 2415
rect -12836 2381 -12802 2413
rect -12836 2311 -12802 2343
rect -12836 2309 -12802 2311
rect -12836 2243 -12802 2271
rect -12836 2237 -12802 2243
rect -12836 2175 -12802 2199
rect -12836 2165 -12802 2175
rect -12836 2107 -12802 2127
rect -12836 2093 -12802 2107
rect -12836 2039 -12802 2055
rect -12836 2021 -12802 2039
rect -12836 1971 -12802 1983
rect -12836 1949 -12802 1971
rect -12836 1903 -12802 1911
rect -12836 1877 -12802 1903
rect -12740 2821 -12706 2847
rect -12740 2813 -12706 2821
rect -12740 2753 -12706 2775
rect -12740 2741 -12706 2753
rect -12740 2685 -12706 2703
rect -12740 2669 -12706 2685
rect -12740 2617 -12706 2631
rect -12740 2597 -12706 2617
rect -12740 2549 -12706 2559
rect -12740 2525 -12706 2549
rect -12740 2481 -12706 2487
rect -12740 2453 -12706 2481
rect -12740 2413 -12706 2415
rect -12740 2381 -12706 2413
rect -12740 2311 -12706 2343
rect -12740 2309 -12706 2311
rect -12740 2243 -12706 2271
rect -12740 2237 -12706 2243
rect -12740 2175 -12706 2199
rect -12740 2165 -12706 2175
rect -12740 2107 -12706 2127
rect -12740 2093 -12706 2107
rect -12740 2039 -12706 2055
rect -12740 2021 -12706 2039
rect -12740 1971 -12706 1983
rect -12740 1949 -12706 1971
rect -12740 1903 -12706 1911
rect -12740 1877 -12706 1903
rect -12644 2821 -12610 2847
rect -12644 2813 -12610 2821
rect -12644 2753 -12610 2775
rect -12644 2741 -12610 2753
rect -12644 2685 -12610 2703
rect -12644 2669 -12610 2685
rect -12644 2617 -12610 2631
rect -12644 2597 -12610 2617
rect -12644 2549 -12610 2559
rect -12644 2525 -12610 2549
rect -12644 2481 -12610 2487
rect -12644 2453 -12610 2481
rect -12644 2413 -12610 2415
rect -12644 2381 -12610 2413
rect -12644 2311 -12610 2343
rect -12644 2309 -12610 2311
rect -12644 2243 -12610 2271
rect -12644 2237 -12610 2243
rect -12644 2175 -12610 2199
rect -12644 2165 -12610 2175
rect -12644 2107 -12610 2127
rect -12644 2093 -12610 2107
rect -12644 2039 -12610 2055
rect -12644 2021 -12610 2039
rect -12644 1971 -12610 1983
rect -12644 1949 -12610 1971
rect -12644 1903 -12610 1911
rect -12644 1877 -12610 1903
rect -12548 2821 -12514 2847
rect -12548 2813 -12514 2821
rect -12548 2753 -12514 2775
rect -12548 2741 -12514 2753
rect -12548 2685 -12514 2703
rect -12548 2669 -12514 2685
rect -12548 2617 -12514 2631
rect -12548 2597 -12514 2617
rect -12548 2549 -12514 2559
rect -12548 2525 -12514 2549
rect -12548 2481 -12514 2487
rect -12548 2453 -12514 2481
rect -12548 2413 -12514 2415
rect -12548 2381 -12514 2413
rect -12548 2311 -12514 2343
rect -12548 2309 -12514 2311
rect -12548 2243 -12514 2271
rect -12548 2237 -12514 2243
rect -12548 2175 -12514 2199
rect -12548 2165 -12514 2175
rect -12548 2107 -12514 2127
rect -12548 2093 -12514 2107
rect -12548 2039 -12514 2055
rect -12548 2021 -12514 2039
rect -12548 1971 -12514 1983
rect -12548 1949 -12514 1971
rect -12548 1903 -12514 1911
rect -12548 1877 -12514 1903
rect -12452 2821 -12418 2847
rect -12452 2813 -12418 2821
rect -12452 2753 -12418 2775
rect -12452 2741 -12418 2753
rect -12452 2685 -12418 2703
rect -12452 2669 -12418 2685
rect -12452 2617 -12418 2631
rect -12452 2597 -12418 2617
rect -12452 2549 -12418 2559
rect -12452 2525 -12418 2549
rect -12452 2481 -12418 2487
rect -12452 2453 -12418 2481
rect -12452 2413 -12418 2415
rect -12452 2381 -12418 2413
rect -12452 2311 -12418 2343
rect -12452 2309 -12418 2311
rect -12452 2243 -12418 2271
rect -12452 2237 -12418 2243
rect -12452 2175 -12418 2199
rect -12452 2165 -12418 2175
rect -12452 2107 -12418 2127
rect -12452 2093 -12418 2107
rect -12452 2039 -12418 2055
rect -12452 2021 -12418 2039
rect -12452 1971 -12418 1983
rect -12452 1949 -12418 1971
rect -12452 1903 -12418 1911
rect -12452 1877 -12418 1903
rect -12356 2821 -12322 2847
rect -12356 2813 -12322 2821
rect -12356 2753 -12322 2775
rect -12356 2741 -12322 2753
rect -12356 2685 -12322 2703
rect -12356 2669 -12322 2685
rect -12356 2617 -12322 2631
rect -12356 2597 -12322 2617
rect -12356 2549 -12322 2559
rect -12356 2525 -12322 2549
rect -12356 2481 -12322 2487
rect -12356 2453 -12322 2481
rect -12356 2413 -12322 2415
rect -12356 2381 -12322 2413
rect -12356 2311 -12322 2343
rect -12356 2309 -12322 2311
rect -12356 2243 -12322 2271
rect -12356 2237 -12322 2243
rect -12356 2175 -12322 2199
rect -12356 2165 -12322 2175
rect -12356 2107 -12322 2127
rect -12356 2093 -12322 2107
rect -12356 2039 -12322 2055
rect -12356 2021 -12322 2039
rect -12356 1971 -12322 1983
rect -12356 1949 -12322 1971
rect -12356 1903 -12322 1911
rect -12356 1877 -12322 1903
rect -12260 2821 -12226 2847
rect -12260 2813 -12226 2821
rect -12260 2753 -12226 2775
rect -12260 2741 -12226 2753
rect -12260 2685 -12226 2703
rect -12260 2669 -12226 2685
rect -12260 2617 -12226 2631
rect -12260 2597 -12226 2617
rect -12260 2549 -12226 2559
rect -12260 2525 -12226 2549
rect -12260 2481 -12226 2487
rect -12260 2453 -12226 2481
rect -12260 2413 -12226 2415
rect -12260 2381 -12226 2413
rect -12260 2311 -12226 2343
rect -12260 2309 -12226 2311
rect -12260 2243 -12226 2271
rect -12260 2237 -12226 2243
rect -12260 2175 -12226 2199
rect -12260 2165 -12226 2175
rect -12260 2107 -12226 2127
rect -12260 2093 -12226 2107
rect -12260 2039 -12226 2055
rect -12260 2021 -12226 2039
rect -12260 1971 -12226 1983
rect -12260 1949 -12226 1971
rect -12260 1903 -12226 1911
rect -12260 1877 -12226 1903
rect -12164 2821 -12130 2847
rect -12164 2813 -12130 2821
rect -12164 2753 -12130 2775
rect -12164 2741 -12130 2753
rect -12164 2685 -12130 2703
rect -12164 2669 -12130 2685
rect -12164 2617 -12130 2631
rect -12164 2597 -12130 2617
rect -12164 2549 -12130 2559
rect -12164 2525 -12130 2549
rect -12164 2481 -12130 2487
rect -12164 2453 -12130 2481
rect -12164 2413 -12130 2415
rect -12164 2381 -12130 2413
rect -12164 2311 -12130 2343
rect -12164 2309 -12130 2311
rect -12164 2243 -12130 2271
rect -12164 2237 -12130 2243
rect -12164 2175 -12130 2199
rect -12164 2165 -12130 2175
rect -12164 2107 -12130 2127
rect -12164 2093 -12130 2107
rect -12164 2039 -12130 2055
rect -12164 2021 -12130 2039
rect -12164 1971 -12130 1983
rect -12164 1949 -12130 1971
rect -12164 1903 -12130 1911
rect -12164 1877 -12130 1903
rect -12068 2821 -12034 2847
rect -12068 2813 -12034 2821
rect -12068 2753 -12034 2775
rect -12068 2741 -12034 2753
rect -12068 2685 -12034 2703
rect -12068 2669 -12034 2685
rect -12068 2617 -12034 2631
rect -12068 2597 -12034 2617
rect -12068 2549 -12034 2559
rect -12068 2525 -12034 2549
rect -12068 2481 -12034 2487
rect -12068 2453 -12034 2481
rect -12068 2413 -12034 2415
rect -12068 2381 -12034 2413
rect -12068 2311 -12034 2343
rect -12068 2309 -12034 2311
rect -12068 2243 -12034 2271
rect -12068 2237 -12034 2243
rect -12068 2175 -12034 2199
rect -12068 2165 -12034 2175
rect -12068 2107 -12034 2127
rect -12068 2093 -12034 2107
rect -12068 2039 -12034 2055
rect -12068 2021 -12034 2039
rect -12068 1971 -12034 1983
rect -12068 1949 -12034 1971
rect -12068 1903 -12034 1911
rect -12068 1877 -12034 1903
rect -6754 3257 -6720 3291
rect -7475 3108 -7441 3142
rect -8420 2992 -8386 3026
rect -5550 3263 -5516 3297
rect -5822 3121 -5788 3155
rect -6752 2994 -6718 3028
rect 16686 3357 16720 3375
rect 16686 3341 16720 3357
rect -1110 3290 -1076 3324
rect -4862 3245 -4828 3279
rect -5006 3123 -4972 3157
rect -5554 3038 -5520 3072
rect -11972 2821 -11938 2847
rect -11972 2813 -11938 2821
rect -11972 2753 -11938 2775
rect -11972 2741 -11938 2753
rect -11972 2685 -11938 2703
rect -11972 2669 -11938 2685
rect -11972 2617 -11938 2631
rect -11972 2597 -11938 2617
rect -11972 2549 -11938 2559
rect -11972 2525 -11938 2549
rect -11972 2481 -11938 2487
rect -11972 2453 -11938 2481
rect -11972 2413 -11938 2415
rect -11972 2381 -11938 2413
rect -11972 2311 -11938 2343
rect -11972 2309 -11938 2311
rect -11972 2243 -11938 2271
rect -11972 2237 -11938 2243
rect -11972 2175 -11938 2199
rect -11972 2165 -11938 2175
rect -11972 2107 -11938 2127
rect -11972 2093 -11938 2107
rect -11972 2039 -11938 2055
rect -11972 2021 -11938 2039
rect -11972 1971 -11938 1983
rect -11972 1949 -11938 1971
rect -11972 1903 -11938 1911
rect -11972 1877 -11938 1903
rect -11876 2821 -11842 2847
rect -11876 2813 -11842 2821
rect -11876 2753 -11842 2775
rect -11876 2741 -11842 2753
rect -11876 2685 -11842 2703
rect -11876 2669 -11842 2685
rect -11876 2617 -11842 2631
rect -11876 2597 -11842 2617
rect -11876 2549 -11842 2559
rect -11876 2525 -11842 2549
rect -11876 2481 -11842 2487
rect -11876 2453 -11842 2481
rect -11876 2413 -11842 2415
rect -11876 2381 -11842 2413
rect -11876 2311 -11842 2343
rect -11876 2309 -11842 2311
rect -11876 2243 -11842 2271
rect -11876 2237 -11842 2243
rect -11876 2175 -11842 2199
rect -11876 2165 -11842 2175
rect -11876 2107 -11842 2127
rect -11876 2093 -11842 2107
rect -11876 2039 -11842 2055
rect -11876 2021 -11842 2039
rect -11876 1971 -11842 1983
rect -11876 1949 -11842 1971
rect -11876 1903 -11842 1911
rect -11876 1877 -11842 1903
rect -11664 2831 -11630 2857
rect -11664 2823 -11630 2831
rect -11664 2763 -11630 2785
rect -11664 2751 -11630 2763
rect -11664 2695 -11630 2713
rect -11664 2679 -11630 2695
rect -11664 2627 -11630 2641
rect -11664 2607 -11630 2627
rect -11664 2559 -11630 2569
rect -11664 2535 -11630 2559
rect -11664 2491 -11630 2497
rect -11664 2463 -11630 2491
rect -11664 2423 -11630 2425
rect -11664 2391 -11630 2423
rect -11664 2321 -11630 2353
rect -11664 2319 -11630 2321
rect -11664 2253 -11630 2281
rect -11664 2247 -11630 2253
rect -11664 2185 -11630 2209
rect -11664 2175 -11630 2185
rect -11664 2117 -11630 2137
rect -11664 2103 -11630 2117
rect -11664 2049 -11630 2065
rect -11664 2031 -11630 2049
rect -11664 1981 -11630 1993
rect -11664 1959 -11630 1981
rect -11664 1913 -11630 1921
rect -11664 1887 -11630 1913
rect -11568 2831 -11534 2857
rect -11568 2823 -11534 2831
rect -11568 2763 -11534 2785
rect -11568 2751 -11534 2763
rect -11568 2695 -11534 2713
rect -11568 2679 -11534 2695
rect -11568 2627 -11534 2641
rect -11568 2607 -11534 2627
rect -11568 2559 -11534 2569
rect -11568 2535 -11534 2559
rect -11568 2491 -11534 2497
rect -11568 2463 -11534 2491
rect -11568 2423 -11534 2425
rect -11568 2391 -11534 2423
rect -11568 2321 -11534 2353
rect -11568 2319 -11534 2321
rect -11568 2253 -11534 2281
rect -11568 2247 -11534 2253
rect -11568 2185 -11534 2209
rect -11568 2175 -11534 2185
rect -11568 2117 -11534 2137
rect -11568 2103 -11534 2117
rect -11568 2049 -11534 2065
rect -11568 2031 -11534 2049
rect -11568 1981 -11534 1993
rect -11568 1959 -11534 1981
rect -11568 1913 -11534 1921
rect -11568 1887 -11534 1913
rect -11472 2831 -11438 2857
rect -11472 2823 -11438 2831
rect -11472 2763 -11438 2785
rect -11472 2751 -11438 2763
rect -11472 2695 -11438 2713
rect -11472 2679 -11438 2695
rect -11472 2627 -11438 2641
rect -11472 2607 -11438 2627
rect -11472 2559 -11438 2569
rect -11472 2535 -11438 2559
rect -11472 2491 -11438 2497
rect -11472 2463 -11438 2491
rect -11472 2423 -11438 2425
rect -11472 2391 -11438 2423
rect -11472 2321 -11438 2353
rect -11472 2319 -11438 2321
rect -11472 2253 -11438 2281
rect -11472 2247 -11438 2253
rect -11472 2185 -11438 2209
rect -11472 2175 -11438 2185
rect -11472 2117 -11438 2137
rect -11472 2103 -11438 2117
rect -11472 2049 -11438 2065
rect -11472 2031 -11438 2049
rect -11472 1981 -11438 1993
rect -11472 1959 -11438 1981
rect -11472 1913 -11438 1921
rect -11472 1887 -11438 1913
rect -11376 2831 -11342 2857
rect -11376 2823 -11342 2831
rect -11376 2763 -11342 2785
rect -11376 2751 -11342 2763
rect -11376 2695 -11342 2713
rect -11376 2679 -11342 2695
rect -11376 2627 -11342 2641
rect -11376 2607 -11342 2627
rect -11376 2559 -11342 2569
rect -11376 2535 -11342 2559
rect -11376 2491 -11342 2497
rect -11376 2463 -11342 2491
rect -11376 2423 -11342 2425
rect -11376 2391 -11342 2423
rect -11376 2321 -11342 2353
rect -11376 2319 -11342 2321
rect -11376 2253 -11342 2281
rect -11376 2247 -11342 2253
rect -11376 2185 -11342 2209
rect -11376 2175 -11342 2185
rect -11376 2117 -11342 2137
rect -11376 2103 -11342 2117
rect -11376 2049 -11342 2065
rect -11376 2031 -11342 2049
rect -11376 1981 -11342 1993
rect -11376 1959 -11342 1981
rect -11376 1913 -11342 1921
rect -11376 1887 -11342 1913
rect -11280 2831 -11246 2857
rect -11280 2823 -11246 2831
rect -11280 2763 -11246 2785
rect -11280 2751 -11246 2763
rect -11280 2695 -11246 2713
rect -11280 2679 -11246 2695
rect -11280 2627 -11246 2641
rect -11280 2607 -11246 2627
rect -11280 2559 -11246 2569
rect -11280 2535 -11246 2559
rect -11280 2491 -11246 2497
rect -11280 2463 -11246 2491
rect -11280 2423 -11246 2425
rect -11280 2391 -11246 2423
rect -11280 2321 -11246 2353
rect -11280 2319 -11246 2321
rect -11280 2253 -11246 2281
rect -11280 2247 -11246 2253
rect -11280 2185 -11246 2209
rect -11280 2175 -11246 2185
rect -11280 2117 -11246 2137
rect -11280 2103 -11246 2117
rect -11280 2049 -11246 2065
rect -11280 2031 -11246 2049
rect -11280 1981 -11246 1993
rect -11280 1959 -11246 1981
rect -11280 1913 -11246 1921
rect -11280 1887 -11246 1913
rect -11184 2831 -11150 2857
rect -11184 2823 -11150 2831
rect -11184 2763 -11150 2785
rect -11184 2751 -11150 2763
rect -11184 2695 -11150 2713
rect -11184 2679 -11150 2695
rect -11184 2627 -11150 2641
rect -11184 2607 -11150 2627
rect -11184 2559 -11150 2569
rect -11184 2535 -11150 2559
rect -11184 2491 -11150 2497
rect -11184 2463 -11150 2491
rect -11184 2423 -11150 2425
rect -11184 2391 -11150 2423
rect -11184 2321 -11150 2353
rect -11184 2319 -11150 2321
rect -11184 2253 -11150 2281
rect -11184 2247 -11150 2253
rect -11184 2185 -11150 2209
rect -11184 2175 -11150 2185
rect -11184 2117 -11150 2137
rect -11184 2103 -11150 2117
rect -11184 2049 -11150 2065
rect -11184 2031 -11150 2049
rect -11184 1981 -11150 1993
rect -11184 1959 -11150 1981
rect -11184 1913 -11150 1921
rect -11184 1887 -11150 1913
rect -10196 2823 -10162 2849
rect -10196 2815 -10162 2823
rect -10196 2755 -10162 2777
rect -10196 2743 -10162 2755
rect -10196 2687 -10162 2705
rect -10196 2671 -10162 2687
rect -10196 2619 -10162 2633
rect -10196 2599 -10162 2619
rect -10196 2551 -10162 2561
rect -10196 2527 -10162 2551
rect -10196 2483 -10162 2489
rect -10196 2455 -10162 2483
rect -10196 2415 -10162 2417
rect -10196 2383 -10162 2415
rect -10196 2313 -10162 2345
rect -10196 2311 -10162 2313
rect -10196 2245 -10162 2273
rect -10196 2239 -10162 2245
rect -10196 2177 -10162 2201
rect -10196 2167 -10162 2177
rect -10196 2109 -10162 2129
rect -10196 2095 -10162 2109
rect -10196 2041 -10162 2057
rect -10196 2023 -10162 2041
rect -10196 1973 -10162 1985
rect -10196 1951 -10162 1973
rect -10196 1905 -10162 1913
rect -10196 1879 -10162 1905
rect -10100 2823 -10066 2849
rect -10100 2815 -10066 2823
rect -10100 2755 -10066 2777
rect -10100 2743 -10066 2755
rect -10100 2687 -10066 2705
rect -10100 2671 -10066 2687
rect -10100 2619 -10066 2633
rect -10100 2599 -10066 2619
rect -10100 2551 -10066 2561
rect -10100 2527 -10066 2551
rect -10100 2483 -10066 2489
rect -10100 2455 -10066 2483
rect -10100 2415 -10066 2417
rect -10100 2383 -10066 2415
rect -10100 2313 -10066 2345
rect -10100 2311 -10066 2313
rect -10100 2245 -10066 2273
rect -10100 2239 -10066 2245
rect -10100 2177 -10066 2201
rect -10100 2167 -10066 2177
rect -10100 2109 -10066 2129
rect -10100 2095 -10066 2109
rect -10100 2041 -10066 2057
rect -10100 2023 -10066 2041
rect -10100 1973 -10066 1985
rect -10100 1951 -10066 1973
rect -10100 1905 -10066 1913
rect -10100 1879 -10066 1905
rect -10004 2823 -9970 2849
rect -10004 2815 -9970 2823
rect -10004 2755 -9970 2777
rect -10004 2743 -9970 2755
rect -10004 2687 -9970 2705
rect -10004 2671 -9970 2687
rect -10004 2619 -9970 2633
rect -10004 2599 -9970 2619
rect -10004 2551 -9970 2561
rect -10004 2527 -9970 2551
rect -10004 2483 -9970 2489
rect -10004 2455 -9970 2483
rect -10004 2415 -9970 2417
rect -10004 2383 -9970 2415
rect -10004 2313 -9970 2345
rect -10004 2311 -9970 2313
rect -10004 2245 -9970 2273
rect -10004 2239 -9970 2245
rect -10004 2177 -9970 2201
rect -10004 2167 -9970 2177
rect -10004 2109 -9970 2129
rect -10004 2095 -9970 2109
rect -10004 2041 -9970 2057
rect -10004 2023 -9970 2041
rect -10004 1973 -9970 1985
rect -10004 1951 -9970 1973
rect -10004 1905 -9970 1913
rect -10004 1879 -9970 1905
rect -9908 2823 -9874 2849
rect -9908 2815 -9874 2823
rect -9908 2755 -9874 2777
rect -9908 2743 -9874 2755
rect -9908 2687 -9874 2705
rect -9908 2671 -9874 2687
rect -9908 2619 -9874 2633
rect -9908 2599 -9874 2619
rect -9908 2551 -9874 2561
rect -9908 2527 -9874 2551
rect -9908 2483 -9874 2489
rect -9908 2455 -9874 2483
rect -9908 2415 -9874 2417
rect -9908 2383 -9874 2415
rect -9908 2313 -9874 2345
rect -9908 2311 -9874 2313
rect -9908 2245 -9874 2273
rect -9908 2239 -9874 2245
rect -9908 2177 -9874 2201
rect -9908 2167 -9874 2177
rect -9908 2109 -9874 2129
rect -9908 2095 -9874 2109
rect -9908 2041 -9874 2057
rect -9908 2023 -9874 2041
rect -9908 1973 -9874 1985
rect -9908 1951 -9874 1973
rect -9908 1905 -9874 1913
rect -9908 1879 -9874 1905
rect -9812 2823 -9778 2849
rect -9812 2815 -9778 2823
rect -9812 2755 -9778 2777
rect -9812 2743 -9778 2755
rect -9812 2687 -9778 2705
rect -9812 2671 -9778 2687
rect -9812 2619 -9778 2633
rect -9812 2599 -9778 2619
rect -9812 2551 -9778 2561
rect -9812 2527 -9778 2551
rect -9812 2483 -9778 2489
rect -9812 2455 -9778 2483
rect -9812 2415 -9778 2417
rect -9812 2383 -9778 2415
rect -9812 2313 -9778 2345
rect -9812 2311 -9778 2313
rect -9812 2245 -9778 2273
rect -9812 2239 -9778 2245
rect -9812 2177 -9778 2201
rect -9812 2167 -9778 2177
rect -9812 2109 -9778 2129
rect -9812 2095 -9778 2109
rect -9812 2041 -9778 2057
rect -9812 2023 -9778 2041
rect -9812 1973 -9778 1985
rect -9812 1951 -9778 1973
rect -9812 1905 -9778 1913
rect -9812 1879 -9778 1905
rect -9716 2823 -9682 2849
rect -9716 2815 -9682 2823
rect -9716 2755 -9682 2777
rect -9716 2743 -9682 2755
rect -9716 2687 -9682 2705
rect -9716 2671 -9682 2687
rect -9716 2619 -9682 2633
rect -9716 2599 -9682 2619
rect -9716 2551 -9682 2561
rect -9716 2527 -9682 2551
rect -9716 2483 -9682 2489
rect -9716 2455 -9682 2483
rect -9716 2415 -9682 2417
rect -9716 2383 -9682 2415
rect -9716 2313 -9682 2345
rect -9716 2311 -9682 2313
rect -9716 2245 -9682 2273
rect -9716 2239 -9682 2245
rect -9716 2177 -9682 2201
rect -9716 2167 -9682 2177
rect -9716 2109 -9682 2129
rect -9716 2095 -9682 2109
rect -9716 2041 -9682 2057
rect -9716 2023 -9682 2041
rect -9716 1973 -9682 1985
rect -9716 1951 -9682 1973
rect -9716 1905 -9682 1913
rect -9716 1879 -9682 1905
rect -9620 2823 -9586 2849
rect -9620 2815 -9586 2823
rect -9620 2755 -9586 2777
rect -9620 2743 -9586 2755
rect -9620 2687 -9586 2705
rect -9620 2671 -9586 2687
rect -9620 2619 -9586 2633
rect -9620 2599 -9586 2619
rect -9620 2551 -9586 2561
rect -9620 2527 -9586 2551
rect -9620 2483 -9586 2489
rect -9620 2455 -9586 2483
rect -9620 2415 -9586 2417
rect -9620 2383 -9586 2415
rect -9620 2313 -9586 2345
rect -9620 2311 -9586 2313
rect -9620 2245 -9586 2273
rect -9620 2239 -9586 2245
rect -9620 2177 -9586 2201
rect -9620 2167 -9586 2177
rect -9620 2109 -9586 2129
rect -9620 2095 -9586 2109
rect -9620 2041 -9586 2057
rect -9620 2023 -9586 2041
rect -9620 1973 -9586 1985
rect -9620 1951 -9586 1973
rect -9620 1905 -9586 1913
rect -9620 1879 -9586 1905
rect -9524 2823 -9490 2849
rect -9524 2815 -9490 2823
rect -9524 2755 -9490 2777
rect -9524 2743 -9490 2755
rect -9524 2687 -9490 2705
rect -9524 2671 -9490 2687
rect -9524 2619 -9490 2633
rect -9524 2599 -9490 2619
rect -9524 2551 -9490 2561
rect -9524 2527 -9490 2551
rect -9524 2483 -9490 2489
rect -9524 2455 -9490 2483
rect -9524 2415 -9490 2417
rect -9524 2383 -9490 2415
rect -9524 2313 -9490 2345
rect -9524 2311 -9490 2313
rect -9524 2245 -9490 2273
rect -9524 2239 -9490 2245
rect -9524 2177 -9490 2201
rect -9524 2167 -9490 2177
rect -9524 2109 -9490 2129
rect -9524 2095 -9490 2109
rect -9524 2041 -9490 2057
rect -9524 2023 -9490 2041
rect -9524 1973 -9490 1985
rect -9524 1951 -9490 1973
rect -9524 1905 -9490 1913
rect -9524 1879 -9490 1905
rect -9428 2823 -9394 2849
rect -9428 2815 -9394 2823
rect -9428 2755 -9394 2777
rect -9428 2743 -9394 2755
rect -9428 2687 -9394 2705
rect -9428 2671 -9394 2687
rect -9428 2619 -9394 2633
rect -9428 2599 -9394 2619
rect -9428 2551 -9394 2561
rect -9428 2527 -9394 2551
rect -9428 2483 -9394 2489
rect -9428 2455 -9394 2483
rect -9428 2415 -9394 2417
rect -9428 2383 -9394 2415
rect -9428 2313 -9394 2345
rect -9428 2311 -9394 2313
rect -9428 2245 -9394 2273
rect -9428 2239 -9394 2245
rect -9428 2177 -9394 2201
rect -9428 2167 -9394 2177
rect -9428 2109 -9394 2129
rect -9428 2095 -9394 2109
rect -9428 2041 -9394 2057
rect -9428 2023 -9394 2041
rect -9428 1973 -9394 1985
rect -9428 1951 -9394 1973
rect -9428 1905 -9394 1913
rect -9428 1879 -9394 1905
rect -9332 2823 -9298 2849
rect -9332 2815 -9298 2823
rect -9332 2755 -9298 2777
rect -9332 2743 -9298 2755
rect -9332 2687 -9298 2705
rect -9332 2671 -9298 2687
rect -9332 2619 -9298 2633
rect -9332 2599 -9298 2619
rect -9332 2551 -9298 2561
rect -9332 2527 -9298 2551
rect -9332 2483 -9298 2489
rect -9332 2455 -9298 2483
rect -9332 2415 -9298 2417
rect -9332 2383 -9298 2415
rect -9332 2313 -9298 2345
rect -9332 2311 -9298 2313
rect -9332 2245 -9298 2273
rect -9332 2239 -9298 2245
rect -9332 2177 -9298 2201
rect -9332 2167 -9298 2177
rect -9332 2109 -9298 2129
rect -9332 2095 -9298 2109
rect -9332 2041 -9298 2057
rect -9332 2023 -9298 2041
rect -9332 1973 -9298 1985
rect -9332 1951 -9298 1973
rect -9332 1905 -9298 1913
rect -9332 1879 -9298 1905
rect -9236 2823 -9202 2849
rect -9236 2815 -9202 2823
rect -9236 2755 -9202 2777
rect -9236 2743 -9202 2755
rect -9236 2687 -9202 2705
rect -9236 2671 -9202 2687
rect -9236 2619 -9202 2633
rect -9236 2599 -9202 2619
rect -9236 2551 -9202 2561
rect -9236 2527 -9202 2551
rect -9236 2483 -9202 2489
rect -9236 2455 -9202 2483
rect -9236 2415 -9202 2417
rect -9236 2383 -9202 2415
rect -9236 2313 -9202 2345
rect -9236 2311 -9202 2313
rect -9236 2245 -9202 2273
rect -9236 2239 -9202 2245
rect -9236 2177 -9202 2201
rect -9236 2167 -9202 2177
rect -9236 2109 -9202 2129
rect -9236 2095 -9202 2109
rect -9236 2041 -9202 2057
rect -9236 2023 -9202 2041
rect -9236 1973 -9202 1985
rect -9236 1951 -9202 1973
rect -9236 1905 -9202 1913
rect -9236 1879 -9202 1905
rect -9140 2823 -9106 2849
rect -9140 2815 -9106 2823
rect -9140 2755 -9106 2777
rect -9140 2743 -9106 2755
rect -9140 2687 -9106 2705
rect -9140 2671 -9106 2687
rect -9140 2619 -9106 2633
rect -9140 2599 -9106 2619
rect -9140 2551 -9106 2561
rect -9140 2527 -9106 2551
rect -9140 2483 -9106 2489
rect -9140 2455 -9106 2483
rect -9140 2415 -9106 2417
rect -9140 2383 -9106 2415
rect -9140 2313 -9106 2345
rect -9140 2311 -9106 2313
rect -9140 2245 -9106 2273
rect -9140 2239 -9106 2245
rect -9140 2177 -9106 2201
rect -9140 2167 -9106 2177
rect -9140 2109 -9106 2129
rect -9140 2095 -9106 2109
rect -9140 2041 -9106 2057
rect -9140 2023 -9106 2041
rect -9140 1973 -9106 1985
rect -9140 1951 -9106 1973
rect -9140 1905 -9106 1913
rect -9140 1879 -9106 1905
rect -9044 2823 -9010 2849
rect -9044 2815 -9010 2823
rect -9044 2755 -9010 2777
rect -9044 2743 -9010 2755
rect -9044 2687 -9010 2705
rect -9044 2671 -9010 2687
rect -9044 2619 -9010 2633
rect -9044 2599 -9010 2619
rect -9044 2551 -9010 2561
rect -9044 2527 -9010 2551
rect -9044 2483 -9010 2489
rect -9044 2455 -9010 2483
rect -9044 2415 -9010 2417
rect -9044 2383 -9010 2415
rect -9044 2313 -9010 2345
rect -9044 2311 -9010 2313
rect -9044 2245 -9010 2273
rect -9044 2239 -9010 2245
rect -9044 2177 -9010 2201
rect -9044 2167 -9010 2177
rect -9044 2109 -9010 2129
rect -9044 2095 -9010 2109
rect -9044 2041 -9010 2057
rect -9044 2023 -9010 2041
rect -9044 1973 -9010 1985
rect -9044 1951 -9010 1973
rect -9044 1905 -9010 1913
rect -9044 1879 -9010 1905
rect -8948 2823 -8914 2849
rect -8948 2815 -8914 2823
rect -8948 2755 -8914 2777
rect -8948 2743 -8914 2755
rect -8948 2687 -8914 2705
rect -8948 2671 -8914 2687
rect -8948 2619 -8914 2633
rect -8948 2599 -8914 2619
rect -8948 2551 -8914 2561
rect -8948 2527 -8914 2551
rect -8948 2483 -8914 2489
rect -8948 2455 -8914 2483
rect -8948 2415 -8914 2417
rect -8948 2383 -8914 2415
rect -8948 2313 -8914 2345
rect -8948 2311 -8914 2313
rect -8948 2245 -8914 2273
rect -8948 2239 -8914 2245
rect -8948 2177 -8914 2201
rect -8948 2167 -8914 2177
rect -8948 2109 -8914 2129
rect -8948 2095 -8914 2109
rect -8948 2041 -8914 2057
rect -8948 2023 -8914 2041
rect -8948 1973 -8914 1985
rect -8948 1951 -8914 1973
rect -8948 1905 -8914 1913
rect -8948 1879 -8914 1905
rect -8852 2823 -8818 2849
rect -8852 2815 -8818 2823
rect -8852 2755 -8818 2777
rect -8852 2743 -8818 2755
rect -8852 2687 -8818 2705
rect -8852 2671 -8818 2687
rect -8852 2619 -8818 2633
rect -8852 2599 -8818 2619
rect -8852 2551 -8818 2561
rect -8852 2527 -8818 2551
rect -8852 2483 -8818 2489
rect -8852 2455 -8818 2483
rect -8852 2415 -8818 2417
rect -8852 2383 -8818 2415
rect -8852 2313 -8818 2345
rect -8852 2311 -8818 2313
rect -8852 2245 -8818 2273
rect -8852 2239 -8818 2245
rect -8852 2177 -8818 2201
rect -8852 2167 -8818 2177
rect -8852 2109 -8818 2129
rect -8852 2095 -8818 2109
rect -8852 2041 -8818 2057
rect -8852 2023 -8818 2041
rect -8852 1973 -8818 1985
rect -8852 1951 -8818 1973
rect -8852 1905 -8818 1913
rect -8852 1879 -8818 1905
rect -8756 2823 -8722 2849
rect -8756 2815 -8722 2823
rect -8756 2755 -8722 2777
rect -8756 2743 -8722 2755
rect -8756 2687 -8722 2705
rect -8756 2671 -8722 2687
rect -8756 2619 -8722 2633
rect -8756 2599 -8722 2619
rect -8756 2551 -8722 2561
rect -8756 2527 -8722 2551
rect -8756 2483 -8722 2489
rect -8756 2455 -8722 2483
rect -8756 2415 -8722 2417
rect -8756 2383 -8722 2415
rect -8756 2313 -8722 2345
rect -8756 2311 -8722 2313
rect -8756 2245 -8722 2273
rect -8756 2239 -8722 2245
rect -8756 2177 -8722 2201
rect -8756 2167 -8722 2177
rect -8756 2109 -8722 2129
rect -8756 2095 -8722 2109
rect -8756 2041 -8722 2057
rect -8756 2023 -8722 2041
rect -8756 1973 -8722 1985
rect -8756 1951 -8722 1973
rect -8756 1905 -8722 1913
rect -8756 1879 -8722 1905
rect -8660 2823 -8626 2849
rect -8660 2815 -8626 2823
rect -8660 2755 -8626 2777
rect -8660 2743 -8626 2755
rect -8660 2687 -8626 2705
rect -8660 2671 -8626 2687
rect -8660 2619 -8626 2633
rect -8660 2599 -8626 2619
rect -8660 2551 -8626 2561
rect -8660 2527 -8626 2551
rect -8660 2483 -8626 2489
rect -8660 2455 -8626 2483
rect -8660 2415 -8626 2417
rect -8660 2383 -8626 2415
rect -8660 2313 -8626 2345
rect -8660 2311 -8626 2313
rect -8660 2245 -8626 2273
rect -8660 2239 -8626 2245
rect -8660 2177 -8626 2201
rect -8660 2167 -8626 2177
rect -8660 2109 -8626 2129
rect -8660 2095 -8626 2109
rect -8660 2041 -8626 2057
rect -8660 2023 -8626 2041
rect -8660 1973 -8626 1985
rect -8660 1951 -8626 1973
rect -8660 1905 -8626 1913
rect -8660 1879 -8626 1905
rect -8564 2823 -8530 2849
rect -8564 2815 -8530 2823
rect -8564 2755 -8530 2777
rect -8564 2743 -8530 2755
rect -8564 2687 -8530 2705
rect -8564 2671 -8530 2687
rect -8564 2619 -8530 2633
rect -8564 2599 -8530 2619
rect -8564 2551 -8530 2561
rect -8564 2527 -8530 2551
rect -8564 2483 -8530 2489
rect -8564 2455 -8530 2483
rect -8564 2415 -8530 2417
rect -8564 2383 -8530 2415
rect -8564 2313 -8530 2345
rect -8564 2311 -8530 2313
rect -8564 2245 -8530 2273
rect -8564 2239 -8530 2245
rect -8564 2177 -8530 2201
rect -8564 2167 -8530 2177
rect -8564 2109 -8530 2129
rect -8564 2095 -8530 2109
rect -8564 2041 -8530 2057
rect -8564 2023 -8530 2041
rect -8564 1973 -8530 1985
rect -8564 1951 -8530 1973
rect -8564 1905 -8530 1913
rect -8564 1879 -8530 1905
rect -8468 2823 -8434 2849
rect -8468 2815 -8434 2823
rect -8468 2755 -8434 2777
rect -8468 2743 -8434 2755
rect -8468 2687 -8434 2705
rect -8468 2671 -8434 2687
rect -8468 2619 -8434 2633
rect -8468 2599 -8434 2619
rect -8468 2551 -8434 2561
rect -8468 2527 -8434 2551
rect -8468 2483 -8434 2489
rect -8468 2455 -8434 2483
rect -8468 2415 -8434 2417
rect -8468 2383 -8434 2415
rect -8468 2313 -8434 2345
rect -8468 2311 -8434 2313
rect -8468 2245 -8434 2273
rect -8468 2239 -8434 2245
rect -8468 2177 -8434 2201
rect -8468 2167 -8434 2177
rect -8468 2109 -8434 2129
rect -8468 2095 -8434 2109
rect -8468 2041 -8434 2057
rect -8468 2023 -8434 2041
rect -8468 1973 -8434 1985
rect -8468 1951 -8434 1973
rect -8468 1905 -8434 1913
rect -8468 1879 -8434 1905
rect -8372 2823 -8338 2849
rect -8372 2815 -8338 2823
rect -8372 2755 -8338 2777
rect -8372 2743 -8338 2755
rect -8372 2687 -8338 2705
rect -8372 2671 -8338 2687
rect -8372 2619 -8338 2633
rect -8372 2599 -8338 2619
rect -8372 2551 -8338 2561
rect -8372 2527 -8338 2551
rect -8372 2483 -8338 2489
rect -8372 2455 -8338 2483
rect -8372 2415 -8338 2417
rect -8372 2383 -8338 2415
rect -8372 2313 -8338 2345
rect -8372 2311 -8338 2313
rect -8372 2245 -8338 2273
rect -8372 2239 -8338 2245
rect -8372 2177 -8338 2201
rect -8372 2167 -8338 2177
rect -8372 2109 -8338 2129
rect -8372 2095 -8338 2109
rect -8372 2041 -8338 2057
rect -8372 2023 -8338 2041
rect -8372 1973 -8338 1985
rect -8372 1951 -8338 1973
rect -8372 1905 -8338 1913
rect -8372 1879 -8338 1905
rect -8276 2823 -8242 2849
rect -8276 2815 -8242 2823
rect -8276 2755 -8242 2777
rect -8276 2743 -8242 2755
rect -8276 2687 -8242 2705
rect -8276 2671 -8242 2687
rect -8276 2619 -8242 2633
rect -8276 2599 -8242 2619
rect -8276 2551 -8242 2561
rect -8276 2527 -8242 2551
rect -8276 2483 -8242 2489
rect -8276 2455 -8242 2483
rect -8276 2415 -8242 2417
rect -8276 2383 -8242 2415
rect -8276 2313 -8242 2345
rect -8276 2311 -8242 2313
rect -8276 2245 -8242 2273
rect -8276 2239 -8242 2245
rect -8276 2177 -8242 2201
rect -8276 2167 -8242 2177
rect -8276 2109 -8242 2129
rect -8276 2095 -8242 2109
rect -8276 2041 -8242 2057
rect -8276 2023 -8242 2041
rect -8276 1973 -8242 1985
rect -8276 1951 -8242 1973
rect -8276 1905 -8242 1913
rect -8276 1879 -8242 1905
rect -8048 2815 -8014 2841
rect -8048 2807 -8014 2815
rect -8048 2747 -8014 2769
rect -8048 2735 -8014 2747
rect -8048 2679 -8014 2697
rect -8048 2663 -8014 2679
rect -8048 2611 -8014 2625
rect -8048 2591 -8014 2611
rect -8048 2543 -8014 2553
rect -8048 2519 -8014 2543
rect -8048 2475 -8014 2481
rect -8048 2447 -8014 2475
rect -8048 2407 -8014 2409
rect -8048 2375 -8014 2407
rect -8048 2305 -8014 2337
rect -8048 2303 -8014 2305
rect -8048 2237 -8014 2265
rect -8048 2231 -8014 2237
rect -8048 2169 -8014 2193
rect -8048 2159 -8014 2169
rect -8048 2101 -8014 2121
rect -8048 2087 -8014 2101
rect -8048 2033 -8014 2049
rect -8048 2015 -8014 2033
rect -8048 1965 -8014 1977
rect -8048 1943 -8014 1965
rect -8048 1897 -8014 1905
rect -8048 1871 -8014 1897
rect -7952 2815 -7918 2841
rect -7952 2807 -7918 2815
rect -7952 2747 -7918 2769
rect -7952 2735 -7918 2747
rect -7952 2679 -7918 2697
rect -7952 2663 -7918 2679
rect -7952 2611 -7918 2625
rect -7952 2591 -7918 2611
rect -7952 2543 -7918 2553
rect -7952 2519 -7918 2543
rect -7952 2475 -7918 2481
rect -7952 2447 -7918 2475
rect -7952 2407 -7918 2409
rect -7952 2375 -7918 2407
rect -7952 2305 -7918 2337
rect -7952 2303 -7918 2305
rect -7952 2237 -7918 2265
rect -7952 2231 -7918 2237
rect -7952 2169 -7918 2193
rect -7952 2159 -7918 2169
rect -7952 2101 -7918 2121
rect -7952 2087 -7918 2101
rect -7952 2033 -7918 2049
rect -7952 2015 -7918 2033
rect -7952 1965 -7918 1977
rect -7952 1943 -7918 1965
rect -7952 1897 -7918 1905
rect -7952 1871 -7918 1897
rect -7856 2815 -7822 2841
rect -7856 2807 -7822 2815
rect -7856 2747 -7822 2769
rect -7856 2735 -7822 2747
rect -7856 2679 -7822 2697
rect -7856 2663 -7822 2679
rect -7856 2611 -7822 2625
rect -7856 2591 -7822 2611
rect -7856 2543 -7822 2553
rect -7856 2519 -7822 2543
rect -7856 2475 -7822 2481
rect -7856 2447 -7822 2475
rect -7856 2407 -7822 2409
rect -7856 2375 -7822 2407
rect -7856 2305 -7822 2337
rect -7856 2303 -7822 2305
rect -7856 2237 -7822 2265
rect -7856 2231 -7822 2237
rect -7856 2169 -7822 2193
rect -7856 2159 -7822 2169
rect -7856 2101 -7822 2121
rect -7856 2087 -7822 2101
rect -7856 2033 -7822 2049
rect -7856 2015 -7822 2033
rect -7856 1965 -7822 1977
rect -7856 1943 -7822 1965
rect -7856 1897 -7822 1905
rect -7856 1871 -7822 1897
rect -7760 2815 -7726 2841
rect -7760 2807 -7726 2815
rect -7760 2747 -7726 2769
rect -7760 2735 -7726 2747
rect -7760 2679 -7726 2697
rect -7760 2663 -7726 2679
rect -7760 2611 -7726 2625
rect -7760 2591 -7726 2611
rect -7760 2543 -7726 2553
rect -7760 2519 -7726 2543
rect -7760 2475 -7726 2481
rect -7760 2447 -7726 2475
rect -7760 2407 -7726 2409
rect -7760 2375 -7726 2407
rect -7760 2305 -7726 2337
rect -7760 2303 -7726 2305
rect -7760 2237 -7726 2265
rect -7760 2231 -7726 2237
rect -7760 2169 -7726 2193
rect -7760 2159 -7726 2169
rect -7760 2101 -7726 2121
rect -7760 2087 -7726 2101
rect -7760 2033 -7726 2049
rect -7760 2015 -7726 2033
rect -7760 1965 -7726 1977
rect -7760 1943 -7726 1965
rect -7760 1897 -7726 1905
rect -7760 1871 -7726 1897
rect -7664 2815 -7630 2841
rect -7664 2807 -7630 2815
rect -7664 2747 -7630 2769
rect -7664 2735 -7630 2747
rect -7664 2679 -7630 2697
rect -7664 2663 -7630 2679
rect -7664 2611 -7630 2625
rect -7664 2591 -7630 2611
rect -7664 2543 -7630 2553
rect -7664 2519 -7630 2543
rect -7664 2475 -7630 2481
rect -7664 2447 -7630 2475
rect -7664 2407 -7630 2409
rect -7664 2375 -7630 2407
rect -7664 2305 -7630 2337
rect -7664 2303 -7630 2305
rect -7664 2237 -7630 2265
rect -7664 2231 -7630 2237
rect -7664 2169 -7630 2193
rect -7664 2159 -7630 2169
rect -7664 2101 -7630 2121
rect -7664 2087 -7630 2101
rect -7664 2033 -7630 2049
rect -7664 2015 -7630 2033
rect -7664 1965 -7630 1977
rect -7664 1943 -7630 1965
rect -7664 1897 -7630 1905
rect -7664 1871 -7630 1897
rect -7568 2815 -7534 2841
rect -7568 2807 -7534 2815
rect -7568 2747 -7534 2769
rect -7568 2735 -7534 2747
rect -7568 2679 -7534 2697
rect -7568 2663 -7534 2679
rect -7568 2611 -7534 2625
rect -7568 2591 -7534 2611
rect -7568 2543 -7534 2553
rect -7568 2519 -7534 2543
rect -7568 2475 -7534 2481
rect -7568 2447 -7534 2475
rect -7568 2407 -7534 2409
rect -7568 2375 -7534 2407
rect -7568 2305 -7534 2337
rect -7568 2303 -7534 2305
rect -7568 2237 -7534 2265
rect -7568 2231 -7534 2237
rect -7568 2169 -7534 2193
rect -7568 2159 -7534 2169
rect -7568 2101 -7534 2121
rect -7568 2087 -7534 2101
rect -7568 2033 -7534 2049
rect -7568 2015 -7534 2033
rect -7568 1965 -7534 1977
rect -7568 1943 -7534 1965
rect -7568 1897 -7534 1905
rect -7568 1871 -7534 1897
rect -7472 2815 -7438 2841
rect -7472 2807 -7438 2815
rect -7472 2747 -7438 2769
rect -7472 2735 -7438 2747
rect -7472 2679 -7438 2697
rect -7472 2663 -7438 2679
rect -7472 2611 -7438 2625
rect -7472 2591 -7438 2611
rect -7472 2543 -7438 2553
rect -7472 2519 -7438 2543
rect -7472 2475 -7438 2481
rect -7472 2447 -7438 2475
rect -7472 2407 -7438 2409
rect -7472 2375 -7438 2407
rect -7472 2305 -7438 2337
rect -7472 2303 -7438 2305
rect -7472 2237 -7438 2265
rect -7472 2231 -7438 2237
rect -7472 2169 -7438 2193
rect -7472 2159 -7438 2169
rect -7472 2101 -7438 2121
rect -7472 2087 -7438 2101
rect -7472 2033 -7438 2049
rect -7472 2015 -7438 2033
rect -7472 1965 -7438 1977
rect -7472 1943 -7438 1965
rect -7472 1897 -7438 1905
rect -7472 1871 -7438 1897
rect -7376 2815 -7342 2841
rect -7376 2807 -7342 2815
rect -7376 2747 -7342 2769
rect -7376 2735 -7342 2747
rect -7376 2679 -7342 2697
rect -7376 2663 -7342 2679
rect -7376 2611 -7342 2625
rect -7376 2591 -7342 2611
rect -7376 2543 -7342 2553
rect -7376 2519 -7342 2543
rect -7376 2475 -7342 2481
rect -7376 2447 -7342 2475
rect -7376 2407 -7342 2409
rect -7376 2375 -7342 2407
rect -7376 2305 -7342 2337
rect -7376 2303 -7342 2305
rect -7376 2237 -7342 2265
rect -7376 2231 -7342 2237
rect -7376 2169 -7342 2193
rect -7376 2159 -7342 2169
rect -7376 2101 -7342 2121
rect -7376 2087 -7342 2101
rect -7376 2033 -7342 2049
rect -7376 2015 -7342 2033
rect -7376 1965 -7342 1977
rect -7376 1943 -7342 1965
rect -7376 1897 -7342 1905
rect -7376 1871 -7342 1897
rect -7280 2815 -7246 2841
rect -7280 2807 -7246 2815
rect -7280 2747 -7246 2769
rect -7280 2735 -7246 2747
rect -7280 2679 -7246 2697
rect -7280 2663 -7246 2679
rect -7280 2611 -7246 2625
rect -7280 2591 -7246 2611
rect -7280 2543 -7246 2553
rect -7280 2519 -7246 2543
rect -7280 2475 -7246 2481
rect -7280 2447 -7246 2475
rect -7280 2407 -7246 2409
rect -7280 2375 -7246 2407
rect -7280 2305 -7246 2337
rect -7280 2303 -7246 2305
rect -7280 2237 -7246 2265
rect -7280 2231 -7246 2237
rect -7280 2169 -7246 2193
rect -7280 2159 -7246 2169
rect -7280 2101 -7246 2121
rect -7280 2087 -7246 2101
rect -7280 2033 -7246 2049
rect -7280 2015 -7246 2033
rect -7280 1965 -7246 1977
rect -7280 1943 -7246 1965
rect -7280 1897 -7246 1905
rect -7280 1871 -7246 1897
rect -7184 2815 -7150 2841
rect -7184 2807 -7150 2815
rect -7184 2747 -7150 2769
rect -7184 2735 -7150 2747
rect -7184 2679 -7150 2697
rect -7184 2663 -7150 2679
rect -7184 2611 -7150 2625
rect -7184 2591 -7150 2611
rect -7184 2543 -7150 2553
rect -7184 2519 -7150 2543
rect -7184 2475 -7150 2481
rect -7184 2447 -7150 2475
rect -7184 2407 -7150 2409
rect -7184 2375 -7150 2407
rect -7184 2305 -7150 2337
rect -7184 2303 -7150 2305
rect -7184 2237 -7150 2265
rect -7184 2231 -7150 2237
rect -7184 2169 -7150 2193
rect -7184 2159 -7150 2169
rect -7184 2101 -7150 2121
rect -7184 2087 -7150 2101
rect -7184 2033 -7150 2049
rect -7184 2015 -7150 2033
rect -7184 1965 -7150 1977
rect -7184 1943 -7150 1965
rect -7184 1897 -7150 1905
rect -7184 1871 -7150 1897
rect -7088 2815 -7054 2841
rect -7088 2807 -7054 2815
rect -7088 2747 -7054 2769
rect -7088 2735 -7054 2747
rect -7088 2679 -7054 2697
rect -7088 2663 -7054 2679
rect -7088 2611 -7054 2625
rect -7088 2591 -7054 2611
rect -7088 2543 -7054 2553
rect -7088 2519 -7054 2543
rect -7088 2475 -7054 2481
rect -7088 2447 -7054 2475
rect -7088 2407 -7054 2409
rect -7088 2375 -7054 2407
rect -7088 2305 -7054 2337
rect -7088 2303 -7054 2305
rect -7088 2237 -7054 2265
rect -7088 2231 -7054 2237
rect -7088 2169 -7054 2193
rect -7088 2159 -7054 2169
rect -7088 2101 -7054 2121
rect -7088 2087 -7054 2101
rect -7088 2033 -7054 2049
rect -7088 2015 -7054 2033
rect -7088 1965 -7054 1977
rect -7088 1943 -7054 1965
rect -7088 1897 -7054 1905
rect -7088 1871 -7054 1897
rect -6992 2815 -6958 2841
rect -6992 2807 -6958 2815
rect -6992 2747 -6958 2769
rect -6992 2735 -6958 2747
rect -6992 2679 -6958 2697
rect -6992 2663 -6958 2679
rect -6992 2611 -6958 2625
rect -6992 2591 -6958 2611
rect -6992 2543 -6958 2553
rect -6992 2519 -6958 2543
rect -6992 2475 -6958 2481
rect -6992 2447 -6958 2475
rect -6992 2407 -6958 2409
rect -6992 2375 -6958 2407
rect -6992 2305 -6958 2337
rect -6992 2303 -6958 2305
rect -6992 2237 -6958 2265
rect -6992 2231 -6958 2237
rect -6992 2169 -6958 2193
rect -6992 2159 -6958 2169
rect -6992 2101 -6958 2121
rect -6992 2087 -6958 2101
rect -6992 2033 -6958 2049
rect -6992 2015 -6958 2033
rect -6992 1965 -6958 1977
rect -6992 1943 -6958 1965
rect -6992 1897 -6958 1905
rect -6992 1871 -6958 1897
rect -6896 2815 -6862 2841
rect -6896 2807 -6862 2815
rect -6896 2747 -6862 2769
rect -6896 2735 -6862 2747
rect -6896 2679 -6862 2697
rect -6896 2663 -6862 2679
rect -6896 2611 -6862 2625
rect -6896 2591 -6862 2611
rect -6896 2543 -6862 2553
rect -6896 2519 -6862 2543
rect -6896 2475 -6862 2481
rect -6896 2447 -6862 2475
rect -6896 2407 -6862 2409
rect -6896 2375 -6862 2407
rect -6896 2305 -6862 2337
rect -6896 2303 -6862 2305
rect -6896 2237 -6862 2265
rect -6896 2231 -6862 2237
rect -6896 2169 -6862 2193
rect -6896 2159 -6862 2169
rect -6896 2101 -6862 2121
rect -6896 2087 -6862 2101
rect -6896 2033 -6862 2049
rect -6896 2015 -6862 2033
rect -6896 1965 -6862 1977
rect -6896 1943 -6862 1965
rect -6896 1897 -6862 1905
rect -6896 1871 -6862 1897
rect -6800 2815 -6766 2841
rect -6800 2807 -6766 2815
rect -6800 2747 -6766 2769
rect -6800 2735 -6766 2747
rect -6800 2679 -6766 2697
rect -6800 2663 -6766 2679
rect -6800 2611 -6766 2625
rect -6800 2591 -6766 2611
rect -6800 2543 -6766 2553
rect -6800 2519 -6766 2543
rect -6800 2475 -6766 2481
rect -6800 2447 -6766 2475
rect -6800 2407 -6766 2409
rect -6800 2375 -6766 2407
rect -6800 2305 -6766 2337
rect -6800 2303 -6766 2305
rect -6800 2237 -6766 2265
rect -6800 2231 -6766 2237
rect -6800 2169 -6766 2193
rect -6800 2159 -6766 2169
rect -6800 2101 -6766 2121
rect -6800 2087 -6766 2101
rect -6800 2033 -6766 2049
rect -6800 2015 -6766 2033
rect -6800 1965 -6766 1977
rect -6800 1943 -6766 1965
rect -6800 1897 -6766 1905
rect -6800 1871 -6766 1897
rect -1686 3195 -1652 3221
rect -1686 3187 -1652 3195
rect -1686 3127 -1652 3149
rect -1686 3115 -1652 3127
rect -1686 3059 -1652 3077
rect -1686 3043 -1652 3059
rect -4862 3008 -4828 3042
rect -1686 2991 -1652 3005
rect -1686 2971 -1652 2991
rect -6704 2815 -6670 2841
rect -6704 2807 -6670 2815
rect -6704 2747 -6670 2769
rect -6704 2735 -6670 2747
rect -6704 2679 -6670 2697
rect -6704 2663 -6670 2679
rect -6704 2611 -6670 2625
rect -6704 2591 -6670 2611
rect -6704 2543 -6670 2553
rect -6704 2519 -6670 2543
rect -6704 2475 -6670 2481
rect -6704 2447 -6670 2475
rect -6704 2407 -6670 2409
rect -6704 2375 -6670 2407
rect -6704 2305 -6670 2337
rect -6704 2303 -6670 2305
rect -6704 2237 -6670 2265
rect -6704 2231 -6670 2237
rect -6704 2169 -6670 2193
rect -6704 2159 -6670 2169
rect -6704 2101 -6670 2121
rect -6704 2087 -6670 2101
rect -6704 2033 -6670 2049
rect -6704 2015 -6670 2033
rect -6704 1965 -6670 1977
rect -6704 1943 -6670 1965
rect -6704 1897 -6670 1905
rect -6704 1871 -6670 1897
rect -6608 2815 -6574 2841
rect -6608 2807 -6574 2815
rect -6608 2747 -6574 2769
rect -6608 2735 -6574 2747
rect -6608 2679 -6574 2697
rect -6608 2663 -6574 2679
rect -6608 2611 -6574 2625
rect -6608 2591 -6574 2611
rect -6608 2543 -6574 2553
rect -6608 2519 -6574 2543
rect -6608 2475 -6574 2481
rect -6608 2447 -6574 2475
rect -6608 2407 -6574 2409
rect -6608 2375 -6574 2407
rect -6608 2305 -6574 2337
rect -6608 2303 -6574 2305
rect -6608 2237 -6574 2265
rect -6608 2231 -6574 2237
rect -6608 2169 -6574 2193
rect -6608 2159 -6574 2169
rect -6608 2101 -6574 2121
rect -6608 2087 -6574 2101
rect -6608 2033 -6574 2049
rect -6608 2015 -6574 2033
rect -6608 1965 -6574 1977
rect -6608 1943 -6574 1965
rect -6608 1897 -6574 1905
rect -6608 1871 -6574 1897
rect -6370 2819 -6336 2845
rect -6370 2811 -6336 2819
rect -6370 2751 -6336 2773
rect -6370 2739 -6336 2751
rect -6370 2683 -6336 2701
rect -6370 2667 -6336 2683
rect -6370 2615 -6336 2629
rect -6370 2595 -6336 2615
rect -6370 2547 -6336 2557
rect -6370 2523 -6336 2547
rect -6370 2479 -6336 2485
rect -6370 2451 -6336 2479
rect -6370 2411 -6336 2413
rect -6370 2379 -6336 2411
rect -6370 2309 -6336 2341
rect -6370 2307 -6336 2309
rect -6370 2241 -6336 2269
rect -6370 2235 -6336 2241
rect -6370 2173 -6336 2197
rect -6370 2163 -6336 2173
rect -6370 2105 -6336 2125
rect -6370 2091 -6336 2105
rect -6370 2037 -6336 2053
rect -6370 2019 -6336 2037
rect -6370 1969 -6336 1981
rect -6370 1947 -6336 1969
rect -6370 1901 -6336 1909
rect -6370 1875 -6336 1901
rect -6274 2819 -6240 2845
rect -6274 2811 -6240 2819
rect -6274 2751 -6240 2773
rect -6274 2739 -6240 2751
rect -6274 2683 -6240 2701
rect -6274 2667 -6240 2683
rect -6274 2615 -6240 2629
rect -6274 2595 -6240 2615
rect -6274 2547 -6240 2557
rect -6274 2523 -6240 2547
rect -6274 2479 -6240 2485
rect -6274 2451 -6240 2479
rect -6274 2411 -6240 2413
rect -6274 2379 -6240 2411
rect -6274 2309 -6240 2341
rect -6274 2307 -6240 2309
rect -6274 2241 -6240 2269
rect -6274 2235 -6240 2241
rect -6274 2173 -6240 2197
rect -6274 2163 -6240 2173
rect -6274 2105 -6240 2125
rect -6274 2091 -6240 2105
rect -6274 2037 -6240 2053
rect -6274 2019 -6240 2037
rect -6274 1969 -6240 1981
rect -6274 1947 -6240 1969
rect -6274 1901 -6240 1909
rect -6274 1875 -6240 1901
rect -6178 2819 -6144 2845
rect -6178 2811 -6144 2819
rect -6178 2751 -6144 2773
rect -6178 2739 -6144 2751
rect -6178 2683 -6144 2701
rect -6178 2667 -6144 2683
rect -6178 2615 -6144 2629
rect -6178 2595 -6144 2615
rect -6178 2547 -6144 2557
rect -6178 2523 -6144 2547
rect -6178 2479 -6144 2485
rect -6178 2451 -6144 2479
rect -6178 2411 -6144 2413
rect -6178 2379 -6144 2411
rect -6178 2309 -6144 2341
rect -6178 2307 -6144 2309
rect -6178 2241 -6144 2269
rect -6178 2235 -6144 2241
rect -6178 2173 -6144 2197
rect -6178 2163 -6144 2173
rect -6178 2105 -6144 2125
rect -6178 2091 -6144 2105
rect -6178 2037 -6144 2053
rect -6178 2019 -6144 2037
rect -6178 1969 -6144 1981
rect -6178 1947 -6144 1969
rect -6178 1901 -6144 1909
rect -6178 1875 -6144 1901
rect -6082 2819 -6048 2845
rect -6082 2811 -6048 2819
rect -6082 2751 -6048 2773
rect -6082 2739 -6048 2751
rect -6082 2683 -6048 2701
rect -6082 2667 -6048 2683
rect -6082 2615 -6048 2629
rect -6082 2595 -6048 2615
rect -6082 2547 -6048 2557
rect -6082 2523 -6048 2547
rect -6082 2479 -6048 2485
rect -6082 2451 -6048 2479
rect -6082 2411 -6048 2413
rect -6082 2379 -6048 2411
rect -6082 2309 -6048 2341
rect -6082 2307 -6048 2309
rect -6082 2241 -6048 2269
rect -6082 2235 -6048 2241
rect -6082 2173 -6048 2197
rect -6082 2163 -6048 2173
rect -6082 2105 -6048 2125
rect -6082 2091 -6048 2105
rect -6082 2037 -6048 2053
rect -6082 2019 -6048 2037
rect -6082 1969 -6048 1981
rect -6082 1947 -6048 1969
rect -6082 1901 -6048 1909
rect -6082 1875 -6048 1901
rect -5986 2819 -5952 2845
rect -5986 2811 -5952 2819
rect -5986 2751 -5952 2773
rect -5986 2739 -5952 2751
rect -5986 2683 -5952 2701
rect -5986 2667 -5952 2683
rect -5986 2615 -5952 2629
rect -5986 2595 -5952 2615
rect -5986 2547 -5952 2557
rect -5986 2523 -5952 2547
rect -5986 2479 -5952 2485
rect -5986 2451 -5952 2479
rect -5986 2411 -5952 2413
rect -5986 2379 -5952 2411
rect -5986 2309 -5952 2341
rect -5986 2307 -5952 2309
rect -5986 2241 -5952 2269
rect -5986 2235 -5952 2241
rect -5986 2173 -5952 2197
rect -5986 2163 -5952 2173
rect -5986 2105 -5952 2125
rect -5986 2091 -5952 2105
rect -5986 2037 -5952 2053
rect -5986 2019 -5952 2037
rect -5986 1969 -5952 1981
rect -5986 1947 -5952 1969
rect -5986 1901 -5952 1909
rect -5986 1875 -5952 1901
rect -5890 2819 -5856 2845
rect -5890 2811 -5856 2819
rect -5890 2751 -5856 2773
rect -5890 2739 -5856 2751
rect -5890 2683 -5856 2701
rect -5890 2667 -5856 2683
rect -5890 2615 -5856 2629
rect -5890 2595 -5856 2615
rect -5890 2547 -5856 2557
rect -5890 2523 -5856 2547
rect -5890 2479 -5856 2485
rect -5890 2451 -5856 2479
rect -5890 2411 -5856 2413
rect -5890 2379 -5856 2411
rect -5890 2309 -5856 2341
rect -5890 2307 -5856 2309
rect -5890 2241 -5856 2269
rect -5890 2235 -5856 2241
rect -5890 2173 -5856 2197
rect -5890 2163 -5856 2173
rect -5890 2105 -5856 2125
rect -5890 2091 -5856 2105
rect -5890 2037 -5856 2053
rect -5890 2019 -5856 2037
rect -5890 1969 -5856 1981
rect -5890 1947 -5856 1969
rect -5890 1901 -5856 1909
rect -5890 1875 -5856 1901
rect -5794 2819 -5760 2845
rect -5794 2811 -5760 2819
rect -5794 2751 -5760 2773
rect -5794 2739 -5760 2751
rect -5794 2683 -5760 2701
rect -5794 2667 -5760 2683
rect -5794 2615 -5760 2629
rect -5794 2595 -5760 2615
rect -5794 2547 -5760 2557
rect -5794 2523 -5760 2547
rect -5794 2479 -5760 2485
rect -5794 2451 -5760 2479
rect -5794 2411 -5760 2413
rect -5794 2379 -5760 2411
rect -5794 2309 -5760 2341
rect -5794 2307 -5760 2309
rect -5794 2241 -5760 2269
rect -5794 2235 -5760 2241
rect -5794 2173 -5760 2197
rect -5794 2163 -5760 2173
rect -5794 2105 -5760 2125
rect -5794 2091 -5760 2105
rect -5794 2037 -5760 2053
rect -5794 2019 -5760 2037
rect -5794 1969 -5760 1981
rect -5794 1947 -5760 1969
rect -5794 1901 -5760 1909
rect -5794 1875 -5760 1901
rect -5698 2819 -5664 2845
rect -5698 2811 -5664 2819
rect -5698 2751 -5664 2773
rect -5698 2739 -5664 2751
rect -5698 2683 -5664 2701
rect -5698 2667 -5664 2683
rect -5698 2615 -5664 2629
rect -5698 2595 -5664 2615
rect -5698 2547 -5664 2557
rect -5698 2523 -5664 2547
rect -5698 2479 -5664 2485
rect -5698 2451 -5664 2479
rect -5698 2411 -5664 2413
rect -5698 2379 -5664 2411
rect -5698 2309 -5664 2341
rect -5698 2307 -5664 2309
rect -5698 2241 -5664 2269
rect -5698 2235 -5664 2241
rect -5698 2173 -5664 2197
rect -5698 2163 -5664 2173
rect -5698 2105 -5664 2125
rect -5698 2091 -5664 2105
rect -5698 2037 -5664 2053
rect -5698 2019 -5664 2037
rect -5698 1969 -5664 1981
rect -5698 1947 -5664 1969
rect -5698 1901 -5664 1909
rect -5698 1875 -5664 1901
rect -5602 2819 -5568 2845
rect -5602 2811 -5568 2819
rect -5602 2751 -5568 2773
rect -5602 2739 -5568 2751
rect -5602 2683 -5568 2701
rect -5602 2667 -5568 2683
rect -5602 2615 -5568 2629
rect -5602 2595 -5568 2615
rect -5602 2547 -5568 2557
rect -5602 2523 -5568 2547
rect -5602 2479 -5568 2485
rect -5602 2451 -5568 2479
rect -5602 2411 -5568 2413
rect -5602 2379 -5568 2411
rect -5602 2309 -5568 2341
rect -5602 2307 -5568 2309
rect -5602 2241 -5568 2269
rect -5602 2235 -5568 2241
rect -5602 2173 -5568 2197
rect -5602 2163 -5568 2173
rect -5602 2105 -5568 2125
rect -5602 2091 -5568 2105
rect -5602 2037 -5568 2053
rect -5602 2019 -5568 2037
rect -5602 1969 -5568 1981
rect -5602 1947 -5568 1969
rect -5602 1901 -5568 1909
rect -5602 1875 -5568 1901
rect -5506 2819 -5472 2845
rect -5506 2811 -5472 2819
rect -5506 2751 -5472 2773
rect -5506 2739 -5472 2751
rect -5506 2683 -5472 2701
rect -5506 2667 -5472 2683
rect -5506 2615 -5472 2629
rect -5506 2595 -5472 2615
rect -5506 2547 -5472 2557
rect -5506 2523 -5472 2547
rect -5506 2479 -5472 2485
rect -5506 2451 -5472 2479
rect -5506 2411 -5472 2413
rect -5506 2379 -5472 2411
rect -5506 2309 -5472 2341
rect -5506 2307 -5472 2309
rect -5506 2241 -5472 2269
rect -5506 2235 -5472 2241
rect -5506 2173 -5472 2197
rect -5506 2163 -5472 2173
rect -5506 2105 -5472 2125
rect -5506 2091 -5472 2105
rect -5506 2037 -5472 2053
rect -5506 2019 -5472 2037
rect -5506 1969 -5472 1981
rect -5506 1947 -5472 1969
rect -5506 1901 -5472 1909
rect -5506 1875 -5472 1901
rect -5410 2819 -5376 2845
rect -5410 2811 -5376 2819
rect -5410 2751 -5376 2773
rect -5410 2739 -5376 2751
rect -5410 2683 -5376 2701
rect -5410 2667 -5376 2683
rect -5410 2615 -5376 2629
rect -5410 2595 -5376 2615
rect -5410 2547 -5376 2557
rect -5410 2523 -5376 2547
rect -5410 2479 -5376 2485
rect -5410 2451 -5376 2479
rect -5410 2411 -5376 2413
rect -5410 2379 -5376 2411
rect -5410 2309 -5376 2341
rect -5410 2307 -5376 2309
rect -5410 2241 -5376 2269
rect -5410 2235 -5376 2241
rect -5410 2173 -5376 2197
rect -5410 2163 -5376 2173
rect -5410 2105 -5376 2125
rect -5410 2091 -5376 2105
rect -5410 2037 -5376 2053
rect -5410 2019 -5376 2037
rect -5410 1969 -5376 1981
rect -5410 1947 -5376 1969
rect -5410 1901 -5376 1909
rect -5410 1875 -5376 1901
rect -5198 2829 -5164 2855
rect -5198 2821 -5164 2829
rect -5198 2761 -5164 2783
rect -5198 2749 -5164 2761
rect -5198 2693 -5164 2711
rect -5198 2677 -5164 2693
rect -5198 2625 -5164 2639
rect -5198 2605 -5164 2625
rect -5198 2557 -5164 2567
rect -5198 2533 -5164 2557
rect -5198 2489 -5164 2495
rect -5198 2461 -5164 2489
rect -5198 2421 -5164 2423
rect -5198 2389 -5164 2421
rect -5198 2319 -5164 2351
rect -5198 2317 -5164 2319
rect -5198 2251 -5164 2279
rect -5198 2245 -5164 2251
rect -5198 2183 -5164 2207
rect -5198 2173 -5164 2183
rect -5198 2115 -5164 2135
rect -5198 2101 -5164 2115
rect -5198 2047 -5164 2063
rect -5198 2029 -5164 2047
rect -5198 1979 -5164 1991
rect -5198 1957 -5164 1979
rect -5198 1911 -5164 1919
rect -5198 1885 -5164 1911
rect -5102 2829 -5068 2855
rect -5102 2821 -5068 2829
rect -5102 2761 -5068 2783
rect -5102 2749 -5068 2761
rect -5102 2693 -5068 2711
rect -5102 2677 -5068 2693
rect -5102 2625 -5068 2639
rect -5102 2605 -5068 2625
rect -5102 2557 -5068 2567
rect -5102 2533 -5068 2557
rect -5102 2489 -5068 2495
rect -5102 2461 -5068 2489
rect -5102 2421 -5068 2423
rect -5102 2389 -5068 2421
rect -5102 2319 -5068 2351
rect -5102 2317 -5068 2319
rect -5102 2251 -5068 2279
rect -5102 2245 -5068 2251
rect -5102 2183 -5068 2207
rect -5102 2173 -5068 2183
rect -5102 2115 -5068 2135
rect -5102 2101 -5068 2115
rect -5102 2047 -5068 2063
rect -5102 2029 -5068 2047
rect -5102 1979 -5068 1991
rect -5102 1957 -5068 1979
rect -5102 1911 -5068 1919
rect -5102 1885 -5068 1911
rect -5006 2829 -4972 2855
rect -5006 2821 -4972 2829
rect -5006 2761 -4972 2783
rect -5006 2749 -4972 2761
rect -5006 2693 -4972 2711
rect -5006 2677 -4972 2693
rect -5006 2625 -4972 2639
rect -5006 2605 -4972 2625
rect -5006 2557 -4972 2567
rect -5006 2533 -4972 2557
rect -5006 2489 -4972 2495
rect -5006 2461 -4972 2489
rect -5006 2421 -4972 2423
rect -5006 2389 -4972 2421
rect -5006 2319 -4972 2351
rect -5006 2317 -4972 2319
rect -5006 2251 -4972 2279
rect -5006 2245 -4972 2251
rect -5006 2183 -4972 2207
rect -5006 2173 -4972 2183
rect -5006 2115 -4972 2135
rect -5006 2101 -4972 2115
rect -5006 2047 -4972 2063
rect -5006 2029 -4972 2047
rect -5006 1979 -4972 1991
rect -5006 1957 -4972 1979
rect -5006 1911 -4972 1919
rect -5006 1885 -4972 1911
rect -4910 2829 -4876 2855
rect -4910 2821 -4876 2829
rect -4910 2761 -4876 2783
rect -4910 2749 -4876 2761
rect -4910 2693 -4876 2711
rect -4910 2677 -4876 2693
rect -4910 2625 -4876 2639
rect -4910 2605 -4876 2625
rect -4910 2557 -4876 2567
rect -4910 2533 -4876 2557
rect -4910 2489 -4876 2495
rect -4910 2461 -4876 2489
rect -4910 2421 -4876 2423
rect -4910 2389 -4876 2421
rect -4910 2319 -4876 2351
rect -4910 2317 -4876 2319
rect -4910 2251 -4876 2279
rect -4910 2245 -4876 2251
rect -4910 2183 -4876 2207
rect -4910 2173 -4876 2183
rect -4910 2115 -4876 2135
rect -4910 2101 -4876 2115
rect -4910 2047 -4876 2063
rect -4910 2029 -4876 2047
rect -4910 1979 -4876 1991
rect -4910 1957 -4876 1979
rect -4910 1911 -4876 1919
rect -4910 1885 -4876 1911
rect -1686 2923 -1652 2933
rect -1686 2899 -1652 2923
rect -4814 2829 -4780 2855
rect -4814 2821 -4780 2829
rect -4814 2761 -4780 2783
rect -4814 2749 -4780 2761
rect -4814 2693 -4780 2711
rect -4814 2677 -4780 2693
rect -4814 2625 -4780 2639
rect -4814 2605 -4780 2625
rect -4814 2557 -4780 2567
rect -4814 2533 -4780 2557
rect -4814 2489 -4780 2495
rect -4814 2461 -4780 2489
rect -4814 2421 -4780 2423
rect -4814 2389 -4780 2421
rect -4814 2319 -4780 2351
rect -4814 2317 -4780 2319
rect -4814 2251 -4780 2279
rect -4814 2245 -4780 2251
rect -4814 2183 -4780 2207
rect -4814 2173 -4780 2183
rect -4814 2115 -4780 2135
rect -4814 2101 -4780 2115
rect -4814 2047 -4780 2063
rect -4814 2029 -4780 2047
rect -4814 1979 -4780 1991
rect -4814 1957 -4780 1979
rect -4814 1911 -4780 1919
rect -4814 1885 -4780 1911
rect -4718 2829 -4684 2855
rect -4718 2821 -4684 2829
rect -4718 2761 -4684 2783
rect -4718 2749 -4684 2761
rect -4718 2693 -4684 2711
rect -4718 2677 -4684 2693
rect -4718 2625 -4684 2639
rect -4718 2605 -4684 2625
rect -4718 2557 -4684 2567
rect -4718 2533 -4684 2557
rect -4718 2489 -4684 2495
rect -4718 2461 -4684 2489
rect -4718 2421 -4684 2423
rect -4718 2389 -4684 2421
rect -4718 2319 -4684 2351
rect -4718 2317 -4684 2319
rect -4718 2251 -4684 2279
rect -4718 2245 -4684 2251
rect -4718 2183 -4684 2207
rect -4718 2173 -4684 2183
rect -1686 2855 -1652 2861
rect -1686 2827 -1652 2855
rect -1686 2787 -1652 2789
rect -1686 2755 -1652 2787
rect -1686 2685 -1652 2717
rect -1686 2683 -1652 2685
rect -1686 2617 -1652 2645
rect -1686 2611 -1652 2617
rect -1686 2549 -1652 2573
rect -1686 2539 -1652 2549
rect -1686 2481 -1652 2501
rect -1686 2467 -1652 2481
rect -1686 2413 -1652 2429
rect -1686 2395 -1652 2413
rect -1686 2345 -1652 2357
rect -1686 2323 -1652 2345
rect -1686 2277 -1652 2285
rect -1686 2251 -1652 2277
rect -1590 3195 -1556 3221
rect -1590 3187 -1556 3195
rect -1590 3127 -1556 3149
rect -1590 3115 -1556 3127
rect -1590 3059 -1556 3077
rect -1590 3043 -1556 3059
rect -1590 2991 -1556 3005
rect -1590 2971 -1556 2991
rect -1590 2923 -1556 2933
rect -1590 2899 -1556 2923
rect -1590 2855 -1556 2861
rect -1590 2827 -1556 2855
rect -1590 2787 -1556 2789
rect -1590 2755 -1556 2787
rect -1590 2685 -1556 2717
rect -1590 2683 -1556 2685
rect -1590 2617 -1556 2645
rect -1590 2611 -1556 2617
rect -1590 2549 -1556 2573
rect -1590 2539 -1556 2549
rect -1590 2481 -1556 2501
rect -1590 2467 -1556 2481
rect -1590 2413 -1556 2429
rect -1590 2395 -1556 2413
rect -1590 2345 -1556 2357
rect -1590 2323 -1556 2345
rect -1590 2277 -1556 2285
rect -1590 2251 -1556 2277
rect -1494 3195 -1460 3221
rect -1494 3187 -1460 3195
rect -1494 3127 -1460 3149
rect -1494 3115 -1460 3127
rect -1494 3059 -1460 3077
rect -1494 3043 -1460 3059
rect -1494 2991 -1460 3005
rect -1494 2971 -1460 2991
rect -1494 2923 -1460 2933
rect -1494 2899 -1460 2923
rect -1494 2855 -1460 2861
rect -1494 2827 -1460 2855
rect -1494 2787 -1460 2789
rect -1494 2755 -1460 2787
rect -1494 2685 -1460 2717
rect -1494 2683 -1460 2685
rect -1494 2617 -1460 2645
rect -1494 2611 -1460 2617
rect -1494 2549 -1460 2573
rect -1494 2539 -1460 2549
rect -1494 2481 -1460 2501
rect -1494 2467 -1460 2481
rect -1494 2413 -1460 2429
rect -1494 2395 -1460 2413
rect -1494 2345 -1460 2357
rect -1494 2323 -1460 2345
rect -1494 2277 -1460 2285
rect -1494 2251 -1460 2277
rect -1398 3195 -1364 3221
rect -1398 3187 -1364 3195
rect -1398 3127 -1364 3149
rect -1398 3115 -1364 3127
rect -1398 3059 -1364 3077
rect -1398 3043 -1364 3059
rect -1398 2991 -1364 3005
rect -1398 2971 -1364 2991
rect -1398 2923 -1364 2933
rect -1398 2899 -1364 2923
rect -1398 2855 -1364 2861
rect -1398 2827 -1364 2855
rect -1398 2787 -1364 2789
rect -1398 2755 -1364 2787
rect -1398 2685 -1364 2717
rect -1398 2683 -1364 2685
rect -1398 2617 -1364 2645
rect -1398 2611 -1364 2617
rect -1398 2549 -1364 2573
rect -1398 2539 -1364 2549
rect -1398 2481 -1364 2501
rect -1398 2467 -1364 2481
rect -1398 2413 -1364 2429
rect -1398 2395 -1364 2413
rect -1398 2345 -1364 2357
rect -1398 2323 -1364 2345
rect -1398 2277 -1364 2285
rect -1398 2251 -1364 2277
rect -1302 3195 -1268 3221
rect -1302 3187 -1268 3195
rect -1302 3127 -1268 3149
rect -1302 3115 -1268 3127
rect -1302 3059 -1268 3077
rect -1302 3043 -1268 3059
rect -1302 2991 -1268 3005
rect -1302 2971 -1268 2991
rect -1302 2923 -1268 2933
rect -1302 2899 -1268 2923
rect -1302 2855 -1268 2861
rect -1302 2827 -1268 2855
rect -1302 2787 -1268 2789
rect -1302 2755 -1268 2787
rect -1302 2685 -1268 2717
rect -1302 2683 -1268 2685
rect -1302 2617 -1268 2645
rect -1302 2611 -1268 2617
rect -1302 2549 -1268 2573
rect -1302 2539 -1268 2549
rect -1302 2481 -1268 2501
rect -1302 2467 -1268 2481
rect -1302 2413 -1268 2429
rect -1302 2395 -1268 2413
rect -1302 2345 -1268 2357
rect -1302 2323 -1268 2345
rect -1302 2277 -1268 2285
rect -1302 2251 -1268 2277
rect -1206 3195 -1172 3221
rect -1206 3187 -1172 3195
rect -1206 3127 -1172 3149
rect -1206 3115 -1172 3127
rect -1206 3059 -1172 3077
rect -1206 3043 -1172 3059
rect -1206 2991 -1172 3005
rect -1206 2971 -1172 2991
rect -1206 2923 -1172 2933
rect -1206 2899 -1172 2923
rect -1206 2855 -1172 2861
rect -1206 2827 -1172 2855
rect -1206 2787 -1172 2789
rect -1206 2755 -1172 2787
rect -1206 2685 -1172 2717
rect -1206 2683 -1172 2685
rect -1206 2617 -1172 2645
rect -1206 2611 -1172 2617
rect -1206 2549 -1172 2573
rect -1206 2539 -1172 2549
rect -1206 2481 -1172 2501
rect -1206 2467 -1172 2481
rect -1206 2413 -1172 2429
rect -1206 2395 -1172 2413
rect -1206 2345 -1172 2357
rect -1206 2323 -1172 2345
rect -1206 2277 -1172 2285
rect -1206 2251 -1172 2277
rect -1110 3195 -1076 3221
rect -1110 3187 -1076 3195
rect -1110 3127 -1076 3149
rect -1110 3115 -1076 3127
rect -1110 3059 -1076 3077
rect -1110 3043 -1076 3059
rect -1110 2991 -1076 3005
rect -1110 2971 -1076 2991
rect -1110 2923 -1076 2933
rect -1110 2899 -1076 2923
rect -1110 2855 -1076 2861
rect -1110 2827 -1076 2855
rect -1110 2787 -1076 2789
rect -1110 2755 -1076 2787
rect -1110 2685 -1076 2717
rect -1110 2683 -1076 2685
rect -1110 2617 -1076 2645
rect -1110 2611 -1076 2617
rect -1110 2549 -1076 2573
rect -1110 2539 -1076 2549
rect -1110 2481 -1076 2501
rect -1110 2467 -1076 2481
rect -1110 2413 -1076 2429
rect -1110 2395 -1076 2413
rect -1110 2345 -1076 2357
rect -1110 2323 -1076 2345
rect -1110 2277 -1076 2285
rect -1110 2251 -1076 2277
rect 16686 3289 16720 3303
rect 16686 3269 16720 3289
rect -1014 3195 -980 3221
rect -1014 3187 -980 3195
rect -1014 3127 -980 3149
rect -1014 3115 -980 3127
rect -1014 3059 -980 3077
rect -1014 3043 -980 3059
rect -1014 2991 -980 3005
rect -1014 2971 -980 2991
rect -1014 2923 -980 2933
rect -1014 2899 -980 2923
rect -1014 2855 -980 2861
rect -1014 2827 -980 2855
rect -1014 2787 -980 2789
rect -1014 2755 -980 2787
rect -1014 2685 -980 2717
rect -1014 2683 -980 2685
rect -1014 2617 -980 2645
rect -1014 2611 -980 2617
rect -1014 2549 -980 2573
rect -1014 2539 -980 2549
rect -1014 2481 -980 2501
rect -1014 2467 -980 2481
rect -1014 2413 -980 2429
rect -1014 2395 -980 2413
rect -1014 2345 -980 2357
rect -1014 2323 -980 2345
rect -1014 2277 -980 2285
rect -1014 2251 -980 2277
rect -918 3195 -884 3221
rect -918 3187 -884 3195
rect -918 3127 -884 3149
rect -918 3115 -884 3127
rect -918 3059 -884 3077
rect -918 3043 -884 3059
rect -918 2991 -884 3005
rect 16686 3221 16720 3231
rect 16686 3197 16720 3221
rect 16686 3153 16720 3159
rect 16686 3125 16720 3153
rect 16686 3085 16720 3087
rect 16686 3053 16720 3085
rect -918 2971 -884 2991
rect 1578 2968 1612 3002
rect -918 2923 -884 2933
rect -918 2899 -884 2923
rect 1674 2960 1708 2994
rect 4534 2952 4568 2986
rect 4630 2944 4664 2978
rect 7564 2952 7598 2986
rect -918 2855 -884 2861
rect -918 2827 -884 2855
rect 7660 2944 7694 2978
rect 10652 2950 10686 2984
rect 16686 2983 16720 3015
rect 16686 2981 16720 2983
rect 10748 2942 10782 2976
rect -918 2787 -884 2789
rect -918 2755 -884 2787
rect -918 2685 -884 2717
rect -918 2683 -884 2685
rect -918 2617 -884 2645
rect -918 2611 -884 2617
rect -918 2549 -884 2573
rect -918 2539 -884 2549
rect -918 2481 -884 2501
rect -918 2467 -884 2481
rect -918 2413 -884 2429
rect -918 2395 -884 2413
rect -918 2345 -884 2357
rect -918 2323 -884 2345
rect -918 2277 -884 2285
rect -918 2251 -884 2277
rect -1097 2138 -1063 2172
rect 1482 2789 1516 2815
rect 1482 2781 1516 2789
rect 1482 2721 1516 2743
rect 1482 2709 1516 2721
rect 1482 2653 1516 2671
rect 1482 2637 1516 2653
rect 1482 2585 1516 2599
rect 1482 2565 1516 2585
rect 1482 2517 1516 2527
rect 1482 2493 1516 2517
rect 1482 2449 1516 2455
rect 1482 2421 1516 2449
rect 1482 2381 1516 2383
rect 1482 2349 1516 2381
rect 1482 2279 1516 2311
rect 1482 2277 1516 2279
rect 1482 2211 1516 2239
rect 1482 2205 1516 2211
rect 1482 2143 1516 2167
rect -4718 2115 -4684 2135
rect -4718 2101 -4684 2115
rect -4718 2047 -4684 2063
rect -4718 2029 -4684 2047
rect -4718 1979 -4684 1991
rect -4718 1957 -4684 1979
rect -4718 1911 -4684 1919
rect -4718 1885 -4684 1911
rect 1482 2133 1516 2143
rect 1482 2075 1516 2095
rect 1482 2061 1516 2075
rect 1482 2007 1516 2023
rect 1482 1989 1516 2007
rect 1482 1939 1516 1951
rect 1482 1917 1516 1939
rect 1482 1871 1516 1879
rect 1482 1845 1516 1871
rect 1578 2789 1612 2815
rect 1578 2781 1612 2789
rect 1578 2721 1612 2743
rect 1578 2709 1612 2721
rect 1578 2653 1612 2671
rect 1578 2637 1612 2653
rect 1578 2585 1612 2599
rect 1578 2565 1612 2585
rect 1578 2517 1612 2527
rect 1578 2493 1612 2517
rect 1578 2449 1612 2455
rect 1578 2421 1612 2449
rect 1578 2381 1612 2383
rect 1578 2349 1612 2381
rect 1578 2279 1612 2311
rect 1578 2277 1612 2279
rect 1578 2211 1612 2239
rect 1578 2205 1612 2211
rect 1578 2143 1612 2167
rect 1578 2133 1612 2143
rect 1578 2075 1612 2095
rect 1578 2061 1612 2075
rect 1578 2007 1612 2023
rect 1578 1989 1612 2007
rect 1578 1939 1612 1951
rect 1578 1917 1612 1939
rect 1578 1871 1612 1879
rect 1578 1845 1612 1871
rect 1674 2789 1708 2815
rect 1674 2781 1708 2789
rect 1674 2721 1708 2743
rect 1674 2709 1708 2721
rect 1674 2653 1708 2671
rect 1674 2637 1708 2653
rect 1674 2585 1708 2599
rect 1674 2565 1708 2585
rect 1674 2517 1708 2527
rect 1674 2493 1708 2517
rect 1674 2449 1708 2455
rect 1674 2421 1708 2449
rect 1674 2381 1708 2383
rect 1674 2349 1708 2381
rect 1674 2279 1708 2311
rect 1674 2277 1708 2279
rect 1674 2211 1708 2239
rect 1674 2205 1708 2211
rect 1674 2143 1708 2167
rect 1674 2133 1708 2143
rect 1674 2075 1708 2095
rect 1674 2061 1708 2075
rect 1674 2007 1708 2023
rect 1674 1989 1708 2007
rect 1674 1939 1708 1951
rect 1674 1917 1708 1939
rect 1674 1871 1708 1879
rect 1674 1845 1708 1871
rect 1770 2789 1804 2815
rect 1770 2781 1804 2789
rect 1770 2721 1804 2743
rect 1770 2709 1804 2721
rect 1770 2653 1804 2671
rect 1770 2637 1804 2653
rect 1770 2585 1804 2599
rect 1770 2565 1804 2585
rect 1770 2517 1804 2527
rect 1770 2493 1804 2517
rect 1770 2449 1804 2455
rect 1770 2421 1804 2449
rect 1770 2381 1804 2383
rect 1770 2349 1804 2381
rect 1770 2279 1804 2311
rect 1770 2277 1804 2279
rect 1770 2211 1804 2239
rect 1770 2205 1804 2211
rect 1770 2143 1804 2167
rect 1770 2133 1804 2143
rect 1770 2075 1804 2095
rect 1770 2061 1804 2075
rect 1770 2007 1804 2023
rect 1770 1989 1804 2007
rect 1770 1939 1804 1951
rect 1770 1917 1804 1939
rect 1770 1871 1804 1879
rect 1770 1845 1804 1871
rect 1866 2789 1900 2815
rect 1866 2781 1900 2789
rect 1866 2721 1900 2743
rect 1866 2709 1900 2721
rect 1866 2653 1900 2671
rect 1866 2637 1900 2653
rect 1866 2585 1900 2599
rect 1866 2565 1900 2585
rect 1866 2517 1900 2527
rect 1866 2493 1900 2517
rect 1866 2449 1900 2455
rect 1866 2421 1900 2449
rect 4438 2773 4472 2799
rect 4438 2765 4472 2773
rect 4438 2705 4472 2727
rect 4438 2693 4472 2705
rect 4438 2637 4472 2655
rect 4438 2621 4472 2637
rect 4438 2569 4472 2583
rect 4438 2549 4472 2569
rect 4438 2501 4472 2511
rect 4438 2477 4472 2501
rect 4438 2433 4472 2439
rect 2579 2394 2613 2428
rect 4438 2405 4472 2433
rect 1866 2381 1900 2383
rect 1866 2349 1900 2381
rect 4438 2365 4472 2367
rect 2392 2316 2426 2350
rect 1866 2279 1900 2311
rect 1866 2277 1900 2279
rect 1866 2211 1900 2239
rect 1866 2205 1900 2211
rect 1866 2143 1900 2167
rect 1866 2133 1900 2143
rect 1866 2075 1900 2095
rect 1866 2061 1900 2075
rect 1866 2007 1900 2023
rect 1866 1989 1900 2007
rect 1866 1939 1900 1951
rect 1866 1917 1900 1939
rect 2500 2227 2534 2229
rect 2500 2195 2534 2227
rect 2500 2125 2534 2157
rect 2500 2123 2534 2125
rect 2658 2227 2692 2229
rect 2658 2195 2692 2227
rect 2658 2125 2692 2157
rect 2658 2123 2692 2125
rect 4438 2333 4472 2365
rect 4438 2263 4472 2295
rect 4438 2261 4472 2263
rect 4438 2195 4472 2223
rect 4438 2189 4472 2195
rect 4438 2127 4472 2151
rect 4438 2117 4472 2127
rect 1866 1871 1900 1879
rect 1866 1845 1900 1871
rect 4438 2059 4472 2079
rect 4438 2045 4472 2059
rect 4438 1991 4472 2007
rect 4438 1973 4472 1991
rect 4438 1923 4472 1935
rect 4438 1901 4472 1923
rect -23029 1522 -22851 1628
rect -21034 1516 -20856 1622
rect -19026 1525 -18848 1631
rect -16546 1533 -16368 1639
rect -14350 1530 -14172 1636
rect -11944 1535 -11766 1641
rect -9379 1531 -9129 1637
rect -7345 1530 -7167 1636
rect -5345 1532 -5167 1638
rect 1578 1662 1612 1696
rect 4438 1855 4472 1863
rect 4438 1829 4472 1855
rect 4534 2773 4568 2799
rect 4534 2765 4568 2773
rect 4534 2705 4568 2727
rect 4534 2693 4568 2705
rect 4534 2637 4568 2655
rect 4534 2621 4568 2637
rect 4534 2569 4568 2583
rect 4534 2549 4568 2569
rect 4534 2501 4568 2511
rect 4534 2477 4568 2501
rect 4534 2433 4568 2439
rect 4534 2405 4568 2433
rect 4534 2365 4568 2367
rect 4534 2333 4568 2365
rect 4534 2263 4568 2295
rect 4534 2261 4568 2263
rect 4534 2195 4568 2223
rect 4534 2189 4568 2195
rect 4534 2127 4568 2151
rect 4534 2117 4568 2127
rect 4534 2059 4568 2079
rect 4534 2045 4568 2059
rect 4534 1991 4568 2007
rect 4534 1973 4568 1991
rect 4534 1923 4568 1935
rect 4534 1901 4568 1923
rect 4534 1855 4568 1863
rect 4534 1829 4568 1855
rect 4630 2773 4664 2799
rect 4630 2765 4664 2773
rect 4630 2705 4664 2727
rect 4630 2693 4664 2705
rect 4630 2637 4664 2655
rect 4630 2621 4664 2637
rect 4630 2569 4664 2583
rect 4630 2549 4664 2569
rect 4630 2501 4664 2511
rect 4630 2477 4664 2501
rect 4630 2433 4664 2439
rect 4630 2405 4664 2433
rect 4630 2365 4664 2367
rect 4630 2333 4664 2365
rect 4630 2263 4664 2295
rect 4630 2261 4664 2263
rect 4630 2195 4664 2223
rect 4630 2189 4664 2195
rect 4630 2127 4664 2151
rect 4630 2117 4664 2127
rect 4630 2059 4664 2079
rect 4630 2045 4664 2059
rect 4630 1991 4664 2007
rect 4630 1973 4664 1991
rect 4630 1923 4664 1935
rect 4630 1901 4664 1923
rect 4630 1855 4664 1863
rect 4630 1829 4664 1855
rect 13808 2924 13842 2958
rect 13904 2916 13938 2950
rect 4726 2773 4760 2799
rect 4726 2765 4760 2773
rect 4726 2705 4760 2727
rect 4726 2693 4760 2705
rect 4726 2637 4760 2655
rect 4726 2621 4760 2637
rect 4726 2569 4760 2583
rect 4726 2549 4760 2569
rect 4726 2501 4760 2511
rect 4726 2477 4760 2501
rect 4726 2433 4760 2439
rect 4726 2405 4760 2433
rect 4726 2365 4760 2367
rect 4726 2333 4760 2365
rect 4726 2263 4760 2295
rect 4726 2261 4760 2263
rect 4726 2195 4760 2223
rect 4726 2189 4760 2195
rect 4726 2127 4760 2151
rect 4726 2117 4760 2127
rect 4726 2059 4760 2079
rect 4726 2045 4760 2059
rect 4726 1991 4760 2007
rect 4726 1973 4760 1991
rect 4726 1923 4760 1935
rect 4726 1901 4760 1923
rect 4726 1855 4760 1863
rect 4726 1829 4760 1855
rect 4822 2773 4856 2799
rect 4822 2765 4856 2773
rect 4822 2705 4856 2727
rect 4822 2693 4856 2705
rect 4822 2637 4856 2655
rect 4822 2621 4856 2637
rect 4822 2569 4856 2583
rect 4822 2549 4856 2569
rect 4822 2501 4856 2511
rect 4822 2477 4856 2501
rect 4822 2433 4856 2439
rect 4822 2405 4856 2433
rect 7468 2773 7502 2799
rect 7468 2765 7502 2773
rect 7468 2705 7502 2727
rect 7468 2693 7502 2705
rect 7468 2637 7502 2655
rect 7468 2621 7502 2637
rect 7468 2569 7502 2583
rect 7468 2549 7502 2569
rect 7468 2501 7502 2511
rect 7468 2477 7502 2501
rect 7468 2433 7502 2439
rect 5579 2394 5613 2428
rect 7468 2405 7502 2433
rect 4822 2365 4856 2367
rect 4822 2333 4856 2365
rect 7468 2365 7502 2367
rect 5392 2316 5426 2350
rect 4822 2263 4856 2295
rect 4822 2261 4856 2263
rect 4822 2195 4856 2223
rect 4822 2189 4856 2195
rect 4822 2127 4856 2151
rect 4822 2117 4856 2127
rect 4822 2059 4856 2079
rect 4822 2045 4856 2059
rect 4822 1991 4856 2007
rect 4822 1973 4856 1991
rect 4822 1923 4856 1935
rect 4822 1901 4856 1923
rect 4822 1855 4856 1863
rect 4822 1829 4856 1855
rect 5500 2227 5534 2229
rect 5500 2195 5534 2227
rect 5500 2125 5534 2157
rect 5500 2123 5534 2125
rect 5658 2227 5692 2229
rect 5658 2195 5692 2227
rect 5658 2125 5692 2157
rect 5658 2123 5692 2125
rect 7468 2333 7502 2365
rect 7468 2263 7502 2295
rect 7468 2261 7502 2263
rect 7468 2195 7502 2223
rect 7468 2189 7502 2195
rect 7468 2127 7502 2151
rect 7468 2117 7502 2127
rect 7468 2059 7502 2079
rect 7468 2045 7502 2059
rect 7468 1991 7502 2007
rect 7468 1973 7502 1991
rect 7468 1923 7502 1935
rect 7468 1901 7502 1923
rect 7468 1855 7502 1863
rect 7468 1829 7502 1855
rect 7564 2773 7598 2799
rect 7564 2765 7598 2773
rect 7564 2705 7598 2727
rect 7564 2693 7598 2705
rect 7564 2637 7598 2655
rect 7564 2621 7598 2637
rect 7564 2569 7598 2583
rect 7564 2549 7598 2569
rect 7564 2501 7598 2511
rect 7564 2477 7598 2501
rect 7564 2433 7598 2439
rect 7564 2405 7598 2433
rect 7564 2365 7598 2367
rect 7564 2333 7598 2365
rect 7564 2263 7598 2295
rect 7564 2261 7598 2263
rect 7564 2195 7598 2223
rect 7564 2189 7598 2195
rect 7564 2127 7598 2151
rect 7564 2117 7598 2127
rect 7564 2059 7598 2079
rect 7564 2045 7598 2059
rect 7564 1991 7598 2007
rect 7564 1973 7598 1991
rect 7564 1923 7598 1935
rect 7564 1901 7598 1923
rect 7564 1855 7598 1863
rect 7564 1829 7598 1855
rect 7660 2773 7694 2799
rect 7660 2765 7694 2773
rect 7660 2705 7694 2727
rect 7660 2693 7694 2705
rect 7660 2637 7694 2655
rect 7660 2621 7694 2637
rect 7660 2569 7694 2583
rect 7660 2549 7694 2569
rect 7660 2501 7694 2511
rect 7660 2477 7694 2501
rect 7660 2433 7694 2439
rect 7660 2405 7694 2433
rect 7660 2365 7694 2367
rect 7660 2333 7694 2365
rect 7660 2263 7694 2295
rect 7660 2261 7694 2263
rect 7660 2195 7694 2223
rect 7660 2189 7694 2195
rect 7660 2127 7694 2151
rect 7660 2117 7694 2127
rect 7660 2059 7694 2079
rect 7660 2045 7694 2059
rect 7660 1991 7694 2007
rect 7660 1973 7694 1991
rect 7660 1923 7694 1935
rect 7660 1901 7694 1923
rect 7660 1855 7694 1863
rect 7660 1829 7694 1855
rect 16686 2915 16720 2943
rect 16686 2909 16720 2915
rect 7756 2773 7790 2799
rect 7756 2765 7790 2773
rect 7756 2705 7790 2727
rect 7756 2693 7790 2705
rect 7756 2637 7790 2655
rect 7756 2621 7790 2637
rect 7756 2569 7790 2583
rect 7756 2549 7790 2569
rect 7756 2501 7790 2511
rect 7756 2477 7790 2501
rect 7756 2433 7790 2439
rect 7756 2405 7790 2433
rect 7756 2365 7790 2367
rect 7756 2333 7790 2365
rect 7756 2263 7790 2295
rect 7756 2261 7790 2263
rect 7756 2195 7790 2223
rect 7756 2189 7790 2195
rect 7756 2127 7790 2151
rect 7756 2117 7790 2127
rect 7756 2059 7790 2079
rect 7756 2045 7790 2059
rect 7756 1991 7790 2007
rect 7756 1973 7790 1991
rect 7756 1923 7790 1935
rect 7756 1901 7790 1923
rect 7756 1855 7790 1863
rect 7756 1829 7790 1855
rect 7852 2773 7886 2799
rect 7852 2765 7886 2773
rect 7852 2705 7886 2727
rect 7852 2693 7886 2705
rect 7852 2637 7886 2655
rect 7852 2621 7886 2637
rect 7852 2569 7886 2583
rect 7852 2549 7886 2569
rect 7852 2501 7886 2511
rect 7852 2477 7886 2501
rect 7852 2433 7886 2439
rect 7852 2405 7886 2433
rect 10556 2771 10590 2797
rect 10556 2763 10590 2771
rect 10556 2703 10590 2725
rect 10556 2691 10590 2703
rect 10556 2635 10590 2653
rect 10556 2619 10590 2635
rect 10556 2567 10590 2581
rect 10556 2547 10590 2567
rect 10556 2499 10590 2509
rect 10556 2475 10590 2499
rect 10556 2431 10590 2437
rect 8579 2394 8613 2428
rect 10556 2403 10590 2431
rect 7852 2365 7886 2367
rect 7852 2333 7886 2365
rect 10556 2363 10590 2365
rect 8392 2316 8426 2350
rect 7852 2263 7886 2295
rect 7852 2261 7886 2263
rect 7852 2195 7886 2223
rect 7852 2189 7886 2195
rect 7852 2127 7886 2151
rect 7852 2117 7886 2127
rect 7852 2059 7886 2079
rect 7852 2045 7886 2059
rect 7852 1991 7886 2007
rect 7852 1973 7886 1991
rect 7852 1923 7886 1935
rect 7852 1901 7886 1923
rect 7852 1855 7886 1863
rect 7852 1829 7886 1855
rect 8500 2227 8534 2229
rect 8500 2195 8534 2227
rect 8500 2125 8534 2157
rect 8500 2123 8534 2125
rect 8658 2227 8692 2229
rect 8658 2195 8692 2227
rect 8658 2125 8692 2157
rect 8658 2123 8692 2125
rect 10556 2331 10590 2363
rect 10556 2261 10590 2293
rect 10556 2259 10590 2261
rect 10556 2193 10590 2221
rect 10556 2187 10590 2193
rect 10556 2125 10590 2149
rect 10556 2115 10590 2125
rect 4534 1646 4568 1680
rect 10556 2057 10590 2077
rect 10556 2043 10590 2057
rect 10556 1989 10590 2005
rect 10556 1971 10590 1989
rect 10556 1921 10590 1933
rect 10556 1899 10590 1921
rect 10556 1853 10590 1861
rect 10556 1827 10590 1853
rect 7564 1646 7598 1680
rect 10652 2771 10686 2797
rect 10652 2763 10686 2771
rect 10652 2703 10686 2725
rect 10652 2691 10686 2703
rect 10652 2635 10686 2653
rect 10652 2619 10686 2635
rect 10652 2567 10686 2581
rect 10652 2547 10686 2567
rect 10652 2499 10686 2509
rect 10652 2475 10686 2499
rect 10652 2431 10686 2437
rect 10652 2403 10686 2431
rect 10652 2363 10686 2365
rect 10652 2331 10686 2363
rect 10652 2261 10686 2293
rect 10652 2259 10686 2261
rect 10652 2193 10686 2221
rect 10652 2187 10686 2193
rect 10652 2125 10686 2149
rect 10652 2115 10686 2125
rect 10652 2057 10686 2077
rect 10652 2043 10686 2057
rect 10652 1989 10686 2005
rect 10652 1971 10686 1989
rect 10652 1921 10686 1933
rect 10652 1899 10686 1921
rect 10652 1853 10686 1861
rect 10652 1827 10686 1853
rect 10748 2771 10782 2797
rect 10748 2763 10782 2771
rect 10748 2703 10782 2725
rect 10748 2691 10782 2703
rect 10748 2635 10782 2653
rect 10748 2619 10782 2635
rect 10748 2567 10782 2581
rect 10748 2547 10782 2567
rect 10748 2499 10782 2509
rect 10748 2475 10782 2499
rect 10748 2431 10782 2437
rect 10748 2403 10782 2431
rect 10748 2363 10782 2365
rect 10748 2331 10782 2363
rect 10748 2261 10782 2293
rect 10748 2259 10782 2261
rect 10748 2193 10782 2221
rect 10748 2187 10782 2193
rect 10748 2125 10782 2149
rect 10748 2115 10782 2125
rect 10748 2057 10782 2077
rect 10748 2043 10782 2057
rect 10748 1989 10782 2005
rect 10748 1971 10782 1989
rect 10748 1921 10782 1933
rect 10748 1899 10782 1921
rect 10748 1853 10782 1861
rect 10748 1827 10782 1853
rect 10844 2771 10878 2797
rect 10844 2763 10878 2771
rect 10844 2703 10878 2725
rect 10844 2691 10878 2703
rect 10844 2635 10878 2653
rect 10844 2619 10878 2635
rect 10844 2567 10878 2581
rect 10844 2547 10878 2567
rect 10844 2499 10878 2509
rect 10844 2475 10878 2499
rect 10844 2431 10878 2437
rect 10844 2403 10878 2431
rect 10844 2363 10878 2365
rect 10844 2331 10878 2363
rect 10844 2261 10878 2293
rect 10844 2259 10878 2261
rect 10844 2193 10878 2221
rect 10844 2187 10878 2193
rect 10844 2125 10878 2149
rect 10844 2115 10878 2125
rect 10844 2057 10878 2077
rect 10844 2043 10878 2057
rect 10844 1989 10878 2005
rect 10844 1971 10878 1989
rect 10844 1921 10878 1933
rect 10844 1899 10878 1921
rect 10844 1853 10878 1861
rect 10844 1827 10878 1853
rect 10940 2771 10974 2797
rect 10940 2763 10974 2771
rect 10940 2703 10974 2725
rect 10940 2691 10974 2703
rect 10940 2635 10974 2653
rect 10940 2619 10974 2635
rect 10940 2567 10974 2581
rect 10940 2547 10974 2567
rect 10940 2499 10974 2509
rect 10940 2475 10974 2499
rect 10940 2431 10974 2437
rect 10940 2403 10974 2431
rect 13712 2745 13746 2771
rect 13712 2737 13746 2745
rect 13712 2677 13746 2699
rect 13712 2665 13746 2677
rect 13712 2609 13746 2627
rect 13712 2593 13746 2609
rect 13712 2541 13746 2555
rect 13712 2521 13746 2541
rect 13712 2473 13746 2483
rect 13712 2449 13746 2473
rect 11579 2394 11613 2428
rect 13712 2405 13746 2411
rect 10940 2363 10974 2365
rect 10940 2331 10974 2363
rect 13712 2377 13746 2405
rect 11392 2316 11426 2350
rect 10940 2261 10974 2293
rect 10940 2259 10974 2261
rect 10940 2193 10974 2221
rect 10940 2187 10974 2193
rect 10940 2125 10974 2149
rect 10940 2115 10974 2125
rect 10940 2057 10974 2077
rect 10940 2043 10974 2057
rect 10940 1989 10974 2005
rect 10940 1971 10974 1989
rect 10940 1921 10974 1933
rect 10940 1899 10974 1921
rect 10940 1853 10974 1861
rect 10940 1827 10974 1853
rect 11500 2227 11534 2229
rect 11500 2195 11534 2227
rect 11500 2125 11534 2157
rect 11500 2123 11534 2125
rect 11658 2227 11692 2229
rect 11658 2195 11692 2227
rect 11658 2125 11692 2157
rect 11658 2123 11692 2125
rect 13712 2337 13746 2339
rect 13712 2305 13746 2337
rect 13712 2235 13746 2267
rect 13712 2233 13746 2235
rect 13712 2167 13746 2195
rect 13712 2161 13746 2167
rect 13712 2099 13746 2123
rect 13712 2089 13746 2099
rect 13712 2031 13746 2051
rect 13712 2017 13746 2031
rect 13712 1963 13746 1979
rect 13712 1945 13746 1963
rect 13712 1895 13746 1907
rect 13712 1873 13746 1895
rect 13712 1827 13746 1835
rect 13712 1801 13746 1827
rect 13808 2745 13842 2771
rect 13808 2737 13842 2745
rect 13808 2677 13842 2699
rect 13808 2665 13842 2677
rect 13808 2609 13842 2627
rect 13808 2593 13842 2609
rect 13808 2541 13842 2555
rect 13808 2521 13842 2541
rect 13808 2473 13842 2483
rect 13808 2449 13842 2473
rect 13808 2405 13842 2411
rect 13808 2377 13842 2405
rect 13808 2337 13842 2339
rect 13808 2305 13842 2337
rect 13808 2235 13842 2267
rect 13808 2233 13842 2235
rect 13808 2167 13842 2195
rect 13808 2161 13842 2167
rect 13808 2099 13842 2123
rect 13808 2089 13842 2099
rect 13808 2031 13842 2051
rect 13808 2017 13842 2031
rect 13808 1963 13842 1979
rect 13808 1945 13842 1963
rect 13808 1895 13842 1907
rect 13808 1873 13842 1895
rect 13808 1827 13842 1835
rect 13808 1801 13842 1827
rect 13904 2745 13938 2771
rect 13904 2737 13938 2745
rect 13904 2677 13938 2699
rect 13904 2665 13938 2677
rect 13904 2609 13938 2627
rect 13904 2593 13938 2609
rect 13904 2541 13938 2555
rect 13904 2521 13938 2541
rect 13904 2473 13938 2483
rect 13904 2449 13938 2473
rect 13904 2405 13938 2411
rect 13904 2377 13938 2405
rect 13904 2337 13938 2339
rect 13904 2305 13938 2337
rect 13904 2235 13938 2267
rect 13904 2233 13938 2235
rect 13904 2167 13938 2195
rect 13904 2161 13938 2167
rect 13904 2099 13938 2123
rect 13904 2089 13938 2099
rect 13904 2031 13938 2051
rect 13904 2017 13938 2031
rect 13904 1963 13938 1979
rect 13904 1945 13938 1963
rect 13904 1895 13938 1907
rect 13904 1873 13938 1895
rect 13904 1827 13938 1835
rect 13904 1801 13938 1827
rect 16686 2847 16720 2871
rect 16686 2837 16720 2847
rect 14000 2745 14034 2771
rect 14000 2737 14034 2745
rect 14000 2677 14034 2699
rect 14000 2665 14034 2677
rect 14000 2609 14034 2627
rect 14000 2593 14034 2609
rect 14000 2541 14034 2555
rect 14000 2521 14034 2541
rect 14000 2473 14034 2483
rect 14000 2449 14034 2473
rect 14000 2405 14034 2411
rect 14000 2377 14034 2405
rect 14000 2337 14034 2339
rect 14000 2305 14034 2337
rect 14000 2235 14034 2267
rect 14000 2233 14034 2235
rect 14000 2167 14034 2195
rect 14000 2161 14034 2167
rect 14000 2099 14034 2123
rect 14000 2089 14034 2099
rect 14000 2031 14034 2051
rect 14000 2017 14034 2031
rect 14000 1963 14034 1979
rect 14000 1945 14034 1963
rect 14000 1895 14034 1907
rect 14000 1873 14034 1895
rect 14000 1827 14034 1835
rect 14000 1801 14034 1827
rect 14096 2745 14130 2771
rect 14096 2737 14130 2745
rect 14096 2677 14130 2699
rect 14096 2665 14130 2677
rect 14096 2609 14130 2627
rect 14096 2593 14130 2609
rect 14096 2541 14130 2555
rect 14096 2521 14130 2541
rect 14096 2473 14130 2483
rect 14096 2449 14130 2473
rect 16686 2779 16720 2799
rect 16686 2765 16720 2779
rect 16686 2711 16720 2727
rect 16686 2693 16720 2711
rect 16686 2643 16720 2655
rect 16686 2621 16720 2643
rect 16686 2575 16720 2583
rect 16686 2549 16720 2575
rect 16782 3493 16816 3519
rect 16782 3485 16816 3493
rect 16782 3425 16816 3447
rect 16782 3413 16816 3425
rect 16782 3357 16816 3375
rect 16782 3341 16816 3357
rect 16782 3289 16816 3303
rect 16782 3269 16816 3289
rect 16782 3221 16816 3231
rect 16782 3197 16816 3221
rect 16782 3153 16816 3159
rect 16782 3125 16816 3153
rect 16782 3085 16816 3087
rect 16782 3053 16816 3085
rect 16782 2983 16816 3015
rect 16782 2981 16816 2983
rect 16782 2915 16816 2943
rect 16782 2909 16816 2915
rect 16782 2847 16816 2871
rect 16782 2837 16816 2847
rect 16782 2779 16816 2799
rect 16782 2765 16816 2779
rect 16782 2711 16816 2727
rect 16782 2693 16816 2711
rect 16782 2643 16816 2655
rect 16782 2621 16816 2643
rect 16782 2575 16816 2583
rect 16782 2549 16816 2575
rect 16878 3493 16912 3519
rect 16878 3485 16912 3493
rect 16878 3425 16912 3447
rect 16878 3413 16912 3425
rect 16878 3357 16912 3375
rect 16878 3341 16912 3357
rect 16878 3289 16912 3303
rect 16878 3269 16912 3289
rect 16878 3221 16912 3231
rect 16878 3197 16912 3221
rect 16878 3153 16912 3159
rect 16878 3125 16912 3153
rect 16878 3085 16912 3087
rect 16878 3053 16912 3085
rect 16878 2983 16912 3015
rect 16878 2981 16912 2983
rect 16878 2915 16912 2943
rect 16878 2909 16912 2915
rect 16878 2847 16912 2871
rect 16878 2837 16912 2847
rect 16878 2779 16912 2799
rect 16878 2765 16912 2779
rect 16878 2711 16912 2727
rect 16878 2693 16912 2711
rect 16878 2643 16912 2655
rect 16878 2621 16912 2643
rect 16878 2575 16912 2583
rect 16878 2549 16912 2575
rect 16974 3493 17008 3519
rect 16974 3485 17008 3493
rect 16974 3425 17008 3447
rect 16974 3413 17008 3425
rect 16974 3357 17008 3375
rect 16974 3341 17008 3357
rect 16974 3289 17008 3303
rect 16974 3269 17008 3289
rect 16974 3221 17008 3231
rect 16974 3197 17008 3221
rect 16974 3153 17008 3159
rect 16974 3125 17008 3153
rect 16974 3085 17008 3087
rect 16974 3053 17008 3085
rect 16974 2983 17008 3015
rect 16974 2981 17008 2983
rect 16974 2915 17008 2943
rect 16974 2909 17008 2915
rect 16974 2847 17008 2871
rect 16974 2837 17008 2847
rect 16974 2779 17008 2799
rect 16974 2765 17008 2779
rect 16974 2711 17008 2727
rect 16974 2693 17008 2711
rect 16974 2643 17008 2655
rect 16974 2621 17008 2643
rect 16974 2575 17008 2583
rect 16974 2549 17008 2575
rect 17070 3493 17104 3519
rect 17070 3485 17104 3493
rect 17070 3425 17104 3447
rect 17070 3413 17104 3425
rect 17070 3357 17104 3375
rect 17070 3341 17104 3357
rect 17070 3289 17104 3303
rect 17070 3269 17104 3289
rect 17070 3221 17104 3231
rect 17070 3197 17104 3221
rect 17070 3153 17104 3159
rect 17070 3125 17104 3153
rect 17070 3085 17104 3087
rect 17070 3053 17104 3085
rect 17070 2983 17104 3015
rect 17070 2981 17104 2983
rect 17070 2915 17104 2943
rect 17070 2909 17104 2915
rect 17070 2847 17104 2871
rect 17070 2837 17104 2847
rect 17070 2779 17104 2799
rect 17070 2765 17104 2779
rect 17070 2711 17104 2727
rect 17070 2693 17104 2711
rect 17070 2643 17104 2655
rect 17070 2621 17104 2643
rect 17070 2575 17104 2583
rect 17070 2549 17104 2575
rect 23318 3907 23352 3941
rect 21646 3770 21680 3804
rect 20388 3656 20422 3690
rect 17166 3493 17200 3519
rect 17166 3485 17200 3493
rect 17166 3425 17200 3447
rect 17166 3413 17200 3425
rect 17166 3357 17200 3375
rect 17166 3341 17200 3357
rect 17166 3289 17200 3303
rect 17166 3269 17200 3289
rect 17166 3221 17200 3231
rect 17166 3197 17200 3221
rect 17166 3153 17200 3159
rect 17166 3125 17200 3153
rect 17166 3085 17200 3087
rect 17166 3053 17200 3085
rect 17166 2983 17200 3015
rect 17166 2981 17200 2983
rect 17166 2915 17200 2943
rect 17166 2909 17200 2915
rect 17166 2847 17200 2871
rect 17166 2837 17200 2847
rect 17166 2779 17200 2799
rect 17166 2765 17200 2779
rect 17166 2711 17200 2727
rect 17166 2693 17200 2711
rect 17166 2643 17200 2655
rect 17166 2621 17200 2643
rect 17166 2575 17200 2583
rect 17166 2549 17200 2575
rect 17378 3483 17412 3509
rect 17378 3475 17412 3483
rect 17378 3415 17412 3437
rect 17378 3403 17412 3415
rect 17378 3347 17412 3365
rect 17378 3331 17412 3347
rect 17378 3279 17412 3293
rect 17378 3259 17412 3279
rect 17378 3211 17412 3221
rect 17378 3187 17412 3211
rect 17378 3143 17412 3149
rect 17378 3115 17412 3143
rect 17378 3075 17412 3077
rect 17378 3043 17412 3075
rect 17378 2973 17412 3005
rect 17378 2971 17412 2973
rect 17378 2905 17412 2933
rect 17378 2899 17412 2905
rect 17378 2837 17412 2861
rect 17378 2827 17412 2837
rect 17378 2769 17412 2789
rect 17378 2755 17412 2769
rect 17378 2701 17412 2717
rect 17378 2683 17412 2701
rect 17378 2633 17412 2645
rect 17378 2611 17412 2633
rect 17378 2565 17412 2573
rect 17378 2539 17412 2565
rect 17474 3483 17508 3509
rect 17474 3475 17508 3483
rect 17474 3415 17508 3437
rect 17474 3403 17508 3415
rect 17474 3347 17508 3365
rect 17474 3331 17508 3347
rect 17474 3279 17508 3293
rect 17474 3259 17508 3279
rect 17474 3211 17508 3221
rect 17474 3187 17508 3211
rect 17474 3143 17508 3149
rect 17474 3115 17508 3143
rect 17474 3075 17508 3077
rect 17474 3043 17508 3075
rect 17474 2973 17508 3005
rect 17474 2971 17508 2973
rect 17474 2905 17508 2933
rect 17474 2899 17508 2905
rect 17474 2837 17508 2861
rect 17474 2827 17508 2837
rect 17474 2769 17508 2789
rect 17474 2755 17508 2769
rect 17474 2701 17508 2717
rect 17474 2683 17508 2701
rect 17474 2633 17508 2645
rect 17474 2611 17508 2633
rect 17474 2565 17508 2573
rect 17474 2539 17508 2565
rect 17570 3483 17604 3509
rect 17570 3475 17604 3483
rect 17570 3415 17604 3437
rect 17570 3403 17604 3415
rect 17570 3347 17604 3365
rect 17570 3331 17604 3347
rect 17570 3279 17604 3293
rect 17570 3259 17604 3279
rect 17570 3211 17604 3221
rect 17570 3187 17604 3211
rect 17570 3143 17604 3149
rect 17570 3115 17604 3143
rect 17570 3075 17604 3077
rect 17570 3043 17604 3075
rect 17570 2973 17604 3005
rect 17570 2971 17604 2973
rect 17570 2905 17604 2933
rect 17570 2899 17604 2905
rect 17570 2837 17604 2861
rect 17570 2827 17604 2837
rect 17570 2769 17604 2789
rect 17570 2755 17604 2769
rect 17570 2701 17604 2717
rect 17570 2683 17604 2701
rect 17570 2633 17604 2645
rect 17570 2611 17604 2633
rect 17570 2565 17604 2573
rect 17570 2539 17604 2565
rect 17666 3483 17700 3509
rect 17666 3475 17700 3483
rect 17666 3415 17700 3437
rect 17666 3403 17700 3415
rect 17666 3347 17700 3365
rect 17666 3331 17700 3347
rect 17666 3279 17700 3293
rect 17666 3259 17700 3279
rect 17666 3211 17700 3221
rect 17666 3187 17700 3211
rect 17666 3143 17700 3149
rect 17666 3115 17700 3143
rect 17666 3075 17700 3077
rect 17666 3043 17700 3075
rect 17666 2973 17700 3005
rect 17666 2971 17700 2973
rect 17666 2905 17700 2933
rect 17666 2899 17700 2905
rect 17666 2837 17700 2861
rect 17666 2827 17700 2837
rect 17666 2769 17700 2789
rect 17666 2755 17700 2769
rect 17666 2701 17700 2717
rect 17666 2683 17700 2701
rect 17666 2633 17700 2645
rect 17666 2611 17700 2633
rect 17666 2565 17700 2573
rect 17666 2539 17700 2565
rect 17762 3483 17796 3509
rect 17762 3475 17796 3483
rect 17762 3415 17796 3437
rect 17762 3403 17796 3415
rect 17762 3347 17796 3365
rect 17762 3331 17796 3347
rect 17762 3279 17796 3293
rect 17762 3259 17796 3279
rect 17762 3211 17796 3221
rect 17762 3187 17796 3211
rect 17762 3143 17796 3149
rect 17762 3115 17796 3143
rect 17762 3075 17796 3077
rect 17762 3043 17796 3075
rect 17762 2973 17796 3005
rect 17762 2971 17796 2973
rect 17762 2905 17796 2933
rect 17762 2899 17796 2905
rect 17762 2837 17796 2861
rect 17762 2827 17796 2837
rect 17762 2769 17796 2789
rect 17762 2755 17796 2769
rect 17762 2701 17796 2717
rect 17762 2683 17796 2701
rect 17762 2633 17796 2645
rect 17762 2611 17796 2633
rect 17762 2565 17796 2573
rect 17762 2539 17796 2565
rect 17858 3483 17892 3509
rect 17858 3475 17892 3483
rect 17858 3415 17892 3437
rect 17858 3403 17892 3415
rect 17858 3347 17892 3365
rect 17858 3331 17892 3347
rect 17858 3279 17892 3293
rect 17858 3259 17892 3279
rect 17858 3211 17892 3221
rect 17858 3187 17892 3211
rect 17858 3143 17892 3149
rect 17858 3115 17892 3143
rect 17858 3075 17892 3077
rect 17858 3043 17892 3075
rect 17858 2973 17892 3005
rect 17858 2971 17892 2973
rect 17858 2905 17892 2933
rect 17858 2899 17892 2905
rect 17858 2837 17892 2861
rect 17858 2827 17892 2837
rect 17858 2769 17892 2789
rect 17858 2755 17892 2769
rect 17858 2701 17892 2717
rect 17858 2683 17892 2701
rect 17858 2633 17892 2645
rect 17858 2611 17892 2633
rect 17858 2565 17892 2573
rect 17858 2539 17892 2565
rect 17954 3483 17988 3509
rect 17954 3475 17988 3483
rect 17954 3415 17988 3437
rect 17954 3403 17988 3415
rect 17954 3347 17988 3365
rect 17954 3331 17988 3347
rect 17954 3279 17988 3293
rect 17954 3259 17988 3279
rect 17954 3211 17988 3221
rect 17954 3187 17988 3211
rect 17954 3143 17988 3149
rect 17954 3115 17988 3143
rect 17954 3075 17988 3077
rect 17954 3043 17988 3075
rect 17954 2973 17988 3005
rect 17954 2971 17988 2973
rect 17954 2905 17988 2933
rect 17954 2899 17988 2905
rect 17954 2837 17988 2861
rect 17954 2827 17988 2837
rect 17954 2769 17988 2789
rect 17954 2755 17988 2769
rect 17954 2701 17988 2717
rect 17954 2683 17988 2701
rect 17954 2633 17988 2645
rect 17954 2611 17988 2633
rect 17954 2565 17988 2573
rect 17954 2539 17988 2565
rect 18050 3483 18084 3509
rect 18050 3475 18084 3483
rect 18050 3415 18084 3437
rect 18050 3403 18084 3415
rect 18050 3347 18084 3365
rect 18050 3331 18084 3347
rect 18050 3279 18084 3293
rect 18050 3259 18084 3279
rect 18050 3211 18084 3221
rect 18050 3187 18084 3211
rect 18050 3143 18084 3149
rect 18050 3115 18084 3143
rect 18050 3075 18084 3077
rect 18050 3043 18084 3075
rect 18050 2973 18084 3005
rect 18050 2971 18084 2973
rect 18050 2905 18084 2933
rect 18050 2899 18084 2905
rect 18050 2837 18084 2861
rect 18050 2827 18084 2837
rect 18050 2769 18084 2789
rect 18050 2755 18084 2769
rect 18050 2701 18084 2717
rect 18050 2683 18084 2701
rect 18050 2633 18084 2645
rect 18050 2611 18084 2633
rect 18050 2565 18084 2573
rect 18050 2539 18084 2565
rect 18146 3483 18180 3509
rect 18146 3475 18180 3483
rect 18146 3415 18180 3437
rect 18146 3403 18180 3415
rect 18146 3347 18180 3365
rect 18146 3331 18180 3347
rect 18146 3279 18180 3293
rect 18146 3259 18180 3279
rect 18146 3211 18180 3221
rect 18146 3187 18180 3211
rect 18146 3143 18180 3149
rect 18146 3115 18180 3143
rect 18146 3075 18180 3077
rect 18146 3043 18180 3075
rect 18146 2973 18180 3005
rect 18146 2971 18180 2973
rect 18146 2905 18180 2933
rect 18146 2899 18180 2905
rect 18146 2837 18180 2861
rect 18146 2827 18180 2837
rect 18146 2769 18180 2789
rect 18146 2755 18180 2769
rect 18146 2701 18180 2717
rect 18146 2683 18180 2701
rect 18146 2633 18180 2645
rect 18146 2611 18180 2633
rect 18146 2565 18180 2573
rect 18146 2539 18180 2565
rect 25354 5079 25388 5105
rect 25354 5071 25388 5079
rect 25354 5011 25388 5033
rect 25354 4999 25388 5011
rect 25354 4943 25388 4961
rect 25354 4927 25388 4943
rect 25354 4875 25388 4889
rect 25354 4855 25388 4875
rect 25354 4807 25388 4817
rect 25354 4783 25388 4807
rect 25354 4739 25388 4745
rect 25354 4711 25388 4739
rect 25354 4671 25388 4673
rect 25354 4639 25388 4671
rect 25354 4569 25388 4601
rect 25354 4567 25388 4569
rect 25354 4501 25388 4529
rect 25354 4495 25388 4501
rect 25354 4433 25388 4457
rect 25354 4423 25388 4433
rect 25354 4365 25388 4385
rect 25354 4351 25388 4365
rect 25354 4297 25388 4313
rect 25354 4279 25388 4297
rect 25354 4229 25388 4241
rect 25354 4207 25388 4229
rect 25354 4161 25388 4169
rect 25354 4135 25388 4161
rect 25450 5079 25484 5105
rect 25450 5071 25484 5079
rect 25450 5011 25484 5033
rect 25450 4999 25484 5011
rect 25450 4943 25484 4961
rect 25450 4927 25484 4943
rect 25450 4875 25484 4889
rect 25450 4855 25484 4875
rect 25450 4807 25484 4817
rect 25450 4783 25484 4807
rect 25450 4739 25484 4745
rect 25450 4711 25484 4739
rect 25450 4671 25484 4673
rect 25450 4639 25484 4671
rect 25450 4569 25484 4601
rect 25450 4567 25484 4569
rect 25450 4501 25484 4529
rect 25450 4495 25484 4501
rect 25450 4433 25484 4457
rect 25450 4423 25484 4433
rect 25450 4365 25484 4385
rect 25450 4351 25484 4365
rect 25450 4297 25484 4313
rect 25450 4279 25484 4297
rect 25450 4229 25484 4241
rect 25450 4207 25484 4229
rect 25450 4161 25484 4169
rect 25450 4135 25484 4161
rect 25546 5079 25580 5105
rect 25546 5071 25580 5079
rect 25546 5011 25580 5033
rect 25546 4999 25580 5011
rect 25546 4943 25580 4961
rect 25546 4927 25580 4943
rect 25546 4875 25580 4889
rect 25546 4855 25580 4875
rect 25546 4807 25580 4817
rect 25546 4783 25580 4807
rect 25546 4739 25580 4745
rect 25546 4711 25580 4739
rect 25546 4671 25580 4673
rect 25546 4639 25580 4671
rect 25546 4569 25580 4601
rect 25546 4567 25580 4569
rect 25546 4501 25580 4529
rect 25546 4495 25580 4501
rect 25546 4433 25580 4457
rect 25546 4423 25580 4433
rect 25546 4365 25580 4385
rect 25546 4351 25580 4365
rect 25546 4297 25580 4313
rect 25546 4279 25580 4297
rect 25546 4229 25580 4241
rect 25546 4207 25580 4229
rect 25546 4161 25580 4169
rect 25546 4135 25580 4161
rect 25642 5079 25676 5105
rect 25642 5071 25676 5079
rect 25642 5011 25676 5033
rect 25642 4999 25676 5011
rect 25642 4943 25676 4961
rect 25642 4927 25676 4943
rect 25642 4875 25676 4889
rect 25642 4855 25676 4875
rect 25642 4807 25676 4817
rect 25642 4783 25676 4807
rect 25642 4739 25676 4745
rect 25642 4711 25676 4739
rect 25642 4671 25676 4673
rect 25642 4639 25676 4671
rect 25642 4569 25676 4601
rect 25642 4567 25676 4569
rect 25642 4501 25676 4529
rect 25642 4495 25676 4501
rect 25642 4433 25676 4457
rect 25642 4423 25676 4433
rect 25642 4365 25676 4385
rect 25642 4351 25676 4365
rect 25642 4297 25676 4313
rect 25642 4279 25676 4297
rect 25642 4229 25676 4241
rect 25642 4207 25676 4229
rect 25642 4161 25676 4169
rect 25642 4135 25676 4161
rect 25738 5079 25772 5105
rect 25738 5071 25772 5079
rect 25738 5011 25772 5033
rect 25738 4999 25772 5011
rect 25738 4943 25772 4961
rect 25738 4927 25772 4943
rect 25738 4875 25772 4889
rect 25738 4855 25772 4875
rect 25738 4807 25772 4817
rect 25738 4783 25772 4807
rect 25738 4739 25772 4745
rect 25738 4711 25772 4739
rect 25738 4671 25772 4673
rect 25738 4639 25772 4671
rect 25738 4569 25772 4601
rect 25738 4567 25772 4569
rect 25738 4501 25772 4529
rect 25738 4495 25772 4501
rect 25738 4433 25772 4457
rect 25738 4423 25772 4433
rect 25738 4365 25772 4385
rect 25738 4351 25772 4365
rect 25738 4297 25772 4313
rect 25738 4279 25772 4297
rect 25738 4229 25772 4241
rect 25738 4207 25772 4229
rect 25738 4161 25772 4169
rect 25738 4135 25772 4161
rect 25834 5079 25868 5105
rect 25834 5071 25868 5079
rect 25834 5011 25868 5033
rect 25834 4999 25868 5011
rect 25834 4943 25868 4961
rect 25834 4927 25868 4943
rect 25834 4875 25868 4889
rect 25834 4855 25868 4875
rect 25834 4807 25868 4817
rect 25834 4783 25868 4807
rect 25834 4739 25868 4745
rect 25834 4711 25868 4739
rect 25834 4671 25868 4673
rect 25834 4639 25868 4671
rect 25834 4569 25868 4601
rect 25834 4567 25868 4569
rect 25834 4501 25868 4529
rect 25834 4495 25868 4501
rect 25834 4433 25868 4457
rect 25834 4423 25868 4433
rect 25834 4365 25868 4385
rect 25834 4351 25868 4365
rect 25834 4297 25868 4313
rect 25834 4279 25868 4297
rect 25834 4229 25868 4241
rect 25834 4207 25868 4229
rect 25834 4161 25868 4169
rect 25834 4135 25868 4161
rect 25930 5079 25964 5105
rect 25930 5071 25964 5079
rect 25930 5011 25964 5033
rect 25930 4999 25964 5011
rect 25930 4943 25964 4961
rect 25930 4927 25964 4943
rect 25930 4875 25964 4889
rect 25930 4855 25964 4875
rect 25930 4807 25964 4817
rect 25930 4783 25964 4807
rect 25930 4739 25964 4745
rect 25930 4711 25964 4739
rect 25930 4671 25964 4673
rect 25930 4639 25964 4671
rect 25930 4569 25964 4601
rect 25930 4567 25964 4569
rect 25930 4501 25964 4529
rect 25930 4495 25964 4501
rect 25930 4433 25964 4457
rect 25930 4423 25964 4433
rect 25930 4365 25964 4385
rect 25930 4351 25964 4365
rect 25930 4297 25964 4313
rect 25930 4279 25964 4297
rect 25930 4229 25964 4241
rect 25930 4207 25964 4229
rect 25930 4161 25964 4169
rect 25930 4135 25964 4161
rect 26026 5079 26060 5105
rect 26026 5071 26060 5079
rect 26026 5011 26060 5033
rect 26026 4999 26060 5011
rect 26026 4943 26060 4961
rect 26026 4927 26060 4943
rect 26026 4875 26060 4889
rect 26026 4855 26060 4875
rect 26026 4807 26060 4817
rect 26026 4783 26060 4807
rect 26026 4739 26060 4745
rect 26026 4711 26060 4739
rect 26026 4671 26060 4673
rect 26026 4639 26060 4671
rect 26026 4569 26060 4601
rect 26026 4567 26060 4569
rect 26026 4501 26060 4529
rect 26026 4495 26060 4501
rect 26026 4433 26060 4457
rect 26026 4423 26060 4433
rect 26026 4365 26060 4385
rect 26026 4351 26060 4365
rect 26026 4297 26060 4313
rect 26026 4279 26060 4297
rect 26026 4229 26060 4241
rect 26026 4207 26060 4229
rect 26026 4161 26060 4169
rect 26026 4135 26060 4161
rect 26122 5079 26156 5105
rect 26122 5071 26156 5079
rect 26122 5011 26156 5033
rect 26122 4999 26156 5011
rect 26122 4943 26156 4961
rect 26122 4927 26156 4943
rect 26122 4875 26156 4889
rect 26122 4855 26156 4875
rect 26122 4807 26156 4817
rect 26122 4783 26156 4807
rect 26122 4739 26156 4745
rect 26122 4711 26156 4739
rect 26122 4671 26156 4673
rect 26122 4639 26156 4671
rect 26122 4569 26156 4601
rect 26122 4567 26156 4569
rect 26122 4501 26156 4529
rect 26122 4495 26156 4501
rect 26122 4433 26156 4457
rect 26122 4423 26156 4433
rect 26122 4365 26156 4385
rect 26122 4351 26156 4365
rect 26122 4297 26156 4313
rect 26122 4279 26156 4297
rect 26122 4229 26156 4241
rect 26122 4207 26156 4229
rect 26122 4161 26156 4169
rect 26122 4135 26156 4161
rect 26218 5079 26252 5105
rect 26218 5071 26252 5079
rect 26218 5011 26252 5033
rect 26218 4999 26252 5011
rect 26218 4943 26252 4961
rect 26218 4927 26252 4943
rect 26218 4875 26252 4889
rect 26218 4855 26252 4875
rect 26218 4807 26252 4817
rect 26218 4783 26252 4807
rect 26218 4739 26252 4745
rect 26218 4711 26252 4739
rect 26218 4671 26252 4673
rect 26218 4639 26252 4671
rect 26218 4569 26252 4601
rect 26218 4567 26252 4569
rect 26218 4501 26252 4529
rect 26218 4495 26252 4501
rect 26218 4433 26252 4457
rect 26218 4423 26252 4433
rect 26218 4365 26252 4385
rect 26218 4351 26252 4365
rect 26218 4297 26252 4313
rect 26218 4279 26252 4297
rect 26218 4229 26252 4241
rect 26218 4207 26252 4229
rect 26218 4161 26252 4169
rect 26218 4135 26252 4161
rect 26314 5079 26348 5105
rect 26314 5071 26348 5079
rect 26314 5011 26348 5033
rect 26314 4999 26348 5011
rect 26314 4943 26348 4961
rect 26314 4927 26348 4943
rect 26314 4875 26348 4889
rect 26314 4855 26348 4875
rect 26314 4807 26348 4817
rect 26314 4783 26348 4807
rect 26314 4739 26348 4745
rect 26314 4711 26348 4739
rect 26314 4671 26348 4673
rect 26314 4639 26348 4671
rect 26314 4569 26348 4601
rect 26314 4567 26348 4569
rect 26314 4501 26348 4529
rect 26314 4495 26348 4501
rect 26314 4433 26348 4457
rect 26314 4423 26348 4433
rect 26314 4365 26348 4385
rect 26314 4351 26348 4365
rect 26314 4297 26348 4313
rect 26314 4279 26348 4297
rect 26314 4229 26348 4241
rect 26314 4207 26348 4229
rect 26314 4161 26348 4169
rect 26314 4135 26348 4161
rect 26410 5079 26444 5105
rect 26410 5071 26444 5079
rect 26410 5011 26444 5033
rect 26410 4999 26444 5011
rect 26410 4943 26444 4961
rect 26410 4927 26444 4943
rect 26410 4875 26444 4889
rect 26410 4855 26444 4875
rect 26410 4807 26444 4817
rect 26410 4783 26444 4807
rect 26410 4739 26444 4745
rect 26410 4711 26444 4739
rect 26410 4671 26444 4673
rect 26410 4639 26444 4671
rect 26410 4569 26444 4601
rect 26410 4567 26444 4569
rect 26410 4501 26444 4529
rect 26410 4495 26444 4501
rect 26410 4433 26444 4457
rect 26410 4423 26444 4433
rect 26410 4365 26444 4385
rect 26410 4351 26444 4365
rect 26410 4297 26444 4313
rect 26410 4279 26444 4297
rect 26410 4229 26444 4241
rect 26410 4207 26444 4229
rect 26410 4161 26444 4169
rect 26410 4135 26444 4161
rect 26506 5079 26540 5105
rect 26506 5071 26540 5079
rect 26506 5011 26540 5033
rect 26506 4999 26540 5011
rect 26506 4943 26540 4961
rect 26506 4927 26540 4943
rect 26506 4875 26540 4889
rect 26506 4855 26540 4875
rect 26506 4807 26540 4817
rect 26506 4783 26540 4807
rect 26506 4739 26540 4745
rect 26506 4711 26540 4739
rect 26506 4671 26540 4673
rect 26506 4639 26540 4671
rect 26506 4569 26540 4601
rect 26506 4567 26540 4569
rect 26506 4501 26540 4529
rect 26506 4495 26540 4501
rect 26506 4433 26540 4457
rect 26506 4423 26540 4433
rect 26506 4365 26540 4385
rect 26506 4351 26540 4365
rect 26506 4297 26540 4313
rect 26506 4279 26540 4297
rect 26506 4229 26540 4241
rect 26506 4207 26540 4229
rect 26506 4161 26540 4169
rect 26506 4135 26540 4161
rect 26602 5079 26636 5105
rect 26602 5071 26636 5079
rect 26602 5011 26636 5033
rect 26602 4999 26636 5011
rect 26602 4943 26636 4961
rect 26602 4927 26636 4943
rect 26602 4875 26636 4889
rect 26602 4855 26636 4875
rect 26602 4807 26636 4817
rect 26602 4783 26636 4807
rect 26602 4739 26636 4745
rect 26602 4711 26636 4739
rect 26602 4671 26636 4673
rect 26602 4639 26636 4671
rect 26602 4569 26636 4601
rect 26602 4567 26636 4569
rect 26602 4501 26636 4529
rect 26602 4495 26636 4501
rect 26602 4433 26636 4457
rect 26602 4423 26636 4433
rect 26602 4365 26636 4385
rect 26602 4351 26636 4365
rect 26602 4297 26636 4313
rect 26602 4279 26636 4297
rect 26602 4229 26636 4241
rect 26602 4207 26636 4229
rect 26602 4161 26636 4169
rect 26602 4135 26636 4161
rect 26826 5073 26860 5099
rect 26826 5065 26860 5073
rect 26826 5005 26860 5027
rect 26826 4993 26860 5005
rect 26826 4937 26860 4955
rect 26826 4921 26860 4937
rect 26826 4869 26860 4883
rect 26826 4849 26860 4869
rect 26826 4801 26860 4811
rect 26826 4777 26860 4801
rect 26826 4733 26860 4739
rect 26826 4705 26860 4733
rect 26826 4665 26860 4667
rect 26826 4633 26860 4665
rect 26826 4563 26860 4595
rect 26826 4561 26860 4563
rect 26826 4495 26860 4523
rect 26826 4489 26860 4495
rect 26826 4427 26860 4451
rect 26826 4417 26860 4427
rect 26826 4359 26860 4379
rect 26826 4345 26860 4359
rect 26826 4291 26860 4307
rect 26826 4273 26860 4291
rect 26826 4223 26860 4235
rect 26826 4201 26860 4223
rect 26826 4155 26860 4163
rect 26826 4129 26860 4155
rect 26922 5073 26956 5099
rect 26922 5065 26956 5073
rect 26922 5005 26956 5027
rect 26922 4993 26956 5005
rect 26922 4937 26956 4955
rect 26922 4921 26956 4937
rect 26922 4869 26956 4883
rect 26922 4849 26956 4869
rect 26922 4801 26956 4811
rect 26922 4777 26956 4801
rect 26922 4733 26956 4739
rect 26922 4705 26956 4733
rect 26922 4665 26956 4667
rect 26922 4633 26956 4665
rect 26922 4563 26956 4595
rect 26922 4561 26956 4563
rect 26922 4495 26956 4523
rect 26922 4489 26956 4495
rect 26922 4427 26956 4451
rect 26922 4417 26956 4427
rect 26922 4359 26956 4379
rect 26922 4345 26956 4359
rect 26922 4291 26956 4307
rect 26922 4273 26956 4291
rect 26922 4223 26956 4235
rect 26922 4201 26956 4223
rect 26922 4155 26956 4163
rect 26922 4129 26956 4155
rect 24006 3925 24040 3959
rect 23462 3785 23496 3819
rect 23318 3670 23352 3704
rect 27018 5073 27052 5099
rect 27018 5065 27052 5073
rect 27018 5005 27052 5027
rect 27018 4993 27052 5005
rect 27018 4937 27052 4955
rect 27018 4921 27052 4937
rect 27018 4869 27052 4883
rect 27018 4849 27052 4869
rect 27018 4801 27052 4811
rect 27018 4777 27052 4801
rect 27018 4733 27052 4739
rect 27018 4705 27052 4733
rect 27018 4665 27052 4667
rect 27018 4633 27052 4665
rect 27018 4563 27052 4595
rect 27018 4561 27052 4563
rect 27018 4495 27052 4523
rect 27018 4489 27052 4495
rect 27018 4427 27052 4451
rect 27018 4417 27052 4427
rect 27018 4359 27052 4379
rect 27018 4345 27052 4359
rect 27018 4291 27052 4307
rect 27018 4273 27052 4291
rect 27018 4223 27052 4235
rect 27018 4201 27052 4223
rect 27018 4155 27052 4163
rect 27018 4129 27052 4155
rect 27114 5073 27148 5099
rect 27114 5065 27148 5073
rect 27114 5005 27148 5027
rect 27114 4993 27148 5005
rect 27114 4937 27148 4955
rect 27114 4921 27148 4937
rect 27114 4869 27148 4883
rect 27114 4849 27148 4869
rect 27114 4801 27148 4811
rect 27114 4777 27148 4801
rect 27114 4733 27148 4739
rect 27114 4705 27148 4733
rect 27114 4665 27148 4667
rect 27114 4633 27148 4665
rect 27114 4563 27148 4595
rect 27114 4561 27148 4563
rect 27114 4495 27148 4523
rect 27114 4489 27148 4495
rect 27114 4427 27148 4451
rect 27114 4417 27148 4427
rect 27114 4359 27148 4379
rect 27114 4345 27148 4359
rect 27114 4291 27148 4307
rect 27114 4273 27148 4291
rect 27114 4223 27148 4235
rect 27114 4201 27148 4223
rect 27114 4155 27148 4163
rect 27114 4129 27148 4155
rect 27210 5073 27244 5099
rect 27210 5065 27244 5073
rect 27210 5005 27244 5027
rect 27210 4993 27244 5005
rect 27210 4937 27244 4955
rect 27210 4921 27244 4937
rect 27210 4869 27244 4883
rect 27210 4849 27244 4869
rect 27210 4801 27244 4811
rect 27210 4777 27244 4801
rect 27210 4733 27244 4739
rect 27210 4705 27244 4733
rect 27210 4665 27244 4667
rect 27210 4633 27244 4665
rect 27210 4563 27244 4595
rect 27210 4561 27244 4563
rect 27210 4495 27244 4523
rect 27210 4489 27244 4495
rect 27210 4427 27244 4451
rect 27210 4417 27244 4427
rect 27210 4359 27244 4379
rect 27210 4345 27244 4359
rect 27210 4291 27244 4307
rect 27210 4273 27244 4291
rect 27210 4223 27244 4235
rect 27210 4201 27244 4223
rect 27210 4155 27244 4163
rect 27210 4129 27244 4155
rect 27306 5073 27340 5099
rect 27306 5065 27340 5073
rect 27306 5005 27340 5027
rect 27306 4993 27340 5005
rect 27306 4937 27340 4955
rect 27306 4921 27340 4937
rect 27306 4869 27340 4883
rect 27306 4849 27340 4869
rect 27306 4801 27340 4811
rect 27306 4777 27340 4801
rect 27306 4733 27340 4739
rect 27306 4705 27340 4733
rect 27306 4665 27340 4667
rect 27306 4633 27340 4665
rect 27306 4563 27340 4595
rect 27306 4561 27340 4563
rect 27306 4495 27340 4523
rect 27306 4489 27340 4495
rect 27306 4427 27340 4451
rect 27306 4417 27340 4427
rect 27306 4359 27340 4379
rect 27306 4345 27340 4359
rect 27306 4291 27340 4307
rect 27306 4273 27340 4291
rect 27306 4223 27340 4235
rect 27306 4201 27340 4223
rect 27306 4155 27340 4163
rect 27306 4129 27340 4155
rect 27402 5073 27436 5099
rect 27402 5065 27436 5073
rect 27402 5005 27436 5027
rect 27402 4993 27436 5005
rect 27402 4937 27436 4955
rect 27402 4921 27436 4937
rect 27402 4869 27436 4883
rect 27402 4849 27436 4869
rect 27402 4801 27436 4811
rect 27402 4777 27436 4801
rect 27402 4733 27436 4739
rect 27402 4705 27436 4733
rect 27402 4665 27436 4667
rect 27402 4633 27436 4665
rect 27402 4563 27436 4595
rect 27402 4561 27436 4563
rect 27402 4495 27436 4523
rect 27402 4489 27436 4495
rect 27402 4427 27436 4451
rect 27402 4417 27436 4427
rect 27402 4359 27436 4379
rect 27402 4345 27436 4359
rect 27402 4291 27436 4307
rect 27402 4273 27436 4291
rect 27402 4223 27436 4235
rect 27402 4201 27436 4223
rect 27402 4155 27436 4163
rect 27402 4129 27436 4155
rect 27498 5073 27532 5099
rect 27498 5065 27532 5073
rect 27498 5005 27532 5027
rect 27498 4993 27532 5005
rect 27498 4937 27532 4955
rect 27498 4921 27532 4937
rect 27498 4869 27532 4883
rect 27498 4849 27532 4869
rect 27498 4801 27532 4811
rect 27498 4777 27532 4801
rect 27498 4733 27532 4739
rect 27498 4705 27532 4733
rect 27498 4665 27532 4667
rect 27498 4633 27532 4665
rect 27498 4563 27532 4595
rect 27498 4561 27532 4563
rect 27498 4495 27532 4523
rect 27498 4489 27532 4495
rect 27498 4427 27532 4451
rect 27498 4417 27532 4427
rect 27498 4359 27532 4379
rect 27498 4345 27532 4359
rect 27498 4291 27532 4307
rect 27498 4273 27532 4291
rect 27498 4223 27532 4235
rect 27498 4201 27532 4223
rect 27498 4155 27532 4163
rect 27498 4129 27532 4155
rect 27594 5073 27628 5099
rect 27594 5065 27628 5073
rect 27594 5005 27628 5027
rect 27594 4993 27628 5005
rect 27594 4937 27628 4955
rect 27594 4921 27628 4937
rect 27594 4869 27628 4883
rect 27594 4849 27628 4869
rect 27594 4801 27628 4811
rect 27594 4777 27628 4801
rect 27594 4733 27628 4739
rect 27594 4705 27628 4733
rect 27594 4665 27628 4667
rect 27594 4633 27628 4665
rect 27594 4563 27628 4595
rect 27594 4561 27628 4563
rect 27594 4495 27628 4523
rect 27594 4489 27628 4495
rect 27594 4427 27628 4451
rect 27594 4417 27628 4427
rect 27594 4359 27628 4379
rect 27594 4345 27628 4359
rect 27594 4291 27628 4307
rect 27594 4273 27628 4291
rect 27594 4223 27628 4235
rect 27594 4201 27628 4223
rect 27594 4155 27628 4163
rect 27594 4129 27628 4155
rect 27690 5073 27724 5099
rect 27690 5065 27724 5073
rect 27690 5005 27724 5027
rect 27690 4993 27724 5005
rect 27690 4937 27724 4955
rect 27690 4921 27724 4937
rect 27690 4869 27724 4883
rect 27690 4849 27724 4869
rect 27690 4801 27724 4811
rect 27690 4777 27724 4801
rect 27690 4733 27724 4739
rect 27690 4705 27724 4733
rect 27690 4665 27724 4667
rect 27690 4633 27724 4665
rect 27690 4563 27724 4595
rect 27690 4561 27724 4563
rect 27690 4495 27724 4523
rect 27690 4489 27724 4495
rect 27690 4427 27724 4451
rect 27690 4417 27724 4427
rect 27690 4359 27724 4379
rect 27690 4345 27724 4359
rect 27690 4291 27724 4307
rect 27690 4273 27724 4291
rect 27690 4223 27724 4235
rect 27690 4201 27724 4223
rect 27690 4155 27724 4163
rect 27690 4129 27724 4155
rect 27786 5073 27820 5099
rect 27786 5065 27820 5073
rect 27786 5005 27820 5027
rect 27786 4993 27820 5005
rect 27786 4937 27820 4955
rect 27786 4921 27820 4937
rect 27786 4869 27820 4883
rect 27786 4849 27820 4869
rect 27786 4801 27820 4811
rect 27786 4777 27820 4801
rect 27786 4733 27820 4739
rect 27786 4705 27820 4733
rect 27786 4665 27820 4667
rect 27786 4633 27820 4665
rect 27786 4563 27820 4595
rect 27786 4561 27820 4563
rect 27786 4495 27820 4523
rect 27786 4489 27820 4495
rect 27786 4427 27820 4451
rect 27786 4417 27820 4427
rect 27786 4359 27820 4379
rect 27786 4345 27820 4359
rect 27786 4291 27820 4307
rect 27786 4273 27820 4291
rect 27786 4223 27820 4235
rect 27786 4201 27820 4223
rect 27786 4155 27820 4163
rect 27786 4129 27820 4155
rect 27882 5073 27916 5099
rect 27882 5065 27916 5073
rect 27882 5005 27916 5027
rect 27882 4993 27916 5005
rect 27882 4937 27916 4955
rect 27882 4921 27916 4937
rect 27882 4869 27916 4883
rect 27882 4849 27916 4869
rect 27882 4801 27916 4811
rect 27882 4777 27916 4801
rect 27882 4733 27916 4739
rect 27882 4705 27916 4733
rect 27882 4665 27916 4667
rect 27882 4633 27916 4665
rect 27882 4563 27916 4595
rect 27882 4561 27916 4563
rect 27882 4495 27916 4523
rect 27882 4489 27916 4495
rect 27882 4427 27916 4451
rect 27882 4417 27916 4427
rect 27882 4359 27916 4379
rect 27882 4345 27916 4359
rect 27882 4291 27916 4307
rect 27882 4273 27916 4291
rect 27882 4223 27916 4235
rect 27882 4201 27916 4223
rect 27882 4155 27916 4163
rect 27882 4129 27916 4155
rect 27978 5073 28012 5099
rect 27978 5065 28012 5073
rect 27978 5005 28012 5027
rect 27978 4993 28012 5005
rect 27978 4937 28012 4955
rect 27978 4921 28012 4937
rect 27978 4869 28012 4883
rect 27978 4849 28012 4869
rect 27978 4801 28012 4811
rect 27978 4777 28012 4801
rect 27978 4733 28012 4739
rect 27978 4705 28012 4733
rect 27978 4665 28012 4667
rect 27978 4633 28012 4665
rect 27978 4563 28012 4595
rect 27978 4561 28012 4563
rect 27978 4495 28012 4523
rect 27978 4489 28012 4495
rect 27978 4427 28012 4451
rect 27978 4417 28012 4427
rect 27978 4359 28012 4379
rect 27978 4345 28012 4359
rect 27978 4291 28012 4307
rect 27978 4273 28012 4291
rect 27978 4223 28012 4235
rect 27978 4201 28012 4223
rect 27978 4155 28012 4163
rect 27978 4129 28012 4155
rect 28074 5073 28108 5099
rect 28074 5065 28108 5073
rect 28074 5005 28108 5027
rect 28074 4993 28108 5005
rect 28074 4937 28108 4955
rect 28074 4921 28108 4937
rect 28074 4869 28108 4883
rect 28074 4849 28108 4869
rect 28074 4801 28108 4811
rect 28074 4777 28108 4801
rect 28074 4733 28108 4739
rect 28074 4705 28108 4733
rect 28074 4665 28108 4667
rect 28074 4633 28108 4665
rect 28074 4563 28108 4595
rect 28074 4561 28108 4563
rect 28074 4495 28108 4523
rect 28074 4489 28108 4495
rect 28074 4427 28108 4451
rect 28074 4417 28108 4427
rect 28074 4359 28108 4379
rect 28074 4345 28108 4359
rect 28074 4291 28108 4307
rect 28074 4273 28108 4291
rect 28074 4223 28108 4235
rect 28074 4201 28108 4223
rect 28074 4155 28108 4163
rect 28074 4129 28108 4155
rect 28170 5073 28204 5099
rect 28170 5065 28204 5073
rect 28170 5005 28204 5027
rect 28170 4993 28204 5005
rect 28170 4937 28204 4955
rect 28170 4921 28204 4937
rect 28170 4869 28204 4883
rect 28170 4849 28204 4869
rect 28170 4801 28204 4811
rect 28170 4777 28204 4801
rect 28170 4733 28204 4739
rect 28170 4705 28204 4733
rect 28170 4665 28204 4667
rect 28170 4633 28204 4665
rect 28170 4563 28204 4595
rect 28170 4561 28204 4563
rect 28170 4495 28204 4523
rect 28170 4489 28204 4495
rect 28170 4427 28204 4451
rect 28170 4417 28204 4427
rect 28170 4359 28204 4379
rect 28170 4345 28204 4359
rect 28170 4291 28204 4307
rect 28170 4273 28204 4291
rect 28170 4223 28204 4235
rect 28170 4201 28204 4223
rect 28170 4155 28204 4163
rect 28170 4129 28204 4155
rect 28266 5073 28300 5099
rect 28266 5065 28300 5073
rect 28266 5005 28300 5027
rect 28266 4993 28300 5005
rect 28266 4937 28300 4955
rect 28266 4921 28300 4937
rect 28266 4869 28300 4883
rect 28266 4849 28300 4869
rect 28266 4801 28300 4811
rect 28266 4777 28300 4801
rect 28266 4733 28300 4739
rect 28266 4705 28300 4733
rect 28266 4665 28300 4667
rect 28266 4633 28300 4665
rect 28266 4563 28300 4595
rect 28266 4561 28300 4563
rect 28266 4495 28300 4523
rect 28266 4489 28300 4495
rect 28266 4427 28300 4451
rect 28266 4417 28300 4427
rect 28266 4359 28300 4379
rect 28266 4345 28300 4359
rect 28266 4291 28300 4307
rect 28266 4273 28300 4291
rect 28266 4223 28300 4235
rect 28266 4201 28300 4223
rect 28266 4155 28300 4163
rect 28266 4129 28300 4155
rect 28362 5073 28396 5099
rect 28362 5065 28396 5073
rect 28362 5005 28396 5027
rect 28362 4993 28396 5005
rect 28362 4937 28396 4955
rect 28362 4921 28396 4937
rect 28362 4869 28396 4883
rect 28362 4849 28396 4869
rect 28362 4801 28396 4811
rect 28362 4777 28396 4801
rect 28362 4733 28396 4739
rect 28362 4705 28396 4733
rect 28362 4665 28396 4667
rect 28362 4633 28396 4665
rect 28362 4563 28396 4595
rect 28362 4561 28396 4563
rect 28362 4495 28396 4523
rect 28362 4489 28396 4495
rect 28362 4427 28396 4451
rect 28362 4417 28396 4427
rect 28362 4359 28396 4379
rect 28362 4345 28396 4359
rect 28362 4291 28396 4307
rect 28362 4273 28396 4291
rect 28362 4223 28396 4235
rect 28362 4201 28396 4223
rect 28362 4155 28396 4163
rect 28362 4129 28396 4155
rect 28458 5073 28492 5099
rect 28458 5065 28492 5073
rect 28458 5005 28492 5027
rect 28458 4993 28492 5005
rect 28458 4937 28492 4955
rect 28458 4921 28492 4937
rect 28458 4869 28492 4883
rect 28458 4849 28492 4869
rect 28458 4801 28492 4811
rect 28458 4777 28492 4801
rect 28458 4733 28492 4739
rect 28458 4705 28492 4733
rect 28458 4665 28492 4667
rect 28458 4633 28492 4665
rect 28458 4563 28492 4595
rect 28458 4561 28492 4563
rect 28458 4495 28492 4523
rect 28458 4489 28492 4495
rect 28458 4427 28492 4451
rect 28458 4417 28492 4427
rect 28458 4359 28492 4379
rect 28458 4345 28492 4359
rect 28458 4291 28492 4307
rect 28458 4273 28492 4291
rect 28458 4223 28492 4235
rect 28458 4201 28492 4223
rect 28458 4155 28492 4163
rect 28458 4129 28492 4155
rect 28554 5073 28588 5099
rect 28554 5065 28588 5073
rect 28554 5005 28588 5027
rect 28554 4993 28588 5005
rect 28554 4937 28588 4955
rect 28554 4921 28588 4937
rect 28554 4869 28588 4883
rect 28554 4849 28588 4869
rect 28554 4801 28588 4811
rect 28554 4777 28588 4801
rect 28554 4733 28588 4739
rect 28554 4705 28588 4733
rect 28554 4665 28588 4667
rect 28554 4633 28588 4665
rect 28554 4563 28588 4595
rect 28554 4561 28588 4563
rect 28554 4495 28588 4523
rect 28554 4489 28588 4495
rect 28554 4427 28588 4451
rect 28554 4417 28588 4427
rect 28554 4359 28588 4379
rect 28554 4345 28588 4359
rect 28554 4291 28588 4307
rect 28554 4273 28588 4291
rect 28554 4223 28588 4235
rect 28554 4201 28588 4223
rect 28554 4155 28588 4163
rect 28554 4129 28588 4155
rect 28650 5073 28684 5099
rect 28650 5065 28684 5073
rect 28650 5005 28684 5027
rect 28650 4993 28684 5005
rect 28650 4937 28684 4955
rect 28650 4921 28684 4937
rect 28650 4869 28684 4883
rect 28650 4849 28684 4869
rect 28650 4801 28684 4811
rect 28650 4777 28684 4801
rect 28650 4733 28684 4739
rect 28650 4705 28684 4733
rect 28650 4665 28684 4667
rect 28650 4633 28684 4665
rect 28650 4563 28684 4595
rect 28650 4561 28684 4563
rect 28650 4495 28684 4523
rect 28650 4489 28684 4495
rect 28650 4427 28684 4451
rect 28650 4417 28684 4427
rect 28650 4359 28684 4379
rect 28650 4345 28684 4359
rect 28650 4291 28684 4307
rect 28650 4273 28684 4291
rect 28650 4223 28684 4235
rect 28650 4201 28684 4223
rect 28650 4155 28684 4163
rect 28650 4129 28684 4155
rect 28746 5073 28780 5099
rect 28746 5065 28780 5073
rect 28746 5005 28780 5027
rect 28746 4993 28780 5005
rect 28746 4937 28780 4955
rect 28746 4921 28780 4937
rect 28746 4869 28780 4883
rect 28746 4849 28780 4869
rect 28746 4801 28780 4811
rect 28746 4777 28780 4801
rect 28746 4733 28780 4739
rect 28746 4705 28780 4733
rect 28746 4665 28780 4667
rect 28746 4633 28780 4665
rect 28746 4563 28780 4595
rect 28746 4561 28780 4563
rect 28746 4495 28780 4523
rect 28746 4489 28780 4495
rect 28746 4427 28780 4451
rect 28746 4417 28780 4427
rect 28746 4359 28780 4379
rect 28746 4345 28780 4359
rect 28746 4291 28780 4307
rect 28746 4273 28780 4291
rect 28746 4223 28780 4235
rect 28746 4201 28780 4223
rect 28746 4155 28780 4163
rect 28746 4129 28780 4155
rect 25210 3919 25244 3953
rect 24278 3783 24312 3817
rect 24010 3700 24044 3734
rect 26874 3913 26908 3947
rect 25931 3770 25965 3804
rect 25208 3656 25242 3690
rect 18242 3483 18276 3509
rect 18242 3475 18276 3483
rect 18242 3415 18276 3437
rect 18242 3403 18276 3415
rect 18242 3347 18276 3365
rect 18242 3331 18276 3347
rect 18242 3279 18276 3293
rect 18242 3259 18276 3279
rect 18242 3211 18276 3221
rect 18242 3187 18276 3211
rect 18242 3143 18276 3149
rect 18242 3115 18276 3143
rect 18242 3075 18276 3077
rect 18242 3043 18276 3075
rect 18242 2973 18276 3005
rect 18242 2971 18276 2973
rect 18242 2905 18276 2933
rect 18242 2899 18276 2905
rect 18242 2837 18276 2861
rect 18242 2827 18276 2837
rect 18242 2769 18276 2789
rect 18242 2755 18276 2769
rect 18242 2701 18276 2717
rect 18242 2683 18276 2701
rect 18242 2633 18276 2645
rect 18242 2611 18276 2633
rect 18242 2565 18276 2573
rect 18242 2539 18276 2565
rect 18338 3483 18372 3509
rect 18338 3475 18372 3483
rect 18338 3415 18372 3437
rect 18338 3403 18372 3415
rect 18338 3347 18372 3365
rect 18338 3331 18372 3347
rect 18338 3279 18372 3293
rect 18338 3259 18372 3279
rect 18338 3211 18372 3221
rect 18338 3187 18372 3211
rect 18338 3143 18372 3149
rect 18338 3115 18372 3143
rect 18338 3075 18372 3077
rect 18338 3043 18372 3075
rect 18338 2973 18372 3005
rect 18338 2971 18372 2973
rect 18338 2905 18372 2933
rect 18338 2899 18372 2905
rect 18338 2837 18372 2861
rect 18338 2827 18372 2837
rect 18338 2769 18372 2789
rect 18338 2755 18372 2769
rect 18338 2701 18372 2717
rect 18338 2683 18372 2701
rect 18338 2633 18372 2645
rect 18338 2611 18372 2633
rect 18338 2565 18372 2573
rect 18338 2539 18372 2565
rect 18576 3479 18610 3505
rect 18576 3471 18610 3479
rect 18576 3411 18610 3433
rect 18576 3399 18610 3411
rect 18576 3343 18610 3361
rect 18576 3327 18610 3343
rect 18576 3275 18610 3289
rect 18576 3255 18610 3275
rect 18576 3207 18610 3217
rect 18576 3183 18610 3207
rect 18576 3139 18610 3145
rect 18576 3111 18610 3139
rect 18576 3071 18610 3073
rect 18576 3039 18610 3071
rect 18576 2969 18610 3001
rect 18576 2967 18610 2969
rect 18576 2901 18610 2929
rect 18576 2895 18610 2901
rect 18576 2833 18610 2857
rect 18576 2823 18610 2833
rect 18576 2765 18610 2785
rect 18576 2751 18610 2765
rect 18576 2697 18610 2713
rect 18576 2679 18610 2697
rect 18576 2629 18610 2641
rect 18576 2607 18610 2629
rect 18576 2561 18610 2569
rect 18576 2535 18610 2561
rect 18672 3479 18706 3505
rect 18672 3471 18706 3479
rect 18672 3411 18706 3433
rect 18672 3399 18706 3411
rect 18672 3343 18706 3361
rect 18672 3327 18706 3343
rect 18672 3275 18706 3289
rect 18672 3255 18706 3275
rect 18672 3207 18706 3217
rect 18672 3183 18706 3207
rect 18672 3139 18706 3145
rect 18672 3111 18706 3139
rect 18672 3071 18706 3073
rect 18672 3039 18706 3071
rect 18672 2969 18706 3001
rect 18672 2967 18706 2969
rect 18672 2901 18706 2929
rect 18672 2895 18706 2901
rect 18672 2833 18706 2857
rect 18672 2823 18706 2833
rect 18672 2765 18706 2785
rect 18672 2751 18706 2765
rect 18672 2697 18706 2713
rect 18672 2679 18706 2697
rect 18672 2629 18706 2641
rect 18672 2607 18706 2629
rect 18672 2561 18706 2569
rect 18672 2535 18706 2561
rect 18768 3479 18802 3505
rect 18768 3471 18802 3479
rect 18768 3411 18802 3433
rect 18768 3399 18802 3411
rect 18768 3343 18802 3361
rect 18768 3327 18802 3343
rect 18768 3275 18802 3289
rect 18768 3255 18802 3275
rect 18768 3207 18802 3217
rect 18768 3183 18802 3207
rect 18768 3139 18802 3145
rect 18768 3111 18802 3139
rect 18768 3071 18802 3073
rect 18768 3039 18802 3071
rect 18768 2969 18802 3001
rect 18768 2967 18802 2969
rect 18768 2901 18802 2929
rect 18768 2895 18802 2901
rect 18768 2833 18802 2857
rect 18768 2823 18802 2833
rect 18768 2765 18802 2785
rect 18768 2751 18802 2765
rect 18768 2697 18802 2713
rect 18768 2679 18802 2697
rect 18768 2629 18802 2641
rect 18768 2607 18802 2629
rect 18768 2561 18802 2569
rect 18768 2535 18802 2561
rect 18864 3479 18898 3505
rect 18864 3471 18898 3479
rect 18864 3411 18898 3433
rect 18864 3399 18898 3411
rect 18864 3343 18898 3361
rect 18864 3327 18898 3343
rect 18864 3275 18898 3289
rect 18864 3255 18898 3275
rect 18864 3207 18898 3217
rect 18864 3183 18898 3207
rect 18864 3139 18898 3145
rect 18864 3111 18898 3139
rect 18864 3071 18898 3073
rect 18864 3039 18898 3071
rect 18864 2969 18898 3001
rect 18864 2967 18898 2969
rect 18864 2901 18898 2929
rect 18864 2895 18898 2901
rect 18864 2833 18898 2857
rect 18864 2823 18898 2833
rect 18864 2765 18898 2785
rect 18864 2751 18898 2765
rect 18864 2697 18898 2713
rect 18864 2679 18898 2697
rect 18864 2629 18898 2641
rect 18864 2607 18898 2629
rect 18864 2561 18898 2569
rect 18864 2535 18898 2561
rect 18960 3479 18994 3505
rect 18960 3471 18994 3479
rect 18960 3411 18994 3433
rect 18960 3399 18994 3411
rect 18960 3343 18994 3361
rect 18960 3327 18994 3343
rect 18960 3275 18994 3289
rect 18960 3255 18994 3275
rect 18960 3207 18994 3217
rect 18960 3183 18994 3207
rect 18960 3139 18994 3145
rect 18960 3111 18994 3139
rect 18960 3071 18994 3073
rect 18960 3039 18994 3071
rect 18960 2969 18994 3001
rect 18960 2967 18994 2969
rect 18960 2901 18994 2929
rect 18960 2895 18994 2901
rect 18960 2833 18994 2857
rect 18960 2823 18994 2833
rect 18960 2765 18994 2785
rect 18960 2751 18994 2765
rect 18960 2697 18994 2713
rect 18960 2679 18994 2697
rect 18960 2629 18994 2641
rect 18960 2607 18994 2629
rect 18960 2561 18994 2569
rect 18960 2535 18994 2561
rect 19056 3479 19090 3505
rect 19056 3471 19090 3479
rect 19056 3411 19090 3433
rect 19056 3399 19090 3411
rect 19056 3343 19090 3361
rect 19056 3327 19090 3343
rect 19056 3275 19090 3289
rect 19056 3255 19090 3275
rect 19056 3207 19090 3217
rect 19056 3183 19090 3207
rect 19056 3139 19090 3145
rect 19056 3111 19090 3139
rect 19056 3071 19090 3073
rect 19056 3039 19090 3071
rect 19056 2969 19090 3001
rect 19056 2967 19090 2969
rect 19056 2901 19090 2929
rect 19056 2895 19090 2901
rect 19056 2833 19090 2857
rect 19056 2823 19090 2833
rect 19056 2765 19090 2785
rect 19056 2751 19090 2765
rect 19056 2697 19090 2713
rect 19056 2679 19090 2697
rect 19056 2629 19090 2641
rect 19056 2607 19090 2629
rect 19056 2561 19090 2569
rect 19056 2535 19090 2561
rect 19152 3479 19186 3505
rect 19152 3471 19186 3479
rect 19152 3411 19186 3433
rect 19152 3399 19186 3411
rect 19152 3343 19186 3361
rect 19152 3327 19186 3343
rect 19152 3275 19186 3289
rect 19152 3255 19186 3275
rect 19152 3207 19186 3217
rect 19152 3183 19186 3207
rect 19152 3139 19186 3145
rect 19152 3111 19186 3139
rect 19152 3071 19186 3073
rect 19152 3039 19186 3071
rect 19152 2969 19186 3001
rect 19152 2967 19186 2969
rect 19152 2901 19186 2929
rect 19152 2895 19186 2901
rect 19152 2833 19186 2857
rect 19152 2823 19186 2833
rect 19152 2765 19186 2785
rect 19152 2751 19186 2765
rect 19152 2697 19186 2713
rect 19152 2679 19186 2697
rect 19152 2629 19186 2641
rect 19152 2607 19186 2629
rect 19152 2561 19186 2569
rect 19152 2535 19186 2561
rect 19248 3479 19282 3505
rect 19248 3471 19282 3479
rect 19248 3411 19282 3433
rect 19248 3399 19282 3411
rect 19248 3343 19282 3361
rect 19248 3327 19282 3343
rect 19248 3275 19282 3289
rect 19248 3255 19282 3275
rect 19248 3207 19282 3217
rect 19248 3183 19282 3207
rect 19248 3139 19282 3145
rect 19248 3111 19282 3139
rect 19248 3071 19282 3073
rect 19248 3039 19282 3071
rect 19248 2969 19282 3001
rect 19248 2967 19282 2969
rect 19248 2901 19282 2929
rect 19248 2895 19282 2901
rect 19248 2833 19282 2857
rect 19248 2823 19282 2833
rect 19248 2765 19282 2785
rect 19248 2751 19282 2765
rect 19248 2697 19282 2713
rect 19248 2679 19282 2697
rect 19248 2629 19282 2641
rect 19248 2607 19282 2629
rect 19248 2561 19282 2569
rect 19248 2535 19282 2561
rect 19344 3479 19378 3505
rect 19344 3471 19378 3479
rect 19344 3411 19378 3433
rect 19344 3399 19378 3411
rect 19344 3343 19378 3361
rect 19344 3327 19378 3343
rect 19344 3275 19378 3289
rect 19344 3255 19378 3275
rect 19344 3207 19378 3217
rect 19344 3183 19378 3207
rect 19344 3139 19378 3145
rect 19344 3111 19378 3139
rect 19344 3071 19378 3073
rect 19344 3039 19378 3071
rect 19344 2969 19378 3001
rect 19344 2967 19378 2969
rect 19344 2901 19378 2929
rect 19344 2895 19378 2901
rect 19344 2833 19378 2857
rect 19344 2823 19378 2833
rect 19344 2765 19378 2785
rect 19344 2751 19378 2765
rect 19344 2697 19378 2713
rect 19344 2679 19378 2697
rect 19344 2629 19378 2641
rect 19344 2607 19378 2629
rect 19344 2561 19378 2569
rect 19344 2535 19378 2561
rect 19440 3479 19474 3505
rect 19440 3471 19474 3479
rect 19440 3411 19474 3433
rect 19440 3399 19474 3411
rect 19440 3343 19474 3361
rect 19440 3327 19474 3343
rect 19440 3275 19474 3289
rect 19440 3255 19474 3275
rect 19440 3207 19474 3217
rect 19440 3183 19474 3207
rect 19440 3139 19474 3145
rect 19440 3111 19474 3139
rect 19440 3071 19474 3073
rect 19440 3039 19474 3071
rect 19440 2969 19474 3001
rect 19440 2967 19474 2969
rect 19440 2901 19474 2929
rect 19440 2895 19474 2901
rect 19440 2833 19474 2857
rect 19440 2823 19474 2833
rect 19440 2765 19474 2785
rect 19440 2751 19474 2765
rect 19440 2697 19474 2713
rect 19440 2679 19474 2697
rect 19440 2629 19474 2641
rect 19440 2607 19474 2629
rect 19440 2561 19474 2569
rect 19440 2535 19474 2561
rect 19536 3479 19570 3505
rect 19536 3471 19570 3479
rect 19536 3411 19570 3433
rect 19536 3399 19570 3411
rect 19536 3343 19570 3361
rect 19536 3327 19570 3343
rect 19536 3275 19570 3289
rect 19536 3255 19570 3275
rect 19536 3207 19570 3217
rect 19536 3183 19570 3207
rect 19536 3139 19570 3145
rect 19536 3111 19570 3139
rect 19536 3071 19570 3073
rect 19536 3039 19570 3071
rect 19536 2969 19570 3001
rect 19536 2967 19570 2969
rect 19536 2901 19570 2929
rect 19536 2895 19570 2901
rect 19536 2833 19570 2857
rect 19536 2823 19570 2833
rect 19536 2765 19570 2785
rect 19536 2751 19570 2765
rect 19536 2697 19570 2713
rect 19536 2679 19570 2697
rect 19536 2629 19570 2641
rect 19536 2607 19570 2629
rect 19536 2561 19570 2569
rect 19536 2535 19570 2561
rect 19632 3479 19666 3505
rect 19632 3471 19666 3479
rect 19632 3411 19666 3433
rect 19632 3399 19666 3411
rect 19632 3343 19666 3361
rect 19632 3327 19666 3343
rect 19632 3275 19666 3289
rect 19632 3255 19666 3275
rect 19632 3207 19666 3217
rect 19632 3183 19666 3207
rect 19632 3139 19666 3145
rect 19632 3111 19666 3139
rect 19632 3071 19666 3073
rect 19632 3039 19666 3071
rect 19632 2969 19666 3001
rect 19632 2967 19666 2969
rect 19632 2901 19666 2929
rect 19632 2895 19666 2901
rect 19632 2833 19666 2857
rect 19632 2823 19666 2833
rect 19632 2765 19666 2785
rect 19632 2751 19666 2765
rect 19632 2697 19666 2713
rect 19632 2679 19666 2697
rect 19632 2629 19666 2641
rect 19632 2607 19666 2629
rect 19632 2561 19666 2569
rect 19632 2535 19666 2561
rect 19728 3479 19762 3505
rect 19728 3471 19762 3479
rect 19728 3411 19762 3433
rect 19728 3399 19762 3411
rect 19728 3343 19762 3361
rect 19728 3327 19762 3343
rect 19728 3275 19762 3289
rect 19728 3255 19762 3275
rect 19728 3207 19762 3217
rect 19728 3183 19762 3207
rect 19728 3139 19762 3145
rect 19728 3111 19762 3139
rect 19728 3071 19762 3073
rect 19728 3039 19762 3071
rect 19728 2969 19762 3001
rect 19728 2967 19762 2969
rect 19728 2901 19762 2929
rect 19728 2895 19762 2901
rect 19728 2833 19762 2857
rect 19728 2823 19762 2833
rect 19728 2765 19762 2785
rect 19728 2751 19762 2765
rect 19728 2697 19762 2713
rect 19728 2679 19762 2697
rect 19728 2629 19762 2641
rect 19728 2607 19762 2629
rect 19728 2561 19762 2569
rect 19728 2535 19762 2561
rect 19824 3479 19858 3505
rect 19824 3471 19858 3479
rect 19824 3411 19858 3433
rect 19824 3399 19858 3411
rect 19824 3343 19858 3361
rect 19824 3327 19858 3343
rect 19824 3275 19858 3289
rect 19824 3255 19858 3275
rect 19824 3207 19858 3217
rect 19824 3183 19858 3207
rect 19824 3139 19858 3145
rect 19824 3111 19858 3139
rect 19824 3071 19858 3073
rect 19824 3039 19858 3071
rect 19824 2969 19858 3001
rect 19824 2967 19858 2969
rect 19824 2901 19858 2929
rect 19824 2895 19858 2901
rect 19824 2833 19858 2857
rect 19824 2823 19858 2833
rect 19824 2765 19858 2785
rect 19824 2751 19858 2765
rect 19824 2697 19858 2713
rect 19824 2679 19858 2697
rect 19824 2629 19858 2641
rect 19824 2607 19858 2629
rect 19824 2561 19858 2569
rect 19824 2535 19858 2561
rect 19920 3479 19954 3505
rect 19920 3471 19954 3479
rect 19920 3411 19954 3433
rect 19920 3399 19954 3411
rect 19920 3343 19954 3361
rect 19920 3327 19954 3343
rect 19920 3275 19954 3289
rect 19920 3255 19954 3275
rect 19920 3207 19954 3217
rect 19920 3183 19954 3207
rect 19920 3139 19954 3145
rect 19920 3111 19954 3139
rect 19920 3071 19954 3073
rect 19920 3039 19954 3071
rect 19920 2969 19954 3001
rect 19920 2967 19954 2969
rect 19920 2901 19954 2929
rect 19920 2895 19954 2901
rect 19920 2833 19954 2857
rect 19920 2823 19954 2833
rect 19920 2765 19954 2785
rect 19920 2751 19954 2765
rect 19920 2697 19954 2713
rect 19920 2679 19954 2697
rect 19920 2629 19954 2641
rect 19920 2607 19954 2629
rect 19920 2561 19954 2569
rect 19920 2535 19954 2561
rect 20016 3479 20050 3505
rect 20016 3471 20050 3479
rect 20016 3411 20050 3433
rect 20016 3399 20050 3411
rect 20016 3343 20050 3361
rect 20016 3327 20050 3343
rect 20016 3275 20050 3289
rect 20016 3255 20050 3275
rect 20016 3207 20050 3217
rect 20016 3183 20050 3207
rect 20016 3139 20050 3145
rect 20016 3111 20050 3139
rect 20016 3071 20050 3073
rect 20016 3039 20050 3071
rect 20016 2969 20050 3001
rect 20016 2967 20050 2969
rect 20016 2901 20050 2929
rect 20016 2895 20050 2901
rect 20016 2833 20050 2857
rect 20016 2823 20050 2833
rect 20016 2765 20050 2785
rect 20016 2751 20050 2765
rect 20016 2697 20050 2713
rect 20016 2679 20050 2697
rect 20016 2629 20050 2641
rect 20016 2607 20050 2629
rect 20016 2561 20050 2569
rect 20016 2535 20050 2561
rect 20244 3487 20278 3513
rect 20244 3479 20278 3487
rect 20244 3419 20278 3441
rect 20244 3407 20278 3419
rect 20244 3351 20278 3369
rect 20244 3335 20278 3351
rect 20244 3283 20278 3297
rect 20244 3263 20278 3283
rect 20244 3215 20278 3225
rect 20244 3191 20278 3215
rect 20244 3147 20278 3153
rect 20244 3119 20278 3147
rect 20244 3079 20278 3081
rect 20244 3047 20278 3079
rect 20244 2977 20278 3009
rect 20244 2975 20278 2977
rect 20244 2909 20278 2937
rect 20244 2903 20278 2909
rect 20244 2841 20278 2865
rect 20244 2831 20278 2841
rect 20244 2773 20278 2793
rect 20244 2759 20278 2773
rect 20244 2705 20278 2721
rect 20244 2687 20278 2705
rect 20244 2637 20278 2649
rect 20244 2615 20278 2637
rect 20244 2569 20278 2577
rect 20244 2543 20278 2569
rect 20340 3487 20374 3513
rect 20340 3479 20374 3487
rect 20340 3419 20374 3441
rect 20340 3407 20374 3419
rect 20340 3351 20374 3369
rect 20340 3335 20374 3351
rect 20340 3283 20374 3297
rect 20340 3263 20374 3283
rect 20340 3215 20374 3225
rect 20340 3191 20374 3215
rect 20340 3147 20374 3153
rect 20340 3119 20374 3147
rect 20340 3079 20374 3081
rect 20340 3047 20374 3079
rect 20340 2977 20374 3009
rect 20340 2975 20374 2977
rect 20340 2909 20374 2937
rect 20340 2903 20374 2909
rect 20340 2841 20374 2865
rect 20340 2831 20374 2841
rect 20340 2773 20374 2793
rect 20340 2759 20374 2773
rect 20340 2705 20374 2721
rect 20340 2687 20374 2705
rect 20340 2637 20374 2649
rect 20340 2615 20374 2637
rect 20340 2569 20374 2577
rect 20340 2543 20374 2569
rect 20436 3487 20470 3513
rect 20436 3479 20470 3487
rect 20436 3419 20470 3441
rect 20436 3407 20470 3419
rect 20436 3351 20470 3369
rect 20436 3335 20470 3351
rect 20436 3283 20470 3297
rect 20436 3263 20470 3283
rect 20436 3215 20470 3225
rect 20436 3191 20470 3215
rect 20436 3147 20470 3153
rect 20436 3119 20470 3147
rect 20436 3079 20470 3081
rect 20436 3047 20470 3079
rect 20436 2977 20470 3009
rect 20436 2975 20470 2977
rect 20436 2909 20470 2937
rect 20436 2903 20470 2909
rect 20436 2841 20470 2865
rect 20436 2831 20470 2841
rect 20436 2773 20470 2793
rect 20436 2759 20470 2773
rect 20436 2705 20470 2721
rect 20436 2687 20470 2705
rect 20436 2637 20470 2649
rect 20436 2615 20470 2637
rect 20436 2569 20470 2577
rect 20436 2543 20470 2569
rect 20532 3487 20566 3513
rect 20532 3479 20566 3487
rect 20532 3419 20566 3441
rect 20532 3407 20566 3419
rect 20532 3351 20566 3369
rect 20532 3335 20566 3351
rect 20532 3283 20566 3297
rect 20532 3263 20566 3283
rect 20532 3215 20566 3225
rect 20532 3191 20566 3215
rect 20532 3147 20566 3153
rect 20532 3119 20566 3147
rect 20532 3079 20566 3081
rect 20532 3047 20566 3079
rect 20532 2977 20566 3009
rect 20532 2975 20566 2977
rect 20532 2909 20566 2937
rect 20532 2903 20566 2909
rect 20532 2841 20566 2865
rect 20532 2831 20566 2841
rect 20532 2773 20566 2793
rect 20532 2759 20566 2773
rect 20532 2705 20566 2721
rect 20532 2687 20566 2705
rect 20532 2637 20566 2649
rect 20532 2615 20566 2637
rect 20532 2569 20566 2577
rect 20532 2543 20566 2569
rect 20628 3487 20662 3513
rect 20628 3479 20662 3487
rect 20628 3419 20662 3441
rect 20628 3407 20662 3419
rect 20628 3351 20662 3369
rect 20628 3335 20662 3351
rect 20628 3283 20662 3297
rect 20628 3263 20662 3283
rect 20628 3215 20662 3225
rect 20628 3191 20662 3215
rect 20628 3147 20662 3153
rect 20628 3119 20662 3147
rect 20628 3079 20662 3081
rect 20628 3047 20662 3079
rect 20628 2977 20662 3009
rect 20628 2975 20662 2977
rect 20628 2909 20662 2937
rect 20628 2903 20662 2909
rect 20628 2841 20662 2865
rect 20628 2831 20662 2841
rect 20628 2773 20662 2793
rect 20628 2759 20662 2773
rect 20628 2705 20662 2721
rect 20628 2687 20662 2705
rect 20628 2637 20662 2649
rect 20628 2615 20662 2637
rect 20628 2569 20662 2577
rect 20628 2543 20662 2569
rect 20724 3487 20758 3513
rect 20724 3479 20758 3487
rect 20724 3419 20758 3441
rect 20724 3407 20758 3419
rect 20724 3351 20758 3369
rect 20724 3335 20758 3351
rect 20724 3283 20758 3297
rect 20724 3263 20758 3283
rect 20724 3215 20758 3225
rect 20724 3191 20758 3215
rect 20724 3147 20758 3153
rect 20724 3119 20758 3147
rect 20724 3079 20758 3081
rect 20724 3047 20758 3079
rect 20724 2977 20758 3009
rect 20724 2975 20758 2977
rect 20724 2909 20758 2937
rect 20724 2903 20758 2909
rect 20724 2841 20758 2865
rect 20724 2831 20758 2841
rect 20724 2773 20758 2793
rect 20724 2759 20758 2773
rect 20724 2705 20758 2721
rect 20724 2687 20758 2705
rect 20724 2637 20758 2649
rect 20724 2615 20758 2637
rect 20724 2569 20758 2577
rect 20724 2543 20758 2569
rect 20820 3487 20854 3513
rect 20820 3479 20854 3487
rect 20820 3419 20854 3441
rect 20820 3407 20854 3419
rect 20820 3351 20854 3369
rect 20820 3335 20854 3351
rect 20820 3283 20854 3297
rect 20820 3263 20854 3283
rect 20820 3215 20854 3225
rect 20820 3191 20854 3215
rect 20820 3147 20854 3153
rect 20820 3119 20854 3147
rect 20820 3079 20854 3081
rect 20820 3047 20854 3079
rect 20820 2977 20854 3009
rect 20820 2975 20854 2977
rect 20820 2909 20854 2937
rect 20820 2903 20854 2909
rect 20820 2841 20854 2865
rect 20820 2831 20854 2841
rect 20820 2773 20854 2793
rect 20820 2759 20854 2773
rect 20820 2705 20854 2721
rect 20820 2687 20854 2705
rect 20820 2637 20854 2649
rect 20820 2615 20854 2637
rect 20820 2569 20854 2577
rect 20820 2543 20854 2569
rect 20916 3487 20950 3513
rect 20916 3479 20950 3487
rect 20916 3419 20950 3441
rect 20916 3407 20950 3419
rect 20916 3351 20950 3369
rect 20916 3335 20950 3351
rect 20916 3283 20950 3297
rect 20916 3263 20950 3283
rect 20916 3215 20950 3225
rect 20916 3191 20950 3215
rect 20916 3147 20950 3153
rect 20916 3119 20950 3147
rect 20916 3079 20950 3081
rect 20916 3047 20950 3079
rect 20916 2977 20950 3009
rect 20916 2975 20950 2977
rect 20916 2909 20950 2937
rect 20916 2903 20950 2909
rect 20916 2841 20950 2865
rect 20916 2831 20950 2841
rect 20916 2773 20950 2793
rect 20916 2759 20950 2773
rect 20916 2705 20950 2721
rect 20916 2687 20950 2705
rect 20916 2637 20950 2649
rect 20916 2615 20950 2637
rect 20916 2569 20950 2577
rect 20916 2543 20950 2569
rect 21012 3487 21046 3513
rect 21012 3479 21046 3487
rect 21012 3419 21046 3441
rect 21012 3407 21046 3419
rect 21012 3351 21046 3369
rect 21012 3335 21046 3351
rect 21012 3283 21046 3297
rect 21012 3263 21046 3283
rect 21012 3215 21046 3225
rect 21012 3191 21046 3215
rect 21012 3147 21046 3153
rect 21012 3119 21046 3147
rect 21012 3079 21046 3081
rect 21012 3047 21046 3079
rect 21012 2977 21046 3009
rect 21012 2975 21046 2977
rect 21012 2909 21046 2937
rect 21012 2903 21046 2909
rect 21012 2841 21046 2865
rect 21012 2831 21046 2841
rect 21012 2773 21046 2793
rect 21012 2759 21046 2773
rect 21012 2705 21046 2721
rect 21012 2687 21046 2705
rect 21012 2637 21046 2649
rect 21012 2615 21046 2637
rect 21012 2569 21046 2577
rect 21012 2543 21046 2569
rect 21108 3487 21142 3513
rect 21108 3479 21142 3487
rect 21108 3419 21142 3441
rect 21108 3407 21142 3419
rect 21108 3351 21142 3369
rect 21108 3335 21142 3351
rect 21108 3283 21142 3297
rect 21108 3263 21142 3283
rect 21108 3215 21142 3225
rect 21108 3191 21142 3215
rect 21108 3147 21142 3153
rect 21108 3119 21142 3147
rect 21108 3079 21142 3081
rect 21108 3047 21142 3079
rect 21108 2977 21142 3009
rect 21108 2975 21142 2977
rect 21108 2909 21142 2937
rect 21108 2903 21142 2909
rect 21108 2841 21142 2865
rect 21108 2831 21142 2841
rect 21108 2773 21142 2793
rect 21108 2759 21142 2773
rect 21108 2705 21142 2721
rect 21108 2687 21142 2705
rect 21108 2637 21142 2649
rect 21108 2615 21142 2637
rect 21108 2569 21142 2577
rect 21108 2543 21142 2569
rect 21204 3487 21238 3513
rect 21204 3479 21238 3487
rect 21204 3419 21238 3441
rect 21204 3407 21238 3419
rect 21204 3351 21238 3369
rect 21204 3335 21238 3351
rect 21204 3283 21238 3297
rect 21204 3263 21238 3283
rect 21204 3215 21238 3225
rect 21204 3191 21238 3215
rect 21204 3147 21238 3153
rect 21204 3119 21238 3147
rect 21204 3079 21238 3081
rect 21204 3047 21238 3079
rect 21204 2977 21238 3009
rect 21204 2975 21238 2977
rect 21204 2909 21238 2937
rect 21204 2903 21238 2909
rect 21204 2841 21238 2865
rect 21204 2831 21238 2841
rect 21204 2773 21238 2793
rect 21204 2759 21238 2773
rect 21204 2705 21238 2721
rect 21204 2687 21238 2705
rect 21204 2637 21238 2649
rect 21204 2615 21238 2637
rect 21204 2569 21238 2577
rect 21204 2543 21238 2569
rect 21300 3487 21334 3513
rect 21300 3479 21334 3487
rect 21300 3419 21334 3441
rect 21300 3407 21334 3419
rect 21300 3351 21334 3369
rect 21300 3335 21334 3351
rect 21300 3283 21334 3297
rect 21300 3263 21334 3283
rect 21300 3215 21334 3225
rect 21300 3191 21334 3215
rect 21300 3147 21334 3153
rect 21300 3119 21334 3147
rect 21300 3079 21334 3081
rect 21300 3047 21334 3079
rect 21300 2977 21334 3009
rect 21300 2975 21334 2977
rect 21300 2909 21334 2937
rect 21300 2903 21334 2909
rect 21300 2841 21334 2865
rect 21300 2831 21334 2841
rect 21300 2773 21334 2793
rect 21300 2759 21334 2773
rect 21300 2705 21334 2721
rect 21300 2687 21334 2705
rect 21300 2637 21334 2649
rect 21300 2615 21334 2637
rect 21300 2569 21334 2577
rect 21300 2543 21334 2569
rect 21396 3487 21430 3513
rect 21396 3479 21430 3487
rect 21396 3419 21430 3441
rect 21396 3407 21430 3419
rect 21396 3351 21430 3369
rect 21396 3335 21430 3351
rect 21396 3283 21430 3297
rect 21396 3263 21430 3283
rect 21396 3215 21430 3225
rect 21396 3191 21430 3215
rect 21396 3147 21430 3153
rect 21396 3119 21430 3147
rect 21396 3079 21430 3081
rect 21396 3047 21430 3079
rect 21396 2977 21430 3009
rect 21396 2975 21430 2977
rect 21396 2909 21430 2937
rect 21396 2903 21430 2909
rect 21396 2841 21430 2865
rect 21396 2831 21430 2841
rect 21396 2773 21430 2793
rect 21396 2759 21430 2773
rect 21396 2705 21430 2721
rect 21396 2687 21430 2705
rect 21396 2637 21430 2649
rect 21396 2615 21430 2637
rect 21396 2569 21430 2577
rect 21396 2543 21430 2569
rect 21492 3487 21526 3513
rect 21492 3479 21526 3487
rect 21492 3419 21526 3441
rect 21492 3407 21526 3419
rect 21492 3351 21526 3369
rect 21492 3335 21526 3351
rect 21492 3283 21526 3297
rect 21492 3263 21526 3283
rect 21492 3215 21526 3225
rect 21492 3191 21526 3215
rect 21492 3147 21526 3153
rect 21492 3119 21526 3147
rect 21492 3079 21526 3081
rect 21492 3047 21526 3079
rect 21492 2977 21526 3009
rect 21492 2975 21526 2977
rect 21492 2909 21526 2937
rect 21492 2903 21526 2909
rect 21492 2841 21526 2865
rect 21492 2831 21526 2841
rect 21492 2773 21526 2793
rect 21492 2759 21526 2773
rect 21492 2705 21526 2721
rect 21492 2687 21526 2705
rect 21492 2637 21526 2649
rect 21492 2615 21526 2637
rect 21492 2569 21526 2577
rect 21492 2543 21526 2569
rect 21588 3487 21622 3513
rect 21588 3479 21622 3487
rect 21588 3419 21622 3441
rect 21588 3407 21622 3419
rect 21588 3351 21622 3369
rect 21588 3335 21622 3351
rect 21588 3283 21622 3297
rect 21588 3263 21622 3283
rect 21588 3215 21622 3225
rect 21588 3191 21622 3215
rect 21588 3147 21622 3153
rect 21588 3119 21622 3147
rect 21588 3079 21622 3081
rect 21588 3047 21622 3079
rect 21588 2977 21622 3009
rect 21588 2975 21622 2977
rect 21588 2909 21622 2937
rect 21588 2903 21622 2909
rect 21588 2841 21622 2865
rect 21588 2831 21622 2841
rect 21588 2773 21622 2793
rect 21588 2759 21622 2773
rect 21588 2705 21622 2721
rect 21588 2687 21622 2705
rect 21588 2637 21622 2649
rect 21588 2615 21622 2637
rect 21588 2569 21622 2577
rect 21588 2543 21622 2569
rect 21684 3487 21718 3513
rect 21684 3479 21718 3487
rect 21684 3419 21718 3441
rect 21684 3407 21718 3419
rect 21684 3351 21718 3369
rect 21684 3335 21718 3351
rect 21684 3283 21718 3297
rect 21684 3263 21718 3283
rect 21684 3215 21718 3225
rect 21684 3191 21718 3215
rect 21684 3147 21718 3153
rect 21684 3119 21718 3147
rect 21684 3079 21718 3081
rect 21684 3047 21718 3079
rect 21684 2977 21718 3009
rect 21684 2975 21718 2977
rect 21684 2909 21718 2937
rect 21684 2903 21718 2909
rect 21684 2841 21718 2865
rect 21684 2831 21718 2841
rect 21684 2773 21718 2793
rect 21684 2759 21718 2773
rect 21684 2705 21718 2721
rect 21684 2687 21718 2705
rect 21684 2637 21718 2649
rect 21684 2615 21718 2637
rect 21684 2569 21718 2577
rect 21684 2543 21718 2569
rect 21780 3487 21814 3513
rect 21780 3479 21814 3487
rect 21780 3419 21814 3441
rect 21780 3407 21814 3419
rect 21780 3351 21814 3369
rect 21780 3335 21814 3351
rect 21780 3283 21814 3297
rect 21780 3263 21814 3283
rect 21780 3215 21814 3225
rect 21780 3191 21814 3215
rect 21780 3147 21814 3153
rect 21780 3119 21814 3147
rect 21780 3079 21814 3081
rect 21780 3047 21814 3079
rect 21780 2977 21814 3009
rect 21780 2975 21814 2977
rect 21780 2909 21814 2937
rect 21780 2903 21814 2909
rect 21780 2841 21814 2865
rect 21780 2831 21814 2841
rect 21780 2773 21814 2793
rect 21780 2759 21814 2773
rect 21780 2705 21814 2721
rect 21780 2687 21814 2705
rect 21780 2637 21814 2649
rect 21780 2615 21814 2637
rect 21780 2569 21814 2577
rect 21780 2543 21814 2569
rect 21876 3487 21910 3513
rect 21876 3479 21910 3487
rect 21876 3419 21910 3441
rect 21876 3407 21910 3419
rect 21876 3351 21910 3369
rect 21876 3335 21910 3351
rect 21876 3283 21910 3297
rect 21876 3263 21910 3283
rect 21876 3215 21910 3225
rect 21876 3191 21910 3215
rect 21876 3147 21910 3153
rect 21876 3119 21910 3147
rect 21876 3079 21910 3081
rect 21876 3047 21910 3079
rect 21876 2977 21910 3009
rect 21876 2975 21910 2977
rect 21876 2909 21910 2937
rect 21876 2903 21910 2909
rect 21876 2841 21910 2865
rect 21876 2831 21910 2841
rect 21876 2773 21910 2793
rect 21876 2759 21910 2773
rect 21876 2705 21910 2721
rect 21876 2687 21910 2705
rect 21876 2637 21910 2649
rect 21876 2615 21910 2637
rect 21876 2569 21910 2577
rect 21876 2543 21910 2569
rect 21972 3487 22006 3513
rect 21972 3479 22006 3487
rect 21972 3419 22006 3441
rect 21972 3407 22006 3419
rect 21972 3351 22006 3369
rect 21972 3335 22006 3351
rect 21972 3283 22006 3297
rect 21972 3263 22006 3283
rect 21972 3215 22006 3225
rect 21972 3191 22006 3215
rect 21972 3147 22006 3153
rect 21972 3119 22006 3147
rect 21972 3079 22006 3081
rect 21972 3047 22006 3079
rect 21972 2977 22006 3009
rect 21972 2975 22006 2977
rect 21972 2909 22006 2937
rect 21972 2903 22006 2909
rect 21972 2841 22006 2865
rect 21972 2831 22006 2841
rect 21972 2773 22006 2793
rect 21972 2759 22006 2773
rect 21972 2705 22006 2721
rect 21972 2687 22006 2705
rect 21972 2637 22006 2649
rect 21972 2615 22006 2637
rect 21972 2569 22006 2577
rect 21972 2543 22006 2569
rect 22068 3487 22102 3513
rect 22068 3479 22102 3487
rect 22068 3419 22102 3441
rect 22068 3407 22102 3419
rect 22068 3351 22102 3369
rect 22068 3335 22102 3351
rect 22068 3283 22102 3297
rect 22068 3263 22102 3283
rect 22068 3215 22102 3225
rect 22068 3191 22102 3215
rect 22068 3147 22102 3153
rect 22068 3119 22102 3147
rect 22068 3079 22102 3081
rect 22068 3047 22102 3079
rect 22068 2977 22102 3009
rect 22068 2975 22102 2977
rect 22068 2909 22102 2937
rect 22068 2903 22102 2909
rect 22068 2841 22102 2865
rect 22068 2831 22102 2841
rect 22068 2773 22102 2793
rect 22068 2759 22102 2773
rect 22068 2705 22102 2721
rect 22068 2687 22102 2705
rect 22068 2637 22102 2649
rect 22068 2615 22102 2637
rect 22068 2569 22102 2577
rect 22068 2543 22102 2569
rect 22164 3487 22198 3513
rect 22164 3479 22198 3487
rect 22164 3419 22198 3441
rect 22164 3407 22198 3419
rect 22164 3351 22198 3369
rect 22164 3335 22198 3351
rect 22164 3283 22198 3297
rect 22164 3263 22198 3283
rect 22164 3215 22198 3225
rect 22164 3191 22198 3215
rect 22164 3147 22198 3153
rect 22164 3119 22198 3147
rect 22164 3079 22198 3081
rect 22164 3047 22198 3079
rect 22164 2977 22198 3009
rect 22164 2975 22198 2977
rect 22164 2909 22198 2937
rect 22164 2903 22198 2909
rect 22164 2841 22198 2865
rect 22164 2831 22198 2841
rect 22164 2773 22198 2793
rect 22164 2759 22198 2773
rect 22164 2705 22198 2721
rect 22164 2687 22198 2705
rect 22164 2637 22198 2649
rect 22164 2615 22198 2637
rect 22164 2569 22198 2577
rect 22164 2543 22198 2569
rect 23174 3491 23208 3517
rect 23174 3483 23208 3491
rect 23174 3423 23208 3445
rect 23174 3411 23208 3423
rect 23174 3355 23208 3373
rect 23174 3339 23208 3355
rect 23174 3287 23208 3301
rect 23174 3267 23208 3287
rect 23174 3219 23208 3229
rect 23174 3195 23208 3219
rect 23174 3151 23208 3157
rect 23174 3123 23208 3151
rect 23174 3083 23208 3085
rect 23174 3051 23208 3083
rect 23174 2981 23208 3013
rect 23174 2979 23208 2981
rect 23174 2913 23208 2941
rect 23174 2907 23208 2913
rect 23174 2845 23208 2869
rect 23174 2835 23208 2845
rect 23174 2777 23208 2797
rect 23174 2763 23208 2777
rect 23174 2709 23208 2725
rect 23174 2691 23208 2709
rect 23174 2641 23208 2653
rect 23174 2619 23208 2641
rect 23174 2573 23208 2581
rect 23174 2547 23208 2573
rect 23270 3491 23304 3517
rect 23270 3483 23304 3491
rect 23270 3423 23304 3445
rect 23270 3411 23304 3423
rect 23270 3355 23304 3373
rect 23270 3339 23304 3355
rect 23270 3287 23304 3301
rect 23270 3267 23304 3287
rect 23270 3219 23304 3229
rect 23270 3195 23304 3219
rect 23270 3151 23304 3157
rect 23270 3123 23304 3151
rect 23270 3083 23304 3085
rect 23270 3051 23304 3083
rect 23270 2981 23304 3013
rect 23270 2979 23304 2981
rect 23270 2913 23304 2941
rect 23270 2907 23304 2913
rect 23270 2845 23304 2869
rect 23270 2835 23304 2845
rect 23270 2777 23304 2797
rect 23270 2763 23304 2777
rect 23270 2709 23304 2725
rect 23270 2691 23304 2709
rect 23270 2641 23304 2653
rect 23270 2619 23304 2641
rect 23270 2573 23304 2581
rect 23270 2547 23304 2573
rect 23366 3491 23400 3517
rect 23366 3483 23400 3491
rect 23366 3423 23400 3445
rect 23366 3411 23400 3423
rect 23366 3355 23400 3373
rect 23366 3339 23400 3355
rect 23366 3287 23400 3301
rect 23366 3267 23400 3287
rect 23366 3219 23400 3229
rect 23366 3195 23400 3219
rect 23366 3151 23400 3157
rect 23366 3123 23400 3151
rect 23366 3083 23400 3085
rect 23366 3051 23400 3083
rect 23366 2981 23400 3013
rect 23366 2979 23400 2981
rect 23366 2913 23400 2941
rect 23366 2907 23400 2913
rect 23366 2845 23400 2869
rect 23366 2835 23400 2845
rect 23366 2777 23400 2797
rect 23366 2763 23400 2777
rect 23366 2709 23400 2725
rect 23366 2691 23400 2709
rect 23366 2641 23400 2653
rect 23366 2619 23400 2641
rect 23366 2573 23400 2581
rect 23366 2547 23400 2573
rect 23462 3491 23496 3517
rect 23462 3483 23496 3491
rect 23462 3423 23496 3445
rect 23462 3411 23496 3423
rect 23462 3355 23496 3373
rect 23462 3339 23496 3355
rect 23462 3287 23496 3301
rect 23462 3267 23496 3287
rect 23462 3219 23496 3229
rect 23462 3195 23496 3219
rect 23462 3151 23496 3157
rect 23462 3123 23496 3151
rect 23462 3083 23496 3085
rect 23462 3051 23496 3083
rect 23462 2981 23496 3013
rect 23462 2979 23496 2981
rect 23462 2913 23496 2941
rect 23462 2907 23496 2913
rect 23462 2845 23496 2869
rect 23462 2835 23496 2845
rect 23462 2777 23496 2797
rect 23462 2763 23496 2777
rect 23462 2709 23496 2725
rect 23462 2691 23496 2709
rect 23462 2641 23496 2653
rect 23462 2619 23496 2641
rect 23462 2573 23496 2581
rect 23462 2547 23496 2573
rect 23558 3491 23592 3517
rect 23558 3483 23592 3491
rect 23558 3423 23592 3445
rect 23558 3411 23592 3423
rect 23558 3355 23592 3373
rect 23558 3339 23592 3355
rect 23558 3287 23592 3301
rect 23558 3267 23592 3287
rect 23558 3219 23592 3229
rect 23558 3195 23592 3219
rect 23558 3151 23592 3157
rect 23558 3123 23592 3151
rect 23558 3083 23592 3085
rect 23558 3051 23592 3083
rect 23558 2981 23592 3013
rect 23558 2979 23592 2981
rect 23558 2913 23592 2941
rect 23558 2907 23592 2913
rect 23558 2845 23592 2869
rect 23558 2835 23592 2845
rect 23558 2777 23592 2797
rect 23558 2763 23592 2777
rect 23558 2709 23592 2725
rect 23558 2691 23592 2709
rect 23558 2641 23592 2653
rect 23558 2619 23592 2641
rect 23558 2573 23592 2581
rect 23558 2547 23592 2573
rect 28134 3768 28168 3802
rect 26876 3654 26910 3688
rect 23654 3491 23688 3517
rect 23654 3483 23688 3491
rect 23654 3423 23688 3445
rect 23654 3411 23688 3423
rect 23654 3355 23688 3373
rect 23654 3339 23688 3355
rect 23654 3287 23688 3301
rect 23654 3267 23688 3287
rect 23654 3219 23688 3229
rect 23654 3195 23688 3219
rect 23654 3151 23688 3157
rect 23654 3123 23688 3151
rect 23654 3083 23688 3085
rect 23654 3051 23688 3083
rect 23654 2981 23688 3013
rect 23654 2979 23688 2981
rect 23654 2913 23688 2941
rect 23654 2907 23688 2913
rect 23654 2845 23688 2869
rect 23654 2835 23688 2845
rect 23654 2777 23688 2797
rect 23654 2763 23688 2777
rect 23654 2709 23688 2725
rect 23654 2691 23688 2709
rect 23654 2641 23688 2653
rect 23654 2619 23688 2641
rect 23654 2573 23688 2581
rect 23654 2547 23688 2573
rect 23866 3481 23900 3507
rect 23866 3473 23900 3481
rect 23866 3413 23900 3435
rect 23866 3401 23900 3413
rect 23866 3345 23900 3363
rect 23866 3329 23900 3345
rect 23866 3277 23900 3291
rect 23866 3257 23900 3277
rect 23866 3209 23900 3219
rect 23866 3185 23900 3209
rect 23866 3141 23900 3147
rect 23866 3113 23900 3141
rect 23866 3073 23900 3075
rect 23866 3041 23900 3073
rect 23866 2971 23900 3003
rect 23866 2969 23900 2971
rect 23866 2903 23900 2931
rect 23866 2897 23900 2903
rect 23866 2835 23900 2859
rect 23866 2825 23900 2835
rect 23866 2767 23900 2787
rect 23866 2753 23900 2767
rect 23866 2699 23900 2715
rect 23866 2681 23900 2699
rect 23866 2631 23900 2643
rect 23866 2609 23900 2631
rect 23866 2563 23900 2571
rect 23866 2537 23900 2563
rect 23962 3481 23996 3507
rect 23962 3473 23996 3481
rect 23962 3413 23996 3435
rect 23962 3401 23996 3413
rect 23962 3345 23996 3363
rect 23962 3329 23996 3345
rect 23962 3277 23996 3291
rect 23962 3257 23996 3277
rect 23962 3209 23996 3219
rect 23962 3185 23996 3209
rect 23962 3141 23996 3147
rect 23962 3113 23996 3141
rect 23962 3073 23996 3075
rect 23962 3041 23996 3073
rect 23962 2971 23996 3003
rect 23962 2969 23996 2971
rect 23962 2903 23996 2931
rect 23962 2897 23996 2903
rect 23962 2835 23996 2859
rect 23962 2825 23996 2835
rect 23962 2767 23996 2787
rect 23962 2753 23996 2767
rect 23962 2699 23996 2715
rect 23962 2681 23996 2699
rect 23962 2631 23996 2643
rect 23962 2609 23996 2631
rect 23962 2563 23996 2571
rect 23962 2537 23996 2563
rect 24058 3481 24092 3507
rect 24058 3473 24092 3481
rect 24058 3413 24092 3435
rect 24058 3401 24092 3413
rect 24058 3345 24092 3363
rect 24058 3329 24092 3345
rect 24058 3277 24092 3291
rect 24058 3257 24092 3277
rect 24058 3209 24092 3219
rect 24058 3185 24092 3209
rect 24058 3141 24092 3147
rect 24058 3113 24092 3141
rect 24058 3073 24092 3075
rect 24058 3041 24092 3073
rect 24058 2971 24092 3003
rect 24058 2969 24092 2971
rect 24058 2903 24092 2931
rect 24058 2897 24092 2903
rect 24058 2835 24092 2859
rect 24058 2825 24092 2835
rect 24058 2767 24092 2787
rect 24058 2753 24092 2767
rect 24058 2699 24092 2715
rect 24058 2681 24092 2699
rect 24058 2631 24092 2643
rect 24058 2609 24092 2631
rect 24058 2563 24092 2571
rect 24058 2537 24092 2563
rect 24154 3481 24188 3507
rect 24154 3473 24188 3481
rect 24154 3413 24188 3435
rect 24154 3401 24188 3413
rect 24154 3345 24188 3363
rect 24154 3329 24188 3345
rect 24154 3277 24188 3291
rect 24154 3257 24188 3277
rect 24154 3209 24188 3219
rect 24154 3185 24188 3209
rect 24154 3141 24188 3147
rect 24154 3113 24188 3141
rect 24154 3073 24188 3075
rect 24154 3041 24188 3073
rect 24154 2971 24188 3003
rect 24154 2969 24188 2971
rect 24154 2903 24188 2931
rect 24154 2897 24188 2903
rect 24154 2835 24188 2859
rect 24154 2825 24188 2835
rect 24154 2767 24188 2787
rect 24154 2753 24188 2767
rect 24154 2699 24188 2715
rect 24154 2681 24188 2699
rect 24154 2631 24188 2643
rect 24154 2609 24188 2631
rect 24154 2563 24188 2571
rect 24154 2537 24188 2563
rect 24250 3481 24284 3507
rect 24250 3473 24284 3481
rect 24250 3413 24284 3435
rect 24250 3401 24284 3413
rect 24250 3345 24284 3363
rect 24250 3329 24284 3345
rect 24250 3277 24284 3291
rect 24250 3257 24284 3277
rect 24250 3209 24284 3219
rect 24250 3185 24284 3209
rect 24250 3141 24284 3147
rect 24250 3113 24284 3141
rect 24250 3073 24284 3075
rect 24250 3041 24284 3073
rect 24250 2971 24284 3003
rect 24250 2969 24284 2971
rect 24250 2903 24284 2931
rect 24250 2897 24284 2903
rect 24250 2835 24284 2859
rect 24250 2825 24284 2835
rect 24250 2767 24284 2787
rect 24250 2753 24284 2767
rect 24250 2699 24284 2715
rect 24250 2681 24284 2699
rect 24250 2631 24284 2643
rect 24250 2609 24284 2631
rect 24250 2563 24284 2571
rect 24250 2537 24284 2563
rect 24346 3481 24380 3507
rect 24346 3473 24380 3481
rect 24346 3413 24380 3435
rect 24346 3401 24380 3413
rect 24346 3345 24380 3363
rect 24346 3329 24380 3345
rect 24346 3277 24380 3291
rect 24346 3257 24380 3277
rect 24346 3209 24380 3219
rect 24346 3185 24380 3209
rect 24346 3141 24380 3147
rect 24346 3113 24380 3141
rect 24346 3073 24380 3075
rect 24346 3041 24380 3073
rect 24346 2971 24380 3003
rect 24346 2969 24380 2971
rect 24346 2903 24380 2931
rect 24346 2897 24380 2903
rect 24346 2835 24380 2859
rect 24346 2825 24380 2835
rect 24346 2767 24380 2787
rect 24346 2753 24380 2767
rect 24346 2699 24380 2715
rect 24346 2681 24380 2699
rect 24346 2631 24380 2643
rect 24346 2609 24380 2631
rect 24346 2563 24380 2571
rect 24346 2537 24380 2563
rect 24442 3481 24476 3507
rect 24442 3473 24476 3481
rect 24442 3413 24476 3435
rect 24442 3401 24476 3413
rect 24442 3345 24476 3363
rect 24442 3329 24476 3345
rect 24442 3277 24476 3291
rect 24442 3257 24476 3277
rect 24442 3209 24476 3219
rect 24442 3185 24476 3209
rect 24442 3141 24476 3147
rect 24442 3113 24476 3141
rect 24442 3073 24476 3075
rect 24442 3041 24476 3073
rect 24442 2971 24476 3003
rect 24442 2969 24476 2971
rect 24442 2903 24476 2931
rect 24442 2897 24476 2903
rect 24442 2835 24476 2859
rect 24442 2825 24476 2835
rect 24442 2767 24476 2787
rect 24442 2753 24476 2767
rect 24442 2699 24476 2715
rect 24442 2681 24476 2699
rect 24442 2631 24476 2643
rect 24442 2609 24476 2631
rect 24442 2563 24476 2571
rect 24442 2537 24476 2563
rect 24538 3481 24572 3507
rect 24538 3473 24572 3481
rect 24538 3413 24572 3435
rect 24538 3401 24572 3413
rect 24538 3345 24572 3363
rect 24538 3329 24572 3345
rect 24538 3277 24572 3291
rect 24538 3257 24572 3277
rect 24538 3209 24572 3219
rect 24538 3185 24572 3209
rect 24538 3141 24572 3147
rect 24538 3113 24572 3141
rect 24538 3073 24572 3075
rect 24538 3041 24572 3073
rect 24538 2971 24572 3003
rect 24538 2969 24572 2971
rect 24538 2903 24572 2931
rect 24538 2897 24572 2903
rect 24538 2835 24572 2859
rect 24538 2825 24572 2835
rect 24538 2767 24572 2787
rect 24538 2753 24572 2767
rect 24538 2699 24572 2715
rect 24538 2681 24572 2699
rect 24538 2631 24572 2643
rect 24538 2609 24572 2631
rect 24538 2563 24572 2571
rect 24538 2537 24572 2563
rect 24634 3481 24668 3507
rect 24634 3473 24668 3481
rect 24634 3413 24668 3435
rect 24634 3401 24668 3413
rect 24634 3345 24668 3363
rect 24634 3329 24668 3345
rect 24634 3277 24668 3291
rect 24634 3257 24668 3277
rect 24634 3209 24668 3219
rect 24634 3185 24668 3209
rect 24634 3141 24668 3147
rect 24634 3113 24668 3141
rect 24634 3073 24668 3075
rect 24634 3041 24668 3073
rect 24634 2971 24668 3003
rect 24634 2969 24668 2971
rect 24634 2903 24668 2931
rect 24634 2897 24668 2903
rect 24634 2835 24668 2859
rect 24634 2825 24668 2835
rect 24634 2767 24668 2787
rect 24634 2753 24668 2767
rect 24634 2699 24668 2715
rect 24634 2681 24668 2699
rect 24634 2631 24668 2643
rect 24634 2609 24668 2631
rect 24634 2563 24668 2571
rect 24634 2537 24668 2563
rect 24730 3481 24764 3507
rect 24730 3473 24764 3481
rect 24730 3413 24764 3435
rect 24730 3401 24764 3413
rect 24730 3345 24764 3363
rect 24730 3329 24764 3345
rect 24730 3277 24764 3291
rect 24730 3257 24764 3277
rect 24730 3209 24764 3219
rect 24730 3185 24764 3209
rect 24730 3141 24764 3147
rect 24730 3113 24764 3141
rect 24730 3073 24764 3075
rect 24730 3041 24764 3073
rect 24730 2971 24764 3003
rect 24730 2969 24764 2971
rect 24730 2903 24764 2931
rect 24730 2897 24764 2903
rect 24730 2835 24764 2859
rect 24730 2825 24764 2835
rect 24730 2767 24764 2787
rect 24730 2753 24764 2767
rect 24730 2699 24764 2715
rect 24730 2681 24764 2699
rect 24730 2631 24764 2643
rect 24730 2609 24764 2631
rect 24730 2563 24764 2571
rect 24730 2537 24764 2563
rect 24826 3481 24860 3507
rect 24826 3473 24860 3481
rect 24826 3413 24860 3435
rect 24826 3401 24860 3413
rect 24826 3345 24860 3363
rect 24826 3329 24860 3345
rect 24826 3277 24860 3291
rect 24826 3257 24860 3277
rect 24826 3209 24860 3219
rect 24826 3185 24860 3209
rect 24826 3141 24860 3147
rect 24826 3113 24860 3141
rect 24826 3073 24860 3075
rect 24826 3041 24860 3073
rect 24826 2971 24860 3003
rect 24826 2969 24860 2971
rect 24826 2903 24860 2931
rect 24826 2897 24860 2903
rect 24826 2835 24860 2859
rect 24826 2825 24860 2835
rect 24826 2767 24860 2787
rect 24826 2753 24860 2767
rect 24826 2699 24860 2715
rect 24826 2681 24860 2699
rect 24826 2631 24860 2643
rect 24826 2609 24860 2631
rect 24826 2563 24860 2571
rect 24826 2537 24860 2563
rect 25064 3477 25098 3503
rect 25064 3469 25098 3477
rect 25064 3409 25098 3431
rect 25064 3397 25098 3409
rect 25064 3341 25098 3359
rect 25064 3325 25098 3341
rect 25064 3273 25098 3287
rect 25064 3253 25098 3273
rect 25064 3205 25098 3215
rect 25064 3181 25098 3205
rect 25064 3137 25098 3143
rect 25064 3109 25098 3137
rect 25064 3069 25098 3071
rect 25064 3037 25098 3069
rect 25064 2967 25098 2999
rect 25064 2965 25098 2967
rect 25064 2899 25098 2927
rect 25064 2893 25098 2899
rect 25064 2831 25098 2855
rect 25064 2821 25098 2831
rect 25064 2763 25098 2783
rect 25064 2749 25098 2763
rect 25064 2695 25098 2711
rect 25064 2677 25098 2695
rect 25064 2627 25098 2639
rect 25064 2605 25098 2627
rect 25064 2559 25098 2567
rect 25064 2533 25098 2559
rect 25160 3477 25194 3503
rect 25160 3469 25194 3477
rect 25160 3409 25194 3431
rect 25160 3397 25194 3409
rect 25160 3341 25194 3359
rect 25160 3325 25194 3341
rect 25160 3273 25194 3287
rect 25160 3253 25194 3273
rect 25160 3205 25194 3215
rect 25160 3181 25194 3205
rect 25160 3137 25194 3143
rect 25160 3109 25194 3137
rect 25160 3069 25194 3071
rect 25160 3037 25194 3069
rect 25160 2967 25194 2999
rect 25160 2965 25194 2967
rect 25160 2899 25194 2927
rect 25160 2893 25194 2899
rect 25160 2831 25194 2855
rect 25160 2821 25194 2831
rect 25160 2763 25194 2783
rect 25160 2749 25194 2763
rect 25160 2695 25194 2711
rect 25160 2677 25194 2695
rect 25160 2627 25194 2639
rect 25160 2605 25194 2627
rect 25160 2559 25194 2567
rect 25160 2533 25194 2559
rect 25256 3477 25290 3503
rect 25256 3469 25290 3477
rect 25256 3409 25290 3431
rect 25256 3397 25290 3409
rect 25256 3341 25290 3359
rect 25256 3325 25290 3341
rect 25256 3273 25290 3287
rect 25256 3253 25290 3273
rect 25256 3205 25290 3215
rect 25256 3181 25290 3205
rect 25256 3137 25290 3143
rect 25256 3109 25290 3137
rect 25256 3069 25290 3071
rect 25256 3037 25290 3069
rect 25256 2967 25290 2999
rect 25256 2965 25290 2967
rect 25256 2899 25290 2927
rect 25256 2893 25290 2899
rect 25256 2831 25290 2855
rect 25256 2821 25290 2831
rect 25256 2763 25290 2783
rect 25256 2749 25290 2763
rect 25256 2695 25290 2711
rect 25256 2677 25290 2695
rect 25256 2627 25290 2639
rect 25256 2605 25290 2627
rect 25256 2559 25290 2567
rect 25256 2533 25290 2559
rect 25352 3477 25386 3503
rect 25352 3469 25386 3477
rect 25352 3409 25386 3431
rect 25352 3397 25386 3409
rect 25352 3341 25386 3359
rect 25352 3325 25386 3341
rect 25352 3273 25386 3287
rect 25352 3253 25386 3273
rect 25352 3205 25386 3215
rect 25352 3181 25386 3205
rect 25352 3137 25386 3143
rect 25352 3109 25386 3137
rect 25352 3069 25386 3071
rect 25352 3037 25386 3069
rect 25352 2967 25386 2999
rect 25352 2965 25386 2967
rect 25352 2899 25386 2927
rect 25352 2893 25386 2899
rect 25352 2831 25386 2855
rect 25352 2821 25386 2831
rect 25352 2763 25386 2783
rect 25352 2749 25386 2763
rect 25352 2695 25386 2711
rect 25352 2677 25386 2695
rect 25352 2627 25386 2639
rect 25352 2605 25386 2627
rect 25352 2559 25386 2567
rect 25352 2533 25386 2559
rect 25448 3477 25482 3503
rect 25448 3469 25482 3477
rect 25448 3409 25482 3431
rect 25448 3397 25482 3409
rect 25448 3341 25482 3359
rect 25448 3325 25482 3341
rect 25448 3273 25482 3287
rect 25448 3253 25482 3273
rect 25448 3205 25482 3215
rect 25448 3181 25482 3205
rect 25448 3137 25482 3143
rect 25448 3109 25482 3137
rect 25448 3069 25482 3071
rect 25448 3037 25482 3069
rect 25448 2967 25482 2999
rect 25448 2965 25482 2967
rect 25448 2899 25482 2927
rect 25448 2893 25482 2899
rect 25448 2831 25482 2855
rect 25448 2821 25482 2831
rect 25448 2763 25482 2783
rect 25448 2749 25482 2763
rect 25448 2695 25482 2711
rect 25448 2677 25482 2695
rect 25448 2627 25482 2639
rect 25448 2605 25482 2627
rect 25448 2559 25482 2567
rect 25448 2533 25482 2559
rect 25544 3477 25578 3503
rect 25544 3469 25578 3477
rect 25544 3409 25578 3431
rect 25544 3397 25578 3409
rect 25544 3341 25578 3359
rect 25544 3325 25578 3341
rect 25544 3273 25578 3287
rect 25544 3253 25578 3273
rect 25544 3205 25578 3215
rect 25544 3181 25578 3205
rect 25544 3137 25578 3143
rect 25544 3109 25578 3137
rect 25544 3069 25578 3071
rect 25544 3037 25578 3069
rect 25544 2967 25578 2999
rect 25544 2965 25578 2967
rect 25544 2899 25578 2927
rect 25544 2893 25578 2899
rect 25544 2831 25578 2855
rect 25544 2821 25578 2831
rect 25544 2763 25578 2783
rect 25544 2749 25578 2763
rect 25544 2695 25578 2711
rect 25544 2677 25578 2695
rect 25544 2627 25578 2639
rect 25544 2605 25578 2627
rect 25544 2559 25578 2567
rect 25544 2533 25578 2559
rect 25640 3477 25674 3503
rect 25640 3469 25674 3477
rect 25640 3409 25674 3431
rect 25640 3397 25674 3409
rect 25640 3341 25674 3359
rect 25640 3325 25674 3341
rect 25640 3273 25674 3287
rect 25640 3253 25674 3273
rect 25640 3205 25674 3215
rect 25640 3181 25674 3205
rect 25640 3137 25674 3143
rect 25640 3109 25674 3137
rect 25640 3069 25674 3071
rect 25640 3037 25674 3069
rect 25640 2967 25674 2999
rect 25640 2965 25674 2967
rect 25640 2899 25674 2927
rect 25640 2893 25674 2899
rect 25640 2831 25674 2855
rect 25640 2821 25674 2831
rect 25640 2763 25674 2783
rect 25640 2749 25674 2763
rect 25640 2695 25674 2711
rect 25640 2677 25674 2695
rect 25640 2627 25674 2639
rect 25640 2605 25674 2627
rect 25640 2559 25674 2567
rect 25640 2533 25674 2559
rect 25736 3477 25770 3503
rect 25736 3469 25770 3477
rect 25736 3409 25770 3431
rect 25736 3397 25770 3409
rect 25736 3341 25770 3359
rect 25736 3325 25770 3341
rect 25736 3273 25770 3287
rect 25736 3253 25770 3273
rect 25736 3205 25770 3215
rect 25736 3181 25770 3205
rect 25736 3137 25770 3143
rect 25736 3109 25770 3137
rect 25736 3069 25770 3071
rect 25736 3037 25770 3069
rect 25736 2967 25770 2999
rect 25736 2965 25770 2967
rect 25736 2899 25770 2927
rect 25736 2893 25770 2899
rect 25736 2831 25770 2855
rect 25736 2821 25770 2831
rect 25736 2763 25770 2783
rect 25736 2749 25770 2763
rect 25736 2695 25770 2711
rect 25736 2677 25770 2695
rect 25736 2627 25770 2639
rect 25736 2605 25770 2627
rect 25736 2559 25770 2567
rect 25736 2533 25770 2559
rect 25832 3477 25866 3503
rect 25832 3469 25866 3477
rect 25832 3409 25866 3431
rect 25832 3397 25866 3409
rect 25832 3341 25866 3359
rect 25832 3325 25866 3341
rect 25832 3273 25866 3287
rect 25832 3253 25866 3273
rect 25832 3205 25866 3215
rect 25832 3181 25866 3205
rect 25832 3137 25866 3143
rect 25832 3109 25866 3137
rect 25832 3069 25866 3071
rect 25832 3037 25866 3069
rect 25832 2967 25866 2999
rect 25832 2965 25866 2967
rect 25832 2899 25866 2927
rect 25832 2893 25866 2899
rect 25832 2831 25866 2855
rect 25832 2821 25866 2831
rect 25832 2763 25866 2783
rect 25832 2749 25866 2763
rect 25832 2695 25866 2711
rect 25832 2677 25866 2695
rect 25832 2627 25866 2639
rect 25832 2605 25866 2627
rect 25832 2559 25866 2567
rect 25832 2533 25866 2559
rect 25928 3477 25962 3503
rect 25928 3469 25962 3477
rect 25928 3409 25962 3431
rect 25928 3397 25962 3409
rect 25928 3341 25962 3359
rect 25928 3325 25962 3341
rect 25928 3273 25962 3287
rect 25928 3253 25962 3273
rect 25928 3205 25962 3215
rect 25928 3181 25962 3205
rect 25928 3137 25962 3143
rect 25928 3109 25962 3137
rect 25928 3069 25962 3071
rect 25928 3037 25962 3069
rect 25928 2967 25962 2999
rect 25928 2965 25962 2967
rect 25928 2899 25962 2927
rect 25928 2893 25962 2899
rect 25928 2831 25962 2855
rect 25928 2821 25962 2831
rect 25928 2763 25962 2783
rect 25928 2749 25962 2763
rect 25928 2695 25962 2711
rect 25928 2677 25962 2695
rect 25928 2627 25962 2639
rect 25928 2605 25962 2627
rect 25928 2559 25962 2567
rect 25928 2533 25962 2559
rect 26024 3477 26058 3503
rect 26024 3469 26058 3477
rect 26024 3409 26058 3431
rect 26024 3397 26058 3409
rect 26024 3341 26058 3359
rect 26024 3325 26058 3341
rect 26024 3273 26058 3287
rect 26024 3253 26058 3273
rect 26024 3205 26058 3215
rect 26024 3181 26058 3205
rect 26024 3137 26058 3143
rect 26024 3109 26058 3137
rect 26024 3069 26058 3071
rect 26024 3037 26058 3069
rect 26024 2967 26058 2999
rect 26024 2965 26058 2967
rect 26024 2899 26058 2927
rect 26024 2893 26058 2899
rect 26024 2831 26058 2855
rect 26024 2821 26058 2831
rect 26024 2763 26058 2783
rect 26024 2749 26058 2763
rect 26024 2695 26058 2711
rect 26024 2677 26058 2695
rect 26024 2627 26058 2639
rect 26024 2605 26058 2627
rect 26024 2559 26058 2567
rect 26024 2533 26058 2559
rect 26120 3477 26154 3503
rect 26120 3469 26154 3477
rect 26120 3409 26154 3431
rect 26120 3397 26154 3409
rect 26120 3341 26154 3359
rect 26120 3325 26154 3341
rect 26120 3273 26154 3287
rect 26120 3253 26154 3273
rect 26120 3205 26154 3215
rect 26120 3181 26154 3205
rect 26120 3137 26154 3143
rect 26120 3109 26154 3137
rect 26120 3069 26154 3071
rect 26120 3037 26154 3069
rect 26120 2967 26154 2999
rect 26120 2965 26154 2967
rect 26120 2899 26154 2927
rect 26120 2893 26154 2899
rect 26120 2831 26154 2855
rect 26120 2821 26154 2831
rect 26120 2763 26154 2783
rect 26120 2749 26154 2763
rect 26120 2695 26154 2711
rect 26120 2677 26154 2695
rect 26120 2627 26154 2639
rect 26120 2605 26154 2627
rect 26120 2559 26154 2567
rect 26120 2533 26154 2559
rect 26216 3477 26250 3503
rect 26216 3469 26250 3477
rect 26216 3409 26250 3431
rect 26216 3397 26250 3409
rect 26216 3341 26250 3359
rect 26216 3325 26250 3341
rect 26216 3273 26250 3287
rect 26216 3253 26250 3273
rect 26216 3205 26250 3215
rect 26216 3181 26250 3205
rect 26216 3137 26250 3143
rect 26216 3109 26250 3137
rect 26216 3069 26250 3071
rect 26216 3037 26250 3069
rect 26216 2967 26250 2999
rect 26216 2965 26250 2967
rect 26216 2899 26250 2927
rect 26216 2893 26250 2899
rect 26216 2831 26250 2855
rect 26216 2821 26250 2831
rect 26216 2763 26250 2783
rect 26216 2749 26250 2763
rect 26216 2695 26250 2711
rect 26216 2677 26250 2695
rect 26216 2627 26250 2639
rect 26216 2605 26250 2627
rect 26216 2559 26250 2567
rect 26216 2533 26250 2559
rect 26312 3477 26346 3503
rect 26312 3469 26346 3477
rect 26312 3409 26346 3431
rect 26312 3397 26346 3409
rect 26312 3341 26346 3359
rect 26312 3325 26346 3341
rect 26312 3273 26346 3287
rect 26312 3253 26346 3273
rect 26312 3205 26346 3215
rect 26312 3181 26346 3205
rect 26312 3137 26346 3143
rect 26312 3109 26346 3137
rect 26312 3069 26346 3071
rect 26312 3037 26346 3069
rect 26312 2967 26346 2999
rect 26312 2965 26346 2967
rect 26312 2899 26346 2927
rect 26312 2893 26346 2899
rect 26312 2831 26346 2855
rect 26312 2821 26346 2831
rect 26312 2763 26346 2783
rect 26312 2749 26346 2763
rect 26312 2695 26346 2711
rect 26312 2677 26346 2695
rect 26312 2627 26346 2639
rect 26312 2605 26346 2627
rect 26312 2559 26346 2567
rect 26312 2533 26346 2559
rect 26408 3477 26442 3503
rect 26408 3469 26442 3477
rect 26408 3409 26442 3431
rect 26408 3397 26442 3409
rect 26408 3341 26442 3359
rect 26408 3325 26442 3341
rect 26408 3273 26442 3287
rect 26408 3253 26442 3273
rect 26408 3205 26442 3215
rect 26408 3181 26442 3205
rect 26408 3137 26442 3143
rect 26408 3109 26442 3137
rect 26408 3069 26442 3071
rect 26408 3037 26442 3069
rect 26408 2967 26442 2999
rect 26408 2965 26442 2967
rect 26408 2899 26442 2927
rect 26408 2893 26442 2899
rect 26408 2831 26442 2855
rect 26408 2821 26442 2831
rect 26408 2763 26442 2783
rect 26408 2749 26442 2763
rect 26408 2695 26442 2711
rect 26408 2677 26442 2695
rect 26408 2627 26442 2639
rect 26408 2605 26442 2627
rect 26408 2559 26442 2567
rect 26408 2533 26442 2559
rect 26504 3477 26538 3503
rect 26504 3469 26538 3477
rect 26504 3409 26538 3431
rect 26504 3397 26538 3409
rect 26504 3341 26538 3359
rect 26504 3325 26538 3341
rect 26504 3273 26538 3287
rect 26504 3253 26538 3273
rect 26504 3205 26538 3215
rect 26504 3181 26538 3205
rect 26504 3137 26538 3143
rect 26504 3109 26538 3137
rect 26504 3069 26538 3071
rect 26504 3037 26538 3069
rect 26504 2967 26538 2999
rect 26504 2965 26538 2967
rect 26504 2899 26538 2927
rect 26504 2893 26538 2899
rect 26504 2831 26538 2855
rect 26504 2821 26538 2831
rect 26504 2763 26538 2783
rect 26504 2749 26538 2763
rect 26504 2695 26538 2711
rect 26504 2677 26538 2695
rect 26504 2627 26538 2639
rect 26504 2605 26538 2627
rect 26504 2559 26538 2567
rect 26504 2533 26538 2559
rect 26732 3485 26766 3511
rect 26732 3477 26766 3485
rect 26732 3417 26766 3439
rect 26732 3405 26766 3417
rect 26732 3349 26766 3367
rect 26732 3333 26766 3349
rect 26732 3281 26766 3295
rect 26732 3261 26766 3281
rect 26732 3213 26766 3223
rect 26732 3189 26766 3213
rect 26732 3145 26766 3151
rect 26732 3117 26766 3145
rect 26732 3077 26766 3079
rect 26732 3045 26766 3077
rect 26732 2975 26766 3007
rect 26732 2973 26766 2975
rect 26732 2907 26766 2935
rect 26732 2901 26766 2907
rect 26732 2839 26766 2863
rect 26732 2829 26766 2839
rect 26732 2771 26766 2791
rect 26732 2757 26766 2771
rect 26732 2703 26766 2719
rect 26732 2685 26766 2703
rect 26732 2635 26766 2647
rect 26732 2613 26766 2635
rect 26732 2567 26766 2575
rect 26732 2541 26766 2567
rect 26828 3485 26862 3511
rect 26828 3477 26862 3485
rect 26828 3417 26862 3439
rect 26828 3405 26862 3417
rect 26828 3349 26862 3367
rect 26828 3333 26862 3349
rect 26828 3281 26862 3295
rect 26828 3261 26862 3281
rect 26828 3213 26862 3223
rect 26828 3189 26862 3213
rect 26828 3145 26862 3151
rect 26828 3117 26862 3145
rect 26828 3077 26862 3079
rect 26828 3045 26862 3077
rect 26828 2975 26862 3007
rect 26828 2973 26862 2975
rect 26828 2907 26862 2935
rect 26828 2901 26862 2907
rect 26828 2839 26862 2863
rect 26828 2829 26862 2839
rect 26828 2771 26862 2791
rect 26828 2757 26862 2771
rect 26828 2703 26862 2719
rect 26828 2685 26862 2703
rect 26828 2635 26862 2647
rect 26828 2613 26862 2635
rect 26828 2567 26862 2575
rect 26828 2541 26862 2567
rect 26924 3485 26958 3511
rect 26924 3477 26958 3485
rect 26924 3417 26958 3439
rect 26924 3405 26958 3417
rect 26924 3349 26958 3367
rect 26924 3333 26958 3349
rect 26924 3281 26958 3295
rect 26924 3261 26958 3281
rect 26924 3213 26958 3223
rect 26924 3189 26958 3213
rect 26924 3145 26958 3151
rect 26924 3117 26958 3145
rect 26924 3077 26958 3079
rect 26924 3045 26958 3077
rect 26924 2975 26958 3007
rect 26924 2973 26958 2975
rect 26924 2907 26958 2935
rect 26924 2901 26958 2907
rect 26924 2839 26958 2863
rect 26924 2829 26958 2839
rect 26924 2771 26958 2791
rect 26924 2757 26958 2771
rect 26924 2703 26958 2719
rect 26924 2685 26958 2703
rect 26924 2635 26958 2647
rect 26924 2613 26958 2635
rect 26924 2567 26958 2575
rect 26924 2541 26958 2567
rect 27020 3485 27054 3511
rect 27020 3477 27054 3485
rect 27020 3417 27054 3439
rect 27020 3405 27054 3417
rect 27020 3349 27054 3367
rect 27020 3333 27054 3349
rect 27020 3281 27054 3295
rect 27020 3261 27054 3281
rect 27020 3213 27054 3223
rect 27020 3189 27054 3213
rect 27020 3145 27054 3151
rect 27020 3117 27054 3145
rect 27020 3077 27054 3079
rect 27020 3045 27054 3077
rect 27020 2975 27054 3007
rect 27020 2973 27054 2975
rect 27020 2907 27054 2935
rect 27020 2901 27054 2907
rect 27020 2839 27054 2863
rect 27020 2829 27054 2839
rect 27020 2771 27054 2791
rect 27020 2757 27054 2771
rect 27020 2703 27054 2719
rect 27020 2685 27054 2703
rect 27020 2635 27054 2647
rect 27020 2613 27054 2635
rect 27020 2567 27054 2575
rect 27020 2541 27054 2567
rect 27116 3485 27150 3511
rect 27116 3477 27150 3485
rect 27116 3417 27150 3439
rect 27116 3405 27150 3417
rect 27116 3349 27150 3367
rect 27116 3333 27150 3349
rect 27116 3281 27150 3295
rect 27116 3261 27150 3281
rect 27116 3213 27150 3223
rect 27116 3189 27150 3213
rect 27116 3145 27150 3151
rect 27116 3117 27150 3145
rect 27116 3077 27150 3079
rect 27116 3045 27150 3077
rect 27116 2975 27150 3007
rect 27116 2973 27150 2975
rect 27116 2907 27150 2935
rect 27116 2901 27150 2907
rect 27116 2839 27150 2863
rect 27116 2829 27150 2839
rect 27116 2771 27150 2791
rect 27116 2757 27150 2771
rect 27116 2703 27150 2719
rect 27116 2685 27150 2703
rect 27116 2635 27150 2647
rect 27116 2613 27150 2635
rect 27116 2567 27150 2575
rect 27116 2541 27150 2567
rect 27212 3485 27246 3511
rect 27212 3477 27246 3485
rect 27212 3417 27246 3439
rect 27212 3405 27246 3417
rect 27212 3349 27246 3367
rect 27212 3333 27246 3349
rect 27212 3281 27246 3295
rect 27212 3261 27246 3281
rect 27212 3213 27246 3223
rect 27212 3189 27246 3213
rect 27212 3145 27246 3151
rect 27212 3117 27246 3145
rect 27212 3077 27246 3079
rect 27212 3045 27246 3077
rect 27212 2975 27246 3007
rect 27212 2973 27246 2975
rect 27212 2907 27246 2935
rect 27212 2901 27246 2907
rect 27212 2839 27246 2863
rect 27212 2829 27246 2839
rect 27212 2771 27246 2791
rect 27212 2757 27246 2771
rect 27212 2703 27246 2719
rect 27212 2685 27246 2703
rect 27212 2635 27246 2647
rect 27212 2613 27246 2635
rect 27212 2567 27246 2575
rect 27212 2541 27246 2567
rect 27308 3485 27342 3511
rect 27308 3477 27342 3485
rect 27308 3417 27342 3439
rect 27308 3405 27342 3417
rect 27308 3349 27342 3367
rect 27308 3333 27342 3349
rect 27308 3281 27342 3295
rect 27308 3261 27342 3281
rect 27308 3213 27342 3223
rect 27308 3189 27342 3213
rect 27308 3145 27342 3151
rect 27308 3117 27342 3145
rect 27308 3077 27342 3079
rect 27308 3045 27342 3077
rect 27308 2975 27342 3007
rect 27308 2973 27342 2975
rect 27308 2907 27342 2935
rect 27308 2901 27342 2907
rect 27308 2839 27342 2863
rect 27308 2829 27342 2839
rect 27308 2771 27342 2791
rect 27308 2757 27342 2771
rect 27308 2703 27342 2719
rect 27308 2685 27342 2703
rect 27308 2635 27342 2647
rect 27308 2613 27342 2635
rect 27308 2567 27342 2575
rect 27308 2541 27342 2567
rect 27404 3485 27438 3511
rect 27404 3477 27438 3485
rect 27404 3417 27438 3439
rect 27404 3405 27438 3417
rect 27404 3349 27438 3367
rect 27404 3333 27438 3349
rect 27404 3281 27438 3295
rect 27404 3261 27438 3281
rect 27404 3213 27438 3223
rect 27404 3189 27438 3213
rect 27404 3145 27438 3151
rect 27404 3117 27438 3145
rect 27404 3077 27438 3079
rect 27404 3045 27438 3077
rect 27404 2975 27438 3007
rect 27404 2973 27438 2975
rect 27404 2907 27438 2935
rect 27404 2901 27438 2907
rect 27404 2839 27438 2863
rect 27404 2829 27438 2839
rect 27404 2771 27438 2791
rect 27404 2757 27438 2771
rect 27404 2703 27438 2719
rect 27404 2685 27438 2703
rect 27404 2635 27438 2647
rect 27404 2613 27438 2635
rect 27404 2567 27438 2575
rect 27404 2541 27438 2567
rect 27500 3485 27534 3511
rect 27500 3477 27534 3485
rect 27500 3417 27534 3439
rect 27500 3405 27534 3417
rect 27500 3349 27534 3367
rect 27500 3333 27534 3349
rect 27500 3281 27534 3295
rect 27500 3261 27534 3281
rect 27500 3213 27534 3223
rect 27500 3189 27534 3213
rect 27500 3145 27534 3151
rect 27500 3117 27534 3145
rect 27500 3077 27534 3079
rect 27500 3045 27534 3077
rect 27500 2975 27534 3007
rect 27500 2973 27534 2975
rect 27500 2907 27534 2935
rect 27500 2901 27534 2907
rect 27500 2839 27534 2863
rect 27500 2829 27534 2839
rect 27500 2771 27534 2791
rect 27500 2757 27534 2771
rect 27500 2703 27534 2719
rect 27500 2685 27534 2703
rect 27500 2635 27534 2647
rect 27500 2613 27534 2635
rect 27500 2567 27534 2575
rect 27500 2541 27534 2567
rect 27596 3485 27630 3511
rect 27596 3477 27630 3485
rect 27596 3417 27630 3439
rect 27596 3405 27630 3417
rect 27596 3349 27630 3367
rect 27596 3333 27630 3349
rect 27596 3281 27630 3295
rect 27596 3261 27630 3281
rect 27596 3213 27630 3223
rect 27596 3189 27630 3213
rect 27596 3145 27630 3151
rect 27596 3117 27630 3145
rect 27596 3077 27630 3079
rect 27596 3045 27630 3077
rect 27596 2975 27630 3007
rect 27596 2973 27630 2975
rect 27596 2907 27630 2935
rect 27596 2901 27630 2907
rect 27596 2839 27630 2863
rect 27596 2829 27630 2839
rect 27596 2771 27630 2791
rect 27596 2757 27630 2771
rect 27596 2703 27630 2719
rect 27596 2685 27630 2703
rect 27596 2635 27630 2647
rect 27596 2613 27630 2635
rect 27596 2567 27630 2575
rect 27596 2541 27630 2567
rect 27692 3485 27726 3511
rect 27692 3477 27726 3485
rect 27692 3417 27726 3439
rect 27692 3405 27726 3417
rect 27692 3349 27726 3367
rect 27692 3333 27726 3349
rect 27692 3281 27726 3295
rect 27692 3261 27726 3281
rect 27692 3213 27726 3223
rect 27692 3189 27726 3213
rect 27692 3145 27726 3151
rect 27692 3117 27726 3145
rect 27692 3077 27726 3079
rect 27692 3045 27726 3077
rect 27692 2975 27726 3007
rect 27692 2973 27726 2975
rect 27692 2907 27726 2935
rect 27692 2901 27726 2907
rect 27692 2839 27726 2863
rect 27692 2829 27726 2839
rect 27692 2771 27726 2791
rect 27692 2757 27726 2771
rect 27692 2703 27726 2719
rect 27692 2685 27726 2703
rect 27692 2635 27726 2647
rect 27692 2613 27726 2635
rect 27692 2567 27726 2575
rect 27692 2541 27726 2567
rect 27788 3485 27822 3511
rect 27788 3477 27822 3485
rect 27788 3417 27822 3439
rect 27788 3405 27822 3417
rect 27788 3349 27822 3367
rect 27788 3333 27822 3349
rect 27788 3281 27822 3295
rect 27788 3261 27822 3281
rect 27788 3213 27822 3223
rect 27788 3189 27822 3213
rect 27788 3145 27822 3151
rect 27788 3117 27822 3145
rect 27788 3077 27822 3079
rect 27788 3045 27822 3077
rect 27788 2975 27822 3007
rect 27788 2973 27822 2975
rect 27788 2907 27822 2935
rect 27788 2901 27822 2907
rect 27788 2839 27822 2863
rect 27788 2829 27822 2839
rect 27788 2771 27822 2791
rect 27788 2757 27822 2771
rect 27788 2703 27822 2719
rect 27788 2685 27822 2703
rect 27788 2635 27822 2647
rect 27788 2613 27822 2635
rect 27788 2567 27822 2575
rect 27788 2541 27822 2567
rect 27884 3485 27918 3511
rect 27884 3477 27918 3485
rect 27884 3417 27918 3439
rect 27884 3405 27918 3417
rect 27884 3349 27918 3367
rect 27884 3333 27918 3349
rect 27884 3281 27918 3295
rect 27884 3261 27918 3281
rect 27884 3213 27918 3223
rect 27884 3189 27918 3213
rect 27884 3145 27918 3151
rect 27884 3117 27918 3145
rect 27884 3077 27918 3079
rect 27884 3045 27918 3077
rect 27884 2975 27918 3007
rect 27884 2973 27918 2975
rect 27884 2907 27918 2935
rect 27884 2901 27918 2907
rect 27884 2839 27918 2863
rect 27884 2829 27918 2839
rect 27884 2771 27918 2791
rect 27884 2757 27918 2771
rect 27884 2703 27918 2719
rect 27884 2685 27918 2703
rect 27884 2635 27918 2647
rect 27884 2613 27918 2635
rect 27884 2567 27918 2575
rect 27884 2541 27918 2567
rect 27980 3485 28014 3511
rect 27980 3477 28014 3485
rect 27980 3417 28014 3439
rect 27980 3405 28014 3417
rect 27980 3349 28014 3367
rect 27980 3333 28014 3349
rect 27980 3281 28014 3295
rect 27980 3261 28014 3281
rect 27980 3213 28014 3223
rect 27980 3189 28014 3213
rect 27980 3145 28014 3151
rect 27980 3117 28014 3145
rect 27980 3077 28014 3079
rect 27980 3045 28014 3077
rect 27980 2975 28014 3007
rect 27980 2973 28014 2975
rect 27980 2907 28014 2935
rect 27980 2901 28014 2907
rect 27980 2839 28014 2863
rect 27980 2829 28014 2839
rect 27980 2771 28014 2791
rect 27980 2757 28014 2771
rect 27980 2703 28014 2719
rect 27980 2685 28014 2703
rect 27980 2635 28014 2647
rect 27980 2613 28014 2635
rect 27980 2567 28014 2575
rect 27980 2541 28014 2567
rect 28076 3485 28110 3511
rect 28076 3477 28110 3485
rect 28076 3417 28110 3439
rect 28076 3405 28110 3417
rect 28076 3349 28110 3367
rect 28076 3333 28110 3349
rect 28076 3281 28110 3295
rect 28076 3261 28110 3281
rect 28076 3213 28110 3223
rect 28076 3189 28110 3213
rect 28076 3145 28110 3151
rect 28076 3117 28110 3145
rect 28076 3077 28110 3079
rect 28076 3045 28110 3077
rect 28076 2975 28110 3007
rect 28076 2973 28110 2975
rect 28076 2907 28110 2935
rect 28076 2901 28110 2907
rect 28076 2839 28110 2863
rect 28076 2829 28110 2839
rect 28076 2771 28110 2791
rect 28076 2757 28110 2771
rect 28076 2703 28110 2719
rect 28076 2685 28110 2703
rect 28076 2635 28110 2647
rect 28076 2613 28110 2635
rect 28076 2567 28110 2575
rect 28076 2541 28110 2567
rect 28172 3485 28206 3511
rect 28172 3477 28206 3485
rect 28172 3417 28206 3439
rect 28172 3405 28206 3417
rect 28172 3349 28206 3367
rect 28172 3333 28206 3349
rect 28172 3281 28206 3295
rect 28172 3261 28206 3281
rect 28172 3213 28206 3223
rect 28172 3189 28206 3213
rect 28172 3145 28206 3151
rect 28172 3117 28206 3145
rect 28172 3077 28206 3079
rect 28172 3045 28206 3077
rect 28172 2975 28206 3007
rect 28172 2973 28206 2975
rect 28172 2907 28206 2935
rect 28172 2901 28206 2907
rect 28172 2839 28206 2863
rect 28172 2829 28206 2839
rect 28172 2771 28206 2791
rect 28172 2757 28206 2771
rect 28172 2703 28206 2719
rect 28172 2685 28206 2703
rect 28172 2635 28206 2647
rect 28172 2613 28206 2635
rect 28172 2567 28206 2575
rect 28172 2541 28206 2567
rect 28268 3485 28302 3511
rect 28268 3477 28302 3485
rect 28268 3417 28302 3439
rect 28268 3405 28302 3417
rect 28268 3349 28302 3367
rect 28268 3333 28302 3349
rect 28268 3281 28302 3295
rect 28268 3261 28302 3281
rect 28268 3213 28302 3223
rect 28268 3189 28302 3213
rect 28268 3145 28302 3151
rect 28268 3117 28302 3145
rect 28268 3077 28302 3079
rect 28268 3045 28302 3077
rect 28268 2975 28302 3007
rect 28268 2973 28302 2975
rect 28268 2907 28302 2935
rect 28268 2901 28302 2907
rect 28268 2839 28302 2863
rect 28268 2829 28302 2839
rect 28268 2771 28302 2791
rect 28268 2757 28302 2771
rect 28268 2703 28302 2719
rect 28268 2685 28302 2703
rect 28268 2635 28302 2647
rect 28268 2613 28302 2635
rect 28268 2567 28302 2575
rect 28268 2541 28302 2567
rect 28364 3485 28398 3511
rect 28364 3477 28398 3485
rect 28364 3417 28398 3439
rect 28364 3405 28398 3417
rect 28364 3349 28398 3367
rect 28364 3333 28398 3349
rect 28364 3281 28398 3295
rect 28364 3261 28398 3281
rect 28364 3213 28398 3223
rect 28364 3189 28398 3213
rect 28364 3145 28398 3151
rect 28364 3117 28398 3145
rect 28364 3077 28398 3079
rect 28364 3045 28398 3077
rect 28364 2975 28398 3007
rect 28364 2973 28398 2975
rect 28364 2907 28398 2935
rect 28364 2901 28398 2907
rect 28364 2839 28398 2863
rect 28364 2829 28398 2839
rect 28364 2771 28398 2791
rect 28364 2757 28398 2771
rect 28364 2703 28398 2719
rect 28364 2685 28398 2703
rect 28364 2635 28398 2647
rect 28364 2613 28398 2635
rect 28364 2567 28398 2575
rect 28364 2541 28398 2567
rect 28460 3485 28494 3511
rect 28460 3477 28494 3485
rect 28460 3417 28494 3439
rect 28460 3405 28494 3417
rect 28460 3349 28494 3367
rect 28460 3333 28494 3349
rect 28460 3281 28494 3295
rect 28460 3261 28494 3281
rect 28460 3213 28494 3223
rect 28460 3189 28494 3213
rect 28460 3145 28494 3151
rect 28460 3117 28494 3145
rect 28460 3077 28494 3079
rect 28460 3045 28494 3077
rect 28460 2975 28494 3007
rect 28460 2973 28494 2975
rect 28460 2907 28494 2935
rect 28460 2901 28494 2907
rect 28460 2839 28494 2863
rect 28460 2829 28494 2839
rect 28460 2771 28494 2791
rect 28460 2757 28494 2771
rect 28460 2703 28494 2719
rect 28460 2685 28494 2703
rect 28460 2635 28494 2647
rect 28460 2613 28494 2635
rect 28460 2567 28494 2575
rect 28460 2541 28494 2567
rect 28556 3485 28590 3511
rect 28556 3477 28590 3485
rect 28556 3417 28590 3439
rect 28556 3405 28590 3417
rect 28556 3349 28590 3367
rect 28556 3333 28590 3349
rect 28556 3281 28590 3295
rect 28556 3261 28590 3281
rect 28556 3213 28590 3223
rect 28556 3189 28590 3213
rect 28556 3145 28590 3151
rect 28556 3117 28590 3145
rect 28556 3077 28590 3079
rect 28556 3045 28590 3077
rect 28556 2975 28590 3007
rect 28556 2973 28590 2975
rect 28556 2907 28590 2935
rect 28556 2901 28590 2907
rect 28556 2839 28590 2863
rect 28556 2829 28590 2839
rect 28556 2771 28590 2791
rect 28556 2757 28590 2771
rect 28556 2703 28590 2719
rect 28556 2685 28590 2703
rect 28556 2635 28590 2647
rect 28556 2613 28590 2635
rect 28556 2567 28590 2575
rect 28556 2541 28590 2567
rect 28652 3485 28686 3511
rect 28652 3477 28686 3485
rect 28652 3417 28686 3439
rect 28652 3405 28686 3417
rect 28652 3349 28686 3367
rect 28652 3333 28686 3349
rect 28652 3281 28686 3295
rect 28652 3261 28686 3281
rect 28652 3213 28686 3223
rect 28652 3189 28686 3213
rect 28652 3145 28686 3151
rect 28652 3117 28686 3145
rect 28652 3077 28686 3079
rect 28652 3045 28686 3077
rect 28652 2975 28686 3007
rect 28652 2973 28686 2975
rect 28652 2907 28686 2935
rect 28652 2901 28686 2907
rect 28652 2839 28686 2863
rect 28652 2829 28686 2839
rect 28652 2771 28686 2791
rect 28652 2757 28686 2771
rect 28652 2703 28686 2719
rect 28652 2685 28686 2703
rect 28652 2635 28686 2647
rect 28652 2613 28686 2635
rect 28652 2567 28686 2575
rect 28652 2541 28686 2567
rect 14096 2405 14130 2411
rect 14096 2377 14130 2405
rect 14579 2394 14613 2428
rect 14096 2337 14130 2339
rect 14096 2305 14130 2337
rect 14392 2316 14426 2350
rect 14096 2235 14130 2267
rect 14096 2233 14130 2235
rect 14096 2167 14130 2195
rect 14096 2161 14130 2167
rect 14096 2099 14130 2123
rect 14096 2089 14130 2099
rect 14096 2031 14130 2051
rect 14096 2017 14130 2031
rect 14096 1963 14130 1979
rect 14096 1945 14130 1963
rect 14096 1895 14130 1907
rect 14096 1873 14130 1895
rect 14096 1827 14130 1835
rect 14096 1801 14130 1827
rect 14500 2227 14534 2229
rect 14500 2195 14534 2227
rect 14500 2125 14534 2157
rect 14500 2123 14534 2125
rect 10652 1644 10686 1678
rect 13808 1618 13842 1652
rect 14658 2227 14692 2229
rect 14658 2195 14692 2227
rect 14658 2125 14692 2157
rect 17947 2193 18125 2299
rect 19954 2193 20132 2299
rect 21949 2196 22127 2302
rect 23302 2191 23480 2297
rect 25305 2190 25483 2296
rect 14658 2123 14692 2125
rect 734 1424 768 1458
rect -1095 1264 -1061 1298
rect -899 1264 -865 1298
rect 158 1227 192 1253
rect 158 1219 192 1227
rect -1686 1025 -1652 1051
rect -1686 1017 -1652 1025
rect -1686 957 -1652 979
rect -1686 945 -1652 957
rect -1686 889 -1652 907
rect -1686 873 -1652 889
rect -1686 821 -1652 835
rect -1686 801 -1652 821
rect -1686 753 -1652 763
rect -1686 729 -1652 753
rect -1686 685 -1652 691
rect -1686 657 -1652 685
rect -1686 617 -1652 619
rect -1686 585 -1652 617
rect -1686 515 -1652 547
rect -1686 513 -1652 515
rect -1686 447 -1652 475
rect -1686 441 -1652 447
rect -1686 379 -1652 403
rect -1686 369 -1652 379
rect -1686 311 -1652 331
rect -1686 297 -1652 311
rect -1686 243 -1652 259
rect -1686 225 -1652 243
rect -1686 175 -1652 187
rect -1686 153 -1652 175
rect -1686 107 -1652 115
rect -1686 81 -1652 107
rect -1588 1025 -1554 1051
rect -1588 1017 -1554 1025
rect -1588 957 -1554 979
rect -1588 945 -1554 957
rect -1588 889 -1554 907
rect -1588 873 -1554 889
rect -1588 821 -1554 835
rect -1588 801 -1554 821
rect -1588 753 -1554 763
rect -1588 729 -1554 753
rect -1588 685 -1554 691
rect -1588 657 -1554 685
rect -1588 617 -1554 619
rect -1588 585 -1554 617
rect -1588 515 -1554 547
rect -1588 513 -1554 515
rect -1588 447 -1554 475
rect -1588 441 -1554 447
rect -1588 379 -1554 403
rect -1588 369 -1554 379
rect -1588 311 -1554 331
rect -1588 297 -1554 311
rect -1588 243 -1554 259
rect -1588 225 -1554 243
rect -1588 175 -1554 187
rect -1588 153 -1554 175
rect -1588 107 -1554 115
rect -1588 81 -1554 107
rect -1490 1025 -1456 1051
rect -1490 1017 -1456 1025
rect -1490 957 -1456 979
rect -1490 945 -1456 957
rect -1490 889 -1456 907
rect -1490 873 -1456 889
rect -1490 821 -1456 835
rect -1490 801 -1456 821
rect -1490 753 -1456 763
rect -1490 729 -1456 753
rect -1490 685 -1456 691
rect -1490 657 -1456 685
rect -1490 617 -1456 619
rect -1490 585 -1456 617
rect -1490 515 -1456 547
rect -1490 513 -1456 515
rect -1490 447 -1456 475
rect -1490 441 -1456 447
rect -1490 379 -1456 403
rect -1490 369 -1456 379
rect -1490 311 -1456 331
rect -1490 297 -1456 311
rect -1490 243 -1456 259
rect -1490 225 -1456 243
rect -1490 175 -1456 187
rect -1490 153 -1456 175
rect -1490 107 -1456 115
rect -1490 81 -1456 107
rect -1392 1025 -1358 1051
rect -1392 1017 -1358 1025
rect -1392 957 -1358 979
rect -1392 945 -1358 957
rect -1392 889 -1358 907
rect -1392 873 -1358 889
rect -1392 821 -1358 835
rect -1392 801 -1358 821
rect -1392 753 -1358 763
rect -1392 729 -1358 753
rect -1392 685 -1358 691
rect -1392 657 -1358 685
rect -1392 617 -1358 619
rect -1392 585 -1358 617
rect -1392 515 -1358 547
rect -1392 513 -1358 515
rect -1392 447 -1358 475
rect -1392 441 -1358 447
rect -1392 379 -1358 403
rect -1392 369 -1358 379
rect -1392 311 -1358 331
rect -1392 297 -1358 311
rect -1392 243 -1358 259
rect -1392 225 -1358 243
rect -1392 175 -1358 187
rect -1392 153 -1358 175
rect -1392 107 -1358 115
rect -1392 81 -1358 107
rect -1294 1025 -1260 1051
rect -1294 1017 -1260 1025
rect -1294 957 -1260 979
rect -1294 945 -1260 957
rect -1294 889 -1260 907
rect -1294 873 -1260 889
rect -1294 821 -1260 835
rect -1294 801 -1260 821
rect -1294 753 -1260 763
rect -1294 729 -1260 753
rect -1294 685 -1260 691
rect -1294 657 -1260 685
rect -1294 617 -1260 619
rect -1294 585 -1260 617
rect -1294 515 -1260 547
rect -1294 513 -1260 515
rect -1294 447 -1260 475
rect -1294 441 -1260 447
rect -1294 379 -1260 403
rect -1294 369 -1260 379
rect -1294 311 -1260 331
rect -1294 297 -1260 311
rect -1294 243 -1260 259
rect -1294 225 -1260 243
rect -1294 175 -1260 187
rect -1294 153 -1260 175
rect -1294 107 -1260 115
rect -1294 81 -1260 107
rect -1196 1025 -1162 1051
rect -1196 1017 -1162 1025
rect -1196 957 -1162 979
rect -1196 945 -1162 957
rect -1196 889 -1162 907
rect -1196 873 -1162 889
rect -1196 821 -1162 835
rect -1196 801 -1162 821
rect -1196 753 -1162 763
rect -1196 729 -1162 753
rect -1196 685 -1162 691
rect -1196 657 -1162 685
rect -1196 617 -1162 619
rect -1196 585 -1162 617
rect -1196 515 -1162 547
rect -1196 513 -1162 515
rect -1196 447 -1162 475
rect -1196 441 -1162 447
rect -1196 379 -1162 403
rect -1196 369 -1162 379
rect -1196 311 -1162 331
rect -1196 297 -1162 311
rect -1196 243 -1162 259
rect -1196 225 -1162 243
rect -1196 175 -1162 187
rect -1196 153 -1162 175
rect -1196 107 -1162 115
rect -1196 81 -1162 107
rect -1098 1025 -1064 1051
rect -1098 1017 -1064 1025
rect -1098 957 -1064 979
rect -1098 945 -1064 957
rect -1098 889 -1064 907
rect -1098 873 -1064 889
rect -1098 821 -1064 835
rect -1098 801 -1064 821
rect -1098 753 -1064 763
rect -1098 729 -1064 753
rect -1098 685 -1064 691
rect -1098 657 -1064 685
rect -1098 617 -1064 619
rect -1098 585 -1064 617
rect -1098 515 -1064 547
rect -1098 513 -1064 515
rect -1098 447 -1064 475
rect -1098 441 -1064 447
rect -1098 379 -1064 403
rect -1098 369 -1064 379
rect -1098 311 -1064 331
rect -1098 297 -1064 311
rect -1098 243 -1064 259
rect -1098 225 -1064 243
rect -1098 175 -1064 187
rect -1098 153 -1064 175
rect -1098 107 -1064 115
rect -1098 81 -1064 107
rect 158 1159 192 1181
rect 158 1147 192 1159
rect 158 1091 192 1109
rect 158 1075 192 1091
rect -1000 1025 -966 1051
rect -1000 1017 -966 1025
rect -1000 957 -966 979
rect -1000 945 -966 957
rect -1000 889 -966 907
rect -1000 873 -966 889
rect -1000 821 -966 835
rect -1000 801 -966 821
rect -1000 753 -966 763
rect -1000 729 -966 753
rect -1000 685 -966 691
rect -1000 657 -966 685
rect -1000 617 -966 619
rect -1000 585 -966 617
rect -1000 515 -966 547
rect -1000 513 -966 515
rect -1000 447 -966 475
rect -1000 441 -966 447
rect -1000 379 -966 403
rect -1000 369 -966 379
rect -1000 311 -966 331
rect -1000 297 -966 311
rect -1000 243 -966 259
rect -1000 225 -966 243
rect -1000 175 -966 187
rect -1000 153 -966 175
rect -1000 107 -966 115
rect -1000 81 -966 107
rect -902 1025 -868 1051
rect -902 1017 -868 1025
rect -902 957 -868 979
rect -902 945 -868 957
rect -902 889 -868 907
rect -902 873 -868 889
rect -902 821 -868 835
rect -902 801 -868 821
rect -902 753 -868 763
rect -902 729 -868 753
rect -902 685 -868 691
rect -902 657 -868 685
rect -902 617 -868 619
rect -902 585 -868 617
rect -902 515 -868 547
rect -902 513 -868 515
rect -902 447 -868 475
rect -902 441 -868 447
rect -902 379 -868 403
rect -902 369 -868 379
rect -902 311 -868 331
rect -902 297 -868 311
rect -902 243 -868 259
rect -902 225 -868 243
rect -902 175 -868 187
rect 158 1023 192 1037
rect 158 1003 192 1023
rect 158 955 192 965
rect 158 931 192 955
rect 158 887 192 893
rect 158 859 192 887
rect 158 819 192 821
rect 158 787 192 819
rect 158 717 192 749
rect 158 715 192 717
rect 158 649 192 677
rect 158 643 192 649
rect 158 581 192 605
rect 158 571 192 581
rect 158 513 192 533
rect 158 499 192 513
rect 158 445 192 461
rect 158 427 192 445
rect 158 377 192 389
rect 158 355 192 377
rect 158 309 192 317
rect 158 283 192 309
rect 254 1227 288 1253
rect 254 1219 288 1227
rect 254 1159 288 1181
rect 254 1147 288 1159
rect 254 1091 288 1109
rect 254 1075 288 1091
rect 254 1023 288 1037
rect 254 1003 288 1023
rect 254 955 288 965
rect 254 931 288 955
rect 254 887 288 893
rect 254 859 288 887
rect 254 819 288 821
rect 254 787 288 819
rect 254 717 288 749
rect 254 715 288 717
rect 254 649 288 677
rect 254 643 288 649
rect 254 581 288 605
rect 254 571 288 581
rect 254 513 288 533
rect 254 499 288 513
rect 254 445 288 461
rect 254 427 288 445
rect 254 377 288 389
rect 254 355 288 377
rect 254 309 288 317
rect 254 283 288 309
rect 350 1227 384 1253
rect 350 1219 384 1227
rect 350 1159 384 1181
rect 350 1147 384 1159
rect 350 1091 384 1109
rect 350 1075 384 1091
rect 350 1023 384 1037
rect 350 1003 384 1023
rect 350 955 384 965
rect 350 931 384 955
rect 350 887 384 893
rect 350 859 384 887
rect 350 819 384 821
rect 350 787 384 819
rect 350 717 384 749
rect 350 715 384 717
rect 350 649 384 677
rect 350 643 384 649
rect 350 581 384 605
rect 350 571 384 581
rect 350 513 384 533
rect 350 499 384 513
rect 350 445 384 461
rect 350 427 384 445
rect 350 377 384 389
rect 350 355 384 377
rect 350 309 384 317
rect 350 283 384 309
rect 446 1227 480 1253
rect 446 1219 480 1227
rect 446 1159 480 1181
rect 446 1147 480 1159
rect 446 1091 480 1109
rect 446 1075 480 1091
rect 446 1023 480 1037
rect 446 1003 480 1023
rect 446 955 480 965
rect 446 931 480 955
rect 446 887 480 893
rect 446 859 480 887
rect 446 819 480 821
rect 446 787 480 819
rect 446 717 480 749
rect 446 715 480 717
rect 446 649 480 677
rect 446 643 480 649
rect 446 581 480 605
rect 446 571 480 581
rect 446 513 480 533
rect 446 499 480 513
rect 446 445 480 461
rect 446 427 480 445
rect 446 377 480 389
rect 446 355 480 377
rect 446 309 480 317
rect 446 283 480 309
rect 542 1227 576 1253
rect 542 1219 576 1227
rect 542 1159 576 1181
rect 542 1147 576 1159
rect 542 1091 576 1109
rect 542 1075 576 1091
rect 542 1023 576 1037
rect 542 1003 576 1023
rect 542 955 576 965
rect 542 931 576 955
rect 542 887 576 893
rect 542 859 576 887
rect 542 819 576 821
rect 542 787 576 819
rect 542 717 576 749
rect 542 715 576 717
rect 542 649 576 677
rect 542 643 576 649
rect 542 581 576 605
rect 542 571 576 581
rect 542 513 576 533
rect 542 499 576 513
rect 542 445 576 461
rect 542 427 576 445
rect 542 377 576 389
rect 542 355 576 377
rect 542 309 576 317
rect 542 283 576 309
rect 638 1227 672 1253
rect 638 1219 672 1227
rect 638 1159 672 1181
rect 638 1147 672 1159
rect 638 1091 672 1109
rect 638 1075 672 1091
rect 638 1023 672 1037
rect 638 1003 672 1023
rect 638 955 672 965
rect 638 931 672 955
rect 638 887 672 893
rect 638 859 672 887
rect 638 819 672 821
rect 638 787 672 819
rect 638 717 672 749
rect 638 715 672 717
rect 638 649 672 677
rect 638 643 672 649
rect 638 581 672 605
rect 638 571 672 581
rect 638 513 672 533
rect 638 499 672 513
rect 638 445 672 461
rect 638 427 672 445
rect 638 377 672 389
rect 638 355 672 377
rect 638 309 672 317
rect 638 283 672 309
rect 734 1227 768 1253
rect 734 1219 768 1227
rect 734 1159 768 1181
rect 734 1147 768 1159
rect 734 1091 768 1109
rect 734 1075 768 1091
rect 734 1023 768 1037
rect 734 1003 768 1023
rect 734 955 768 965
rect 734 931 768 955
rect 734 887 768 893
rect 734 859 768 887
rect 734 819 768 821
rect 734 787 768 819
rect 734 717 768 749
rect 734 715 768 717
rect 734 649 768 677
rect 734 643 768 649
rect 734 581 768 605
rect 734 571 768 581
rect 734 513 768 533
rect 734 499 768 513
rect 734 445 768 461
rect 734 427 768 445
rect 734 377 768 389
rect 734 355 768 377
rect 734 309 768 317
rect 734 283 768 309
rect 830 1227 864 1253
rect 830 1219 864 1227
rect 830 1159 864 1181
rect 830 1147 864 1159
rect 830 1091 864 1109
rect 830 1075 864 1091
rect 830 1023 864 1037
rect 830 1003 864 1023
rect 830 955 864 965
rect 830 931 864 955
rect 830 887 864 893
rect 830 859 864 887
rect 830 819 864 821
rect 830 787 864 819
rect 830 717 864 749
rect 830 715 864 717
rect 830 649 864 677
rect 830 643 864 649
rect 830 581 864 605
rect 830 571 864 581
rect 830 513 864 533
rect 830 499 864 513
rect 830 445 864 461
rect 830 427 864 445
rect 830 377 864 389
rect 830 355 864 377
rect 830 309 864 317
rect 830 283 864 309
rect 926 1227 960 1253
rect 926 1219 960 1227
rect 926 1159 960 1181
rect 926 1147 960 1159
rect 926 1091 960 1109
rect 926 1075 960 1091
rect 926 1023 960 1037
rect 926 1003 960 1023
rect 926 955 960 965
rect 926 931 960 955
rect 926 887 960 893
rect 926 859 960 887
rect 926 819 960 821
rect 926 787 960 819
rect 926 717 960 749
rect 926 715 960 717
rect 926 649 960 677
rect 926 643 960 649
rect 926 581 960 605
rect 926 571 960 581
rect 926 513 960 533
rect 926 499 960 513
rect 926 445 960 461
rect 926 427 960 445
rect 926 377 960 389
rect 926 355 960 377
rect 926 309 960 317
rect 926 283 960 309
rect 1022 1227 1056 1253
rect 1022 1219 1056 1227
rect 1022 1159 1056 1181
rect 1022 1147 1056 1159
rect 1022 1091 1056 1109
rect 1022 1075 1056 1091
rect 1022 1023 1056 1037
rect 1022 1003 1056 1023
rect 1022 955 1056 965
rect 1022 931 1056 955
rect 1022 887 1056 893
rect 1022 859 1056 887
rect 1022 819 1056 821
rect 1022 787 1056 819
rect 1022 717 1056 749
rect 1022 715 1056 717
rect 1022 649 1056 677
rect 1022 643 1056 649
rect 1022 581 1056 605
rect 1022 571 1056 581
rect 1022 513 1056 533
rect 1022 499 1056 513
rect 1022 445 1056 461
rect 1022 427 1056 445
rect 1022 377 1056 389
rect 1022 355 1056 377
rect 1022 309 1056 317
rect 1022 283 1056 309
rect 1118 1227 1152 1253
rect 1118 1219 1152 1227
rect 1118 1159 1152 1181
rect 1118 1147 1152 1159
rect 1118 1091 1152 1109
rect 1118 1075 1152 1091
rect 1118 1023 1152 1037
rect 1118 1003 1152 1023
rect 1118 955 1152 965
rect 1118 931 1152 955
rect 1118 887 1152 893
rect 1118 859 1152 887
rect 1118 819 1152 821
rect 1118 787 1152 819
rect 1118 717 1152 749
rect 1118 715 1152 717
rect 1118 649 1152 677
rect 1118 643 1152 649
rect 1118 581 1152 605
rect 1118 571 1152 581
rect 1118 513 1152 533
rect 1118 499 1152 513
rect 1118 445 1152 461
rect 1118 427 1152 445
rect 1118 377 1152 389
rect 1118 355 1152 377
rect 1118 309 1152 317
rect 1118 283 1152 309
rect 1214 1227 1248 1253
rect 1214 1219 1248 1227
rect 1214 1159 1248 1181
rect 1214 1147 1248 1159
rect 1214 1091 1248 1109
rect 1214 1075 1248 1091
rect 1214 1023 1248 1037
rect 1214 1003 1248 1023
rect 1214 955 1248 965
rect 1214 931 1248 955
rect 1214 887 1248 893
rect 1214 859 1248 887
rect 1214 819 1248 821
rect 1214 787 1248 819
rect 1214 717 1248 749
rect 1214 715 1248 717
rect 1214 649 1248 677
rect 1214 643 1248 649
rect 1214 581 1248 605
rect 1214 571 1248 581
rect 1214 513 1248 533
rect 1214 499 1248 513
rect 1214 445 1248 461
rect 1214 427 1248 445
rect 1214 377 1248 389
rect 1214 355 1248 377
rect 1214 309 1248 317
rect 1214 283 1248 309
rect 1310 1227 1344 1253
rect 1310 1219 1344 1227
rect 1310 1159 1344 1181
rect 1310 1147 1344 1159
rect 1310 1091 1344 1109
rect 1310 1075 1344 1091
rect 1310 1023 1344 1037
rect 1310 1003 1344 1023
rect 1310 955 1344 965
rect 1310 931 1344 955
rect 1310 887 1344 893
rect 1310 859 1344 887
rect 1310 819 1344 821
rect 1310 787 1344 819
rect 1310 717 1344 749
rect 1310 715 1344 717
rect 1310 649 1344 677
rect 1310 643 1344 649
rect 1310 581 1344 605
rect 1310 571 1344 581
rect 1310 513 1344 533
rect 1310 499 1344 513
rect 1310 445 1344 461
rect 1310 427 1344 445
rect 1310 377 1344 389
rect 1310 355 1344 377
rect 1310 309 1344 317
rect 1310 283 1344 309
rect -902 153 -868 175
rect -902 107 -868 115
rect -902 81 -868 107
rect 156 96 190 130
rect 830 86 864 120
rect 2400 1418 2434 1452
rect 3690 1408 3724 1442
rect 1926 1227 1960 1253
rect 1926 1219 1960 1227
rect 1926 1159 1960 1181
rect 1926 1147 1960 1159
rect 1926 1091 1960 1109
rect 1926 1075 1960 1091
rect 1926 1023 1960 1037
rect 1926 1003 1960 1023
rect 1926 955 1960 965
rect 1926 931 1960 955
rect 1926 887 1960 893
rect 1926 859 1960 887
rect 1926 819 1960 821
rect 1926 787 1960 819
rect 1926 717 1960 749
rect 1926 715 1960 717
rect 1926 649 1960 677
rect 1926 643 1960 649
rect 1926 581 1960 605
rect 1926 571 1960 581
rect 1926 513 1960 533
rect 1926 499 1960 513
rect 1926 445 1960 461
rect 1926 427 1960 445
rect 1926 377 1960 389
rect 1926 355 1960 377
rect 1926 309 1960 317
rect 1926 283 1960 309
rect 2022 1227 2056 1253
rect 2022 1219 2056 1227
rect 2022 1159 2056 1181
rect 2022 1147 2056 1159
rect 2022 1091 2056 1109
rect 2022 1075 2056 1091
rect 2022 1023 2056 1037
rect 2022 1003 2056 1023
rect 2022 955 2056 965
rect 2022 931 2056 955
rect 2022 887 2056 893
rect 2022 859 2056 887
rect 2022 819 2056 821
rect 2022 787 2056 819
rect 2022 717 2056 749
rect 2022 715 2056 717
rect 2022 649 2056 677
rect 2022 643 2056 649
rect 2022 581 2056 605
rect 2022 571 2056 581
rect 2022 513 2056 533
rect 2022 499 2056 513
rect 2022 445 2056 461
rect 2022 427 2056 445
rect 2022 377 2056 389
rect 2022 355 2056 377
rect 2022 309 2056 317
rect 2022 283 2056 309
rect 2118 1227 2152 1253
rect 2118 1219 2152 1227
rect 2118 1159 2152 1181
rect 2118 1147 2152 1159
rect 2118 1091 2152 1109
rect 2118 1075 2152 1091
rect 2118 1023 2152 1037
rect 2118 1003 2152 1023
rect 2118 955 2152 965
rect 2118 931 2152 955
rect 2118 887 2152 893
rect 2118 859 2152 887
rect 2118 819 2152 821
rect 2118 787 2152 819
rect 2118 717 2152 749
rect 2118 715 2152 717
rect 2118 649 2152 677
rect 2118 643 2152 649
rect 2118 581 2152 605
rect 2118 571 2152 581
rect 2118 513 2152 533
rect 2118 499 2152 513
rect 2118 445 2152 461
rect 2118 427 2152 445
rect 2118 377 2152 389
rect 2118 355 2152 377
rect 2118 309 2152 317
rect 2118 283 2152 309
rect 2214 1227 2248 1253
rect 2214 1219 2248 1227
rect 2214 1159 2248 1181
rect 2214 1147 2248 1159
rect 2214 1091 2248 1109
rect 2214 1075 2248 1091
rect 2214 1023 2248 1037
rect 2214 1003 2248 1023
rect 2214 955 2248 965
rect 2214 931 2248 955
rect 2214 887 2248 893
rect 2214 859 2248 887
rect 2214 819 2248 821
rect 2214 787 2248 819
rect 2214 717 2248 749
rect 2214 715 2248 717
rect 2214 649 2248 677
rect 2214 643 2248 649
rect 2214 581 2248 605
rect 2214 571 2248 581
rect 2214 513 2248 533
rect 2214 499 2248 513
rect 2214 445 2248 461
rect 2214 427 2248 445
rect 2214 377 2248 389
rect 2214 355 2248 377
rect 2214 309 2248 317
rect 2214 283 2248 309
rect 2310 1227 2344 1253
rect 2310 1219 2344 1227
rect 2310 1159 2344 1181
rect 2310 1147 2344 1159
rect 2310 1091 2344 1109
rect 2310 1075 2344 1091
rect 2310 1023 2344 1037
rect 2310 1003 2344 1023
rect 2310 955 2344 965
rect 2310 931 2344 955
rect 2310 887 2344 893
rect 2310 859 2344 887
rect 2310 819 2344 821
rect 2310 787 2344 819
rect 2310 717 2344 749
rect 2310 715 2344 717
rect 2310 649 2344 677
rect 2310 643 2344 649
rect 2310 581 2344 605
rect 2310 571 2344 581
rect 2310 513 2344 533
rect 2310 499 2344 513
rect 2310 445 2344 461
rect 2310 427 2344 445
rect 2310 377 2344 389
rect 2310 355 2344 377
rect 2310 309 2344 317
rect 2310 283 2344 309
rect 2406 1227 2440 1253
rect 2406 1219 2440 1227
rect 2406 1159 2440 1181
rect 2406 1147 2440 1159
rect 2406 1091 2440 1109
rect 2406 1075 2440 1091
rect 2406 1023 2440 1037
rect 2406 1003 2440 1023
rect 2406 955 2440 965
rect 2406 931 2440 955
rect 2406 887 2440 893
rect 2406 859 2440 887
rect 2406 819 2440 821
rect 2406 787 2440 819
rect 2406 717 2440 749
rect 2406 715 2440 717
rect 2406 649 2440 677
rect 2406 643 2440 649
rect 2406 581 2440 605
rect 2406 571 2440 581
rect 2406 513 2440 533
rect 2406 499 2440 513
rect 2406 445 2440 461
rect 2406 427 2440 445
rect 2406 377 2440 389
rect 2406 355 2440 377
rect 2406 309 2440 317
rect 2406 283 2440 309
rect 2502 1227 2536 1253
rect 2502 1219 2536 1227
rect 2502 1159 2536 1181
rect 2502 1147 2536 1159
rect 2502 1091 2536 1109
rect 2502 1075 2536 1091
rect 2502 1023 2536 1037
rect 2502 1003 2536 1023
rect 2502 955 2536 965
rect 2502 931 2536 955
rect 2502 887 2536 893
rect 2502 859 2536 887
rect 2502 819 2536 821
rect 2502 787 2536 819
rect 2502 717 2536 749
rect 2502 715 2536 717
rect 2502 649 2536 677
rect 2502 643 2536 649
rect 2502 581 2536 605
rect 2502 571 2536 581
rect 2502 513 2536 533
rect 2502 499 2536 513
rect 2502 445 2536 461
rect 2502 427 2536 445
rect 2502 377 2536 389
rect 2502 355 2536 377
rect 2502 309 2536 317
rect 2502 283 2536 309
rect 2598 1227 2632 1253
rect 2598 1219 2632 1227
rect 2598 1159 2632 1181
rect 2598 1147 2632 1159
rect 2598 1091 2632 1109
rect 2598 1075 2632 1091
rect 2598 1023 2632 1037
rect 2598 1003 2632 1023
rect 2598 955 2632 965
rect 2598 931 2632 955
rect 2598 887 2632 893
rect 2598 859 2632 887
rect 2598 819 2632 821
rect 2598 787 2632 819
rect 2598 717 2632 749
rect 2598 715 2632 717
rect 2598 649 2632 677
rect 2598 643 2632 649
rect 2598 581 2632 605
rect 2598 571 2632 581
rect 2598 513 2632 533
rect 2598 499 2632 513
rect 2598 445 2632 461
rect 2598 427 2632 445
rect 2598 377 2632 389
rect 2598 355 2632 377
rect 2598 309 2632 317
rect 2598 283 2632 309
rect 2694 1227 2728 1253
rect 2694 1219 2728 1227
rect 2694 1159 2728 1181
rect 2694 1147 2728 1159
rect 2694 1091 2728 1109
rect 2694 1075 2728 1091
rect 2694 1023 2728 1037
rect 2694 1003 2728 1023
rect 2694 955 2728 965
rect 2694 931 2728 955
rect 2694 887 2728 893
rect 2694 859 2728 887
rect 2694 819 2728 821
rect 2694 787 2728 819
rect 2694 717 2728 749
rect 2694 715 2728 717
rect 2694 649 2728 677
rect 2694 643 2728 649
rect 2694 581 2728 605
rect 2694 571 2728 581
rect 2694 513 2728 533
rect 2694 499 2728 513
rect 2694 445 2728 461
rect 2694 427 2728 445
rect 2694 377 2728 389
rect 2694 355 2728 377
rect 2694 309 2728 317
rect 2694 283 2728 309
rect 2790 1227 2824 1253
rect 2790 1219 2824 1227
rect 2790 1159 2824 1181
rect 2790 1147 2824 1159
rect 2790 1091 2824 1109
rect 2790 1075 2824 1091
rect 2790 1023 2824 1037
rect 2790 1003 2824 1023
rect 2790 955 2824 965
rect 2790 931 2824 955
rect 2790 887 2824 893
rect 2790 859 2824 887
rect 2790 819 2824 821
rect 2790 787 2824 819
rect 2790 717 2824 749
rect 2790 715 2824 717
rect 2790 649 2824 677
rect 2790 643 2824 649
rect 2790 581 2824 605
rect 2790 571 2824 581
rect 2790 513 2824 533
rect 2790 499 2824 513
rect 2790 445 2824 461
rect 2790 427 2824 445
rect 2790 377 2824 389
rect 2790 355 2824 377
rect 2790 309 2824 317
rect 2790 283 2824 309
rect 2886 1227 2920 1253
rect 2886 1219 2920 1227
rect 2886 1159 2920 1181
rect 2886 1147 2920 1159
rect 2886 1091 2920 1109
rect 2886 1075 2920 1091
rect 2886 1023 2920 1037
rect 2886 1003 2920 1023
rect 2886 955 2920 965
rect 2886 931 2920 955
rect 2886 887 2920 893
rect 2886 859 2920 887
rect 2886 819 2920 821
rect 2886 787 2920 819
rect 2886 717 2920 749
rect 2886 715 2920 717
rect 2886 649 2920 677
rect 2886 643 2920 649
rect 2886 581 2920 605
rect 2886 571 2920 581
rect 2886 513 2920 533
rect 2886 499 2920 513
rect 2886 445 2920 461
rect 2886 427 2920 445
rect 2886 377 2920 389
rect 2886 355 2920 377
rect 2886 309 2920 317
rect 2886 283 2920 309
rect 2982 1227 3016 1253
rect 2982 1219 3016 1227
rect 2982 1159 3016 1181
rect 2982 1147 3016 1159
rect 2982 1091 3016 1109
rect 2982 1075 3016 1091
rect 2982 1023 3016 1037
rect 2982 1003 3016 1023
rect 2982 955 3016 965
rect 2982 931 3016 955
rect 2982 887 3016 893
rect 2982 859 3016 887
rect 2982 819 3016 821
rect 2982 787 3016 819
rect 2982 717 3016 749
rect 2982 715 3016 717
rect 2982 649 3016 677
rect 2982 643 3016 649
rect 2982 581 3016 605
rect 2982 571 3016 581
rect 2982 513 3016 533
rect 2982 499 3016 513
rect 2982 445 3016 461
rect 2982 427 3016 445
rect 2982 377 3016 389
rect 2982 355 3016 377
rect 2982 309 3016 317
rect 2982 283 3016 309
rect 3114 1211 3148 1237
rect 3114 1203 3148 1211
rect 3114 1143 3148 1165
rect 3114 1131 3148 1143
rect 3114 1075 3148 1093
rect 3114 1059 3148 1075
rect 3114 1007 3148 1021
rect 3114 987 3148 1007
rect 3114 939 3148 949
rect 3114 915 3148 939
rect 3114 871 3148 877
rect 3114 843 3148 871
rect 3114 803 3148 805
rect 3114 771 3148 803
rect 3114 701 3148 733
rect 3114 699 3148 701
rect 3114 633 3148 661
rect 3114 627 3148 633
rect 3114 565 3148 589
rect 3114 555 3148 565
rect 3114 497 3148 517
rect 3114 483 3148 497
rect 3114 429 3148 445
rect 3114 411 3148 429
rect 3114 361 3148 373
rect 3114 339 3148 361
rect 3114 293 3148 301
rect 3114 267 3148 293
rect 3210 1211 3244 1237
rect 3210 1203 3244 1211
rect 3210 1143 3244 1165
rect 3210 1131 3244 1143
rect 3210 1075 3244 1093
rect 3210 1059 3244 1075
rect 3210 1007 3244 1021
rect 3210 987 3244 1007
rect 3210 939 3244 949
rect 3210 915 3244 939
rect 3210 871 3244 877
rect 3210 843 3244 871
rect 3210 803 3244 805
rect 3210 771 3244 803
rect 3210 701 3244 733
rect 3210 699 3244 701
rect 3210 633 3244 661
rect 3210 627 3244 633
rect 3210 565 3244 589
rect 3210 555 3244 565
rect 3210 497 3244 517
rect 3210 483 3244 497
rect 3210 429 3244 445
rect 3210 411 3244 429
rect 3210 361 3244 373
rect 3210 339 3244 361
rect 3210 293 3244 301
rect 3210 267 3244 293
rect 3306 1211 3340 1237
rect 3306 1203 3340 1211
rect 3306 1143 3340 1165
rect 3306 1131 3340 1143
rect 3306 1075 3340 1093
rect 3306 1059 3340 1075
rect 3306 1007 3340 1021
rect 3306 987 3340 1007
rect 3306 939 3340 949
rect 3306 915 3340 939
rect 3306 871 3340 877
rect 3306 843 3340 871
rect 3306 803 3340 805
rect 3306 771 3340 803
rect 3306 701 3340 733
rect 3306 699 3340 701
rect 3306 633 3340 661
rect 3306 627 3340 633
rect 3306 565 3340 589
rect 3306 555 3340 565
rect 3306 497 3340 517
rect 3306 483 3340 497
rect 3306 429 3340 445
rect 3306 411 3340 429
rect 3306 361 3340 373
rect 3306 339 3340 361
rect 3306 293 3340 301
rect 3306 267 3340 293
rect 3402 1211 3436 1237
rect 3402 1203 3436 1211
rect 3402 1143 3436 1165
rect 3402 1131 3436 1143
rect 3402 1075 3436 1093
rect 3402 1059 3436 1075
rect 3402 1007 3436 1021
rect 3402 987 3436 1007
rect 3402 939 3436 949
rect 3402 915 3436 939
rect 3402 871 3436 877
rect 3402 843 3436 871
rect 3402 803 3436 805
rect 3402 771 3436 803
rect 3402 701 3436 733
rect 3402 699 3436 701
rect 3402 633 3436 661
rect 3402 627 3436 633
rect 3402 565 3436 589
rect 3402 555 3436 565
rect 3402 497 3436 517
rect 3402 483 3436 497
rect 3402 429 3436 445
rect 3402 411 3436 429
rect 3402 361 3436 373
rect 3402 339 3436 361
rect 3402 293 3436 301
rect 3402 267 3436 293
rect 3498 1211 3532 1237
rect 3498 1203 3532 1211
rect 3498 1143 3532 1165
rect 3498 1131 3532 1143
rect 3498 1075 3532 1093
rect 3498 1059 3532 1075
rect 3498 1007 3532 1021
rect 3498 987 3532 1007
rect 3498 939 3532 949
rect 3498 915 3532 939
rect 3498 871 3532 877
rect 3498 843 3532 871
rect 3498 803 3532 805
rect 3498 771 3532 803
rect 3498 701 3532 733
rect 3498 699 3532 701
rect 3498 633 3532 661
rect 3498 627 3532 633
rect 3498 565 3532 589
rect 3498 555 3532 565
rect 3498 497 3532 517
rect 3498 483 3532 497
rect 3498 429 3532 445
rect 3498 411 3532 429
rect 3498 361 3532 373
rect 3498 339 3532 361
rect 3498 293 3532 301
rect 3498 267 3532 293
rect 3594 1211 3628 1237
rect 3594 1203 3628 1211
rect 3594 1143 3628 1165
rect 3594 1131 3628 1143
rect 3594 1075 3628 1093
rect 3594 1059 3628 1075
rect 3594 1007 3628 1021
rect 3594 987 3628 1007
rect 3594 939 3628 949
rect 3594 915 3628 939
rect 3594 871 3628 877
rect 3594 843 3628 871
rect 3594 803 3628 805
rect 3594 771 3628 803
rect 3594 701 3628 733
rect 3594 699 3628 701
rect 3594 633 3628 661
rect 3594 627 3628 633
rect 3594 565 3628 589
rect 3594 555 3628 565
rect 3594 497 3628 517
rect 3594 483 3628 497
rect 3594 429 3628 445
rect 3594 411 3628 429
rect 3594 361 3628 373
rect 3594 339 3628 361
rect 3594 293 3628 301
rect 3594 267 3628 293
rect 3690 1211 3724 1237
rect 3690 1203 3724 1211
rect 3690 1143 3724 1165
rect 3690 1131 3724 1143
rect 3690 1075 3724 1093
rect 3690 1059 3724 1075
rect 3690 1007 3724 1021
rect 3690 987 3724 1007
rect 3690 939 3724 949
rect 3690 915 3724 939
rect 3690 871 3724 877
rect 3690 843 3724 871
rect 3690 803 3724 805
rect 3690 771 3724 803
rect 3690 701 3724 733
rect 3690 699 3724 701
rect 3690 633 3724 661
rect 3690 627 3724 633
rect 3690 565 3724 589
rect 3690 555 3724 565
rect 3690 497 3724 517
rect 3690 483 3724 497
rect 3690 429 3724 445
rect 3690 411 3724 429
rect 3690 361 3724 373
rect 3690 339 3724 361
rect 3690 293 3724 301
rect 3690 267 3724 293
rect 3786 1211 3820 1237
rect 3786 1203 3820 1211
rect 3786 1143 3820 1165
rect 3786 1131 3820 1143
rect 3786 1075 3820 1093
rect 3786 1059 3820 1075
rect 3786 1007 3820 1021
rect 3786 987 3820 1007
rect 3786 939 3820 949
rect 3786 915 3820 939
rect 3786 871 3820 877
rect 3786 843 3820 871
rect 3786 803 3820 805
rect 3786 771 3820 803
rect 3786 701 3820 733
rect 3786 699 3820 701
rect 3786 633 3820 661
rect 3786 627 3820 633
rect 3786 565 3820 589
rect 3786 555 3820 565
rect 3786 497 3820 517
rect 3786 483 3820 497
rect 3786 429 3820 445
rect 3786 411 3820 429
rect 3786 361 3820 373
rect 3786 339 3820 361
rect 3786 293 3820 301
rect 3786 267 3820 293
rect 3882 1211 3916 1237
rect 3882 1203 3916 1211
rect 3882 1143 3916 1165
rect 3882 1131 3916 1143
rect 3882 1075 3916 1093
rect 3882 1059 3916 1075
rect 3882 1007 3916 1021
rect 3882 987 3916 1007
rect 3882 939 3916 949
rect 3882 915 3916 939
rect 3882 871 3916 877
rect 3882 843 3916 871
rect 3882 803 3916 805
rect 3882 771 3916 803
rect 3882 701 3916 733
rect 3882 699 3916 701
rect 3882 633 3916 661
rect 3882 627 3916 633
rect 3882 565 3916 589
rect 3882 555 3916 565
rect 3882 497 3916 517
rect 3882 483 3916 497
rect 3882 429 3916 445
rect 3882 411 3916 429
rect 3882 361 3916 373
rect 3882 339 3916 361
rect 3882 293 3916 301
rect 3882 267 3916 293
rect 3978 1211 4012 1237
rect 3978 1203 4012 1211
rect 3978 1143 4012 1165
rect 3978 1131 4012 1143
rect 3978 1075 4012 1093
rect 3978 1059 4012 1075
rect 3978 1007 4012 1021
rect 3978 987 4012 1007
rect 3978 939 4012 949
rect 3978 915 4012 939
rect 3978 871 4012 877
rect 3978 843 4012 871
rect 3978 803 4012 805
rect 3978 771 4012 803
rect 3978 701 4012 733
rect 3978 699 4012 701
rect 3978 633 4012 661
rect 3978 627 4012 633
rect 3978 565 4012 589
rect 3978 555 4012 565
rect 3978 497 4012 517
rect 3978 483 4012 497
rect 3978 429 4012 445
rect 3978 411 4012 429
rect 3978 361 4012 373
rect 3978 339 4012 361
rect 3978 293 4012 301
rect 3978 267 4012 293
rect 4074 1211 4108 1237
rect 4074 1203 4108 1211
rect 4074 1143 4108 1165
rect 4074 1131 4108 1143
rect 4074 1075 4108 1093
rect 4074 1059 4108 1075
rect 4074 1007 4108 1021
rect 4074 987 4108 1007
rect 4074 939 4108 949
rect 4074 915 4108 939
rect 4074 871 4108 877
rect 4074 843 4108 871
rect 4074 803 4108 805
rect 4074 771 4108 803
rect 4074 701 4108 733
rect 4074 699 4108 701
rect 4074 633 4108 661
rect 4074 627 4108 633
rect 4074 565 4108 589
rect 4074 555 4108 565
rect 4074 497 4108 517
rect 4074 483 4108 497
rect 4074 429 4108 445
rect 4074 411 4108 429
rect 4074 361 4108 373
rect 4074 339 4108 361
rect 4074 293 4108 301
rect 4074 267 4108 293
rect 4170 1211 4204 1237
rect 4170 1203 4204 1211
rect 4170 1143 4204 1165
rect 4170 1131 4204 1143
rect 4170 1075 4204 1093
rect 4170 1059 4204 1075
rect 4170 1007 4204 1021
rect 4170 987 4204 1007
rect 4170 939 4204 949
rect 4170 915 4204 939
rect 4170 871 4204 877
rect 4170 843 4204 871
rect 4170 803 4204 805
rect 4170 771 4204 803
rect 4170 701 4204 733
rect 4170 699 4204 701
rect 4170 633 4204 661
rect 4170 627 4204 633
rect 4170 565 4204 589
rect 4170 555 4204 565
rect 4170 497 4204 517
rect 4170 483 4204 497
rect 4170 429 4204 445
rect 4170 411 4204 429
rect 4170 361 4204 373
rect 4170 339 4204 361
rect 4170 293 4204 301
rect 4170 267 4204 293
rect 4266 1211 4300 1237
rect 4266 1203 4300 1211
rect 4266 1143 4300 1165
rect 4266 1131 4300 1143
rect 4266 1075 4300 1093
rect 4266 1059 4300 1075
rect 4266 1007 4300 1021
rect 4266 987 4300 1007
rect 4266 939 4300 949
rect 4266 915 4300 939
rect 4266 871 4300 877
rect 4266 843 4300 871
rect 4266 803 4300 805
rect 4266 771 4300 803
rect 4266 701 4300 733
rect 4266 699 4300 701
rect 4266 633 4300 661
rect 4266 627 4300 633
rect 4266 565 4300 589
rect 4266 555 4300 565
rect 4266 497 4300 517
rect 4266 483 4300 497
rect 4266 429 4300 445
rect 4266 411 4300 429
rect 4266 361 4300 373
rect 4266 339 4300 361
rect 4266 293 4300 301
rect 4266 267 4300 293
rect 2494 112 2528 146
rect 2788 96 2822 130
rect 3112 80 3146 114
rect 3786 70 3820 104
rect 1498 -6 1720 30
rect 5356 1402 5390 1436
rect 6720 1408 6754 1442
rect 4882 1211 4916 1237
rect 4882 1203 4916 1211
rect 4882 1143 4916 1165
rect 4882 1131 4916 1143
rect 4882 1075 4916 1093
rect 4882 1059 4916 1075
rect 4882 1007 4916 1021
rect 4882 987 4916 1007
rect 4882 939 4916 949
rect 4882 915 4916 939
rect 4882 871 4916 877
rect 4882 843 4916 871
rect 4882 803 4916 805
rect 4882 771 4916 803
rect 4882 701 4916 733
rect 4882 699 4916 701
rect 4882 633 4916 661
rect 4882 627 4916 633
rect 4882 565 4916 589
rect 4882 555 4916 565
rect 4882 497 4916 517
rect 4882 483 4916 497
rect 4882 429 4916 445
rect 4882 411 4916 429
rect 4882 361 4916 373
rect 4882 339 4916 361
rect 4882 293 4916 301
rect 4882 267 4916 293
rect 4978 1211 5012 1237
rect 4978 1203 5012 1211
rect 4978 1143 5012 1165
rect 4978 1131 5012 1143
rect 4978 1075 5012 1093
rect 4978 1059 5012 1075
rect 4978 1007 5012 1021
rect 4978 987 5012 1007
rect 4978 939 5012 949
rect 4978 915 5012 939
rect 4978 871 5012 877
rect 4978 843 5012 871
rect 4978 803 5012 805
rect 4978 771 5012 803
rect 4978 701 5012 733
rect 4978 699 5012 701
rect 4978 633 5012 661
rect 4978 627 5012 633
rect 4978 565 5012 589
rect 4978 555 5012 565
rect 4978 497 5012 517
rect 4978 483 5012 497
rect 4978 429 5012 445
rect 4978 411 5012 429
rect 4978 361 5012 373
rect 4978 339 5012 361
rect 4978 293 5012 301
rect 4978 267 5012 293
rect 5074 1211 5108 1237
rect 5074 1203 5108 1211
rect 5074 1143 5108 1165
rect 5074 1131 5108 1143
rect 5074 1075 5108 1093
rect 5074 1059 5108 1075
rect 5074 1007 5108 1021
rect 5074 987 5108 1007
rect 5074 939 5108 949
rect 5074 915 5108 939
rect 5074 871 5108 877
rect 5074 843 5108 871
rect 5074 803 5108 805
rect 5074 771 5108 803
rect 5074 701 5108 733
rect 5074 699 5108 701
rect 5074 633 5108 661
rect 5074 627 5108 633
rect 5074 565 5108 589
rect 5074 555 5108 565
rect 5074 497 5108 517
rect 5074 483 5108 497
rect 5074 429 5108 445
rect 5074 411 5108 429
rect 5074 361 5108 373
rect 5074 339 5108 361
rect 5074 293 5108 301
rect 5074 267 5108 293
rect 5170 1211 5204 1237
rect 5170 1203 5204 1211
rect 5170 1143 5204 1165
rect 5170 1131 5204 1143
rect 5170 1075 5204 1093
rect 5170 1059 5204 1075
rect 5170 1007 5204 1021
rect 5170 987 5204 1007
rect 5170 939 5204 949
rect 5170 915 5204 939
rect 5170 871 5204 877
rect 5170 843 5204 871
rect 5170 803 5204 805
rect 5170 771 5204 803
rect 5170 701 5204 733
rect 5170 699 5204 701
rect 5170 633 5204 661
rect 5170 627 5204 633
rect 5170 565 5204 589
rect 5170 555 5204 565
rect 5170 497 5204 517
rect 5170 483 5204 497
rect 5170 429 5204 445
rect 5170 411 5204 429
rect 5170 361 5204 373
rect 5170 339 5204 361
rect 5170 293 5204 301
rect 5170 267 5204 293
rect 5266 1211 5300 1237
rect 5266 1203 5300 1211
rect 5266 1143 5300 1165
rect 5266 1131 5300 1143
rect 5266 1075 5300 1093
rect 5266 1059 5300 1075
rect 5266 1007 5300 1021
rect 5266 987 5300 1007
rect 5266 939 5300 949
rect 5266 915 5300 939
rect 5266 871 5300 877
rect 5266 843 5300 871
rect 5266 803 5300 805
rect 5266 771 5300 803
rect 5266 701 5300 733
rect 5266 699 5300 701
rect 5266 633 5300 661
rect 5266 627 5300 633
rect 5266 565 5300 589
rect 5266 555 5300 565
rect 5266 497 5300 517
rect 5266 483 5300 497
rect 5266 429 5300 445
rect 5266 411 5300 429
rect 5266 361 5300 373
rect 5266 339 5300 361
rect 5266 293 5300 301
rect 5266 267 5300 293
rect 5362 1211 5396 1237
rect 5362 1203 5396 1211
rect 5362 1143 5396 1165
rect 5362 1131 5396 1143
rect 5362 1075 5396 1093
rect 5362 1059 5396 1075
rect 5362 1007 5396 1021
rect 5362 987 5396 1007
rect 5362 939 5396 949
rect 5362 915 5396 939
rect 5362 871 5396 877
rect 5362 843 5396 871
rect 5362 803 5396 805
rect 5362 771 5396 803
rect 5362 701 5396 733
rect 5362 699 5396 701
rect 5362 633 5396 661
rect 5362 627 5396 633
rect 5362 565 5396 589
rect 5362 555 5396 565
rect 5362 497 5396 517
rect 5362 483 5396 497
rect 5362 429 5396 445
rect 5362 411 5396 429
rect 5362 361 5396 373
rect 5362 339 5396 361
rect 5362 293 5396 301
rect 5362 267 5396 293
rect 5458 1211 5492 1237
rect 5458 1203 5492 1211
rect 5458 1143 5492 1165
rect 5458 1131 5492 1143
rect 5458 1075 5492 1093
rect 5458 1059 5492 1075
rect 5458 1007 5492 1021
rect 5458 987 5492 1007
rect 5458 939 5492 949
rect 5458 915 5492 939
rect 5458 871 5492 877
rect 5458 843 5492 871
rect 5458 803 5492 805
rect 5458 771 5492 803
rect 5458 701 5492 733
rect 5458 699 5492 701
rect 5458 633 5492 661
rect 5458 627 5492 633
rect 5458 565 5492 589
rect 5458 555 5492 565
rect 5458 497 5492 517
rect 5458 483 5492 497
rect 5458 429 5492 445
rect 5458 411 5492 429
rect 5458 361 5492 373
rect 5458 339 5492 361
rect 5458 293 5492 301
rect 5458 267 5492 293
rect 5554 1211 5588 1237
rect 5554 1203 5588 1211
rect 5554 1143 5588 1165
rect 5554 1131 5588 1143
rect 5554 1075 5588 1093
rect 5554 1059 5588 1075
rect 5554 1007 5588 1021
rect 5554 987 5588 1007
rect 5554 939 5588 949
rect 5554 915 5588 939
rect 5554 871 5588 877
rect 5554 843 5588 871
rect 5554 803 5588 805
rect 5554 771 5588 803
rect 5554 701 5588 733
rect 5554 699 5588 701
rect 5554 633 5588 661
rect 5554 627 5588 633
rect 5554 565 5588 589
rect 5554 555 5588 565
rect 5554 497 5588 517
rect 5554 483 5588 497
rect 5554 429 5588 445
rect 5554 411 5588 429
rect 5554 361 5588 373
rect 5554 339 5588 361
rect 5554 293 5588 301
rect 5554 267 5588 293
rect 5650 1211 5684 1237
rect 5650 1203 5684 1211
rect 5650 1143 5684 1165
rect 5650 1131 5684 1143
rect 5650 1075 5684 1093
rect 5650 1059 5684 1075
rect 5650 1007 5684 1021
rect 5650 987 5684 1007
rect 5650 939 5684 949
rect 5650 915 5684 939
rect 5650 871 5684 877
rect 5650 843 5684 871
rect 5650 803 5684 805
rect 5650 771 5684 803
rect 5650 701 5684 733
rect 5650 699 5684 701
rect 5650 633 5684 661
rect 5650 627 5684 633
rect 5650 565 5684 589
rect 5650 555 5684 565
rect 5650 497 5684 517
rect 5650 483 5684 497
rect 5650 429 5684 445
rect 5650 411 5684 429
rect 5650 361 5684 373
rect 5650 339 5684 361
rect 5650 293 5684 301
rect 5650 267 5684 293
rect 5746 1211 5780 1237
rect 5746 1203 5780 1211
rect 5746 1143 5780 1165
rect 5746 1131 5780 1143
rect 5746 1075 5780 1093
rect 5746 1059 5780 1075
rect 5746 1007 5780 1021
rect 5746 987 5780 1007
rect 5746 939 5780 949
rect 5746 915 5780 939
rect 5746 871 5780 877
rect 5746 843 5780 871
rect 5746 803 5780 805
rect 5746 771 5780 803
rect 5746 701 5780 733
rect 5746 699 5780 701
rect 5746 633 5780 661
rect 5746 627 5780 633
rect 5746 565 5780 589
rect 5746 555 5780 565
rect 5746 497 5780 517
rect 5746 483 5780 497
rect 5746 429 5780 445
rect 5746 411 5780 429
rect 5746 361 5780 373
rect 5746 339 5780 361
rect 5746 293 5780 301
rect 5746 267 5780 293
rect 5842 1211 5876 1237
rect 5842 1203 5876 1211
rect 5842 1143 5876 1165
rect 5842 1131 5876 1143
rect 5842 1075 5876 1093
rect 5842 1059 5876 1075
rect 5842 1007 5876 1021
rect 5842 987 5876 1007
rect 5842 939 5876 949
rect 5842 915 5876 939
rect 5842 871 5876 877
rect 5842 843 5876 871
rect 5842 803 5876 805
rect 5842 771 5876 803
rect 5842 701 5876 733
rect 5842 699 5876 701
rect 5842 633 5876 661
rect 5842 627 5876 633
rect 5842 565 5876 589
rect 5842 555 5876 565
rect 5842 497 5876 517
rect 5842 483 5876 497
rect 5842 429 5876 445
rect 5842 411 5876 429
rect 5842 361 5876 373
rect 5842 339 5876 361
rect 5842 293 5876 301
rect 5842 267 5876 293
rect 5938 1211 5972 1237
rect 5938 1203 5972 1211
rect 5938 1143 5972 1165
rect 5938 1131 5972 1143
rect 5938 1075 5972 1093
rect 5938 1059 5972 1075
rect 5938 1007 5972 1021
rect 5938 987 5972 1007
rect 5938 939 5972 949
rect 5938 915 5972 939
rect 5938 871 5972 877
rect 5938 843 5972 871
rect 5938 803 5972 805
rect 5938 771 5972 803
rect 5938 701 5972 733
rect 5938 699 5972 701
rect 5938 633 5972 661
rect 5938 627 5972 633
rect 5938 565 5972 589
rect 5938 555 5972 565
rect 5938 497 5972 517
rect 5938 483 5972 497
rect 5938 429 5972 445
rect 5938 411 5972 429
rect 5938 361 5972 373
rect 5938 339 5972 361
rect 5938 293 5972 301
rect 5938 267 5972 293
rect 6144 1211 6178 1237
rect 6144 1203 6178 1211
rect 6144 1143 6178 1165
rect 6144 1131 6178 1143
rect 6144 1075 6178 1093
rect 6144 1059 6178 1075
rect 6144 1007 6178 1021
rect 6144 987 6178 1007
rect 6144 939 6178 949
rect 6144 915 6178 939
rect 6144 871 6178 877
rect 6144 843 6178 871
rect 6144 803 6178 805
rect 6144 771 6178 803
rect 6144 701 6178 733
rect 6144 699 6178 701
rect 6144 633 6178 661
rect 6144 627 6178 633
rect 6144 565 6178 589
rect 6144 555 6178 565
rect 6144 497 6178 517
rect 6144 483 6178 497
rect 6144 429 6178 445
rect 6144 411 6178 429
rect 6144 361 6178 373
rect 6144 339 6178 361
rect 6144 293 6178 301
rect 6144 267 6178 293
rect 6240 1211 6274 1237
rect 6240 1203 6274 1211
rect 6240 1143 6274 1165
rect 6240 1131 6274 1143
rect 6240 1075 6274 1093
rect 6240 1059 6274 1075
rect 6240 1007 6274 1021
rect 6240 987 6274 1007
rect 6240 939 6274 949
rect 6240 915 6274 939
rect 6240 871 6274 877
rect 6240 843 6274 871
rect 6240 803 6274 805
rect 6240 771 6274 803
rect 6240 701 6274 733
rect 6240 699 6274 701
rect 6240 633 6274 661
rect 6240 627 6274 633
rect 6240 565 6274 589
rect 6240 555 6274 565
rect 6240 497 6274 517
rect 6240 483 6274 497
rect 6240 429 6274 445
rect 6240 411 6274 429
rect 6240 361 6274 373
rect 6240 339 6274 361
rect 6240 293 6274 301
rect 6240 267 6274 293
rect 6336 1211 6370 1237
rect 6336 1203 6370 1211
rect 6336 1143 6370 1165
rect 6336 1131 6370 1143
rect 6336 1075 6370 1093
rect 6336 1059 6370 1075
rect 6336 1007 6370 1021
rect 6336 987 6370 1007
rect 6336 939 6370 949
rect 6336 915 6370 939
rect 6336 871 6370 877
rect 6336 843 6370 871
rect 6336 803 6370 805
rect 6336 771 6370 803
rect 6336 701 6370 733
rect 6336 699 6370 701
rect 6336 633 6370 661
rect 6336 627 6370 633
rect 6336 565 6370 589
rect 6336 555 6370 565
rect 6336 497 6370 517
rect 6336 483 6370 497
rect 6336 429 6370 445
rect 6336 411 6370 429
rect 6336 361 6370 373
rect 6336 339 6370 361
rect 6336 293 6370 301
rect 6336 267 6370 293
rect 6432 1211 6466 1237
rect 6432 1203 6466 1211
rect 6432 1143 6466 1165
rect 6432 1131 6466 1143
rect 6432 1075 6466 1093
rect 6432 1059 6466 1075
rect 6432 1007 6466 1021
rect 6432 987 6466 1007
rect 6432 939 6466 949
rect 6432 915 6466 939
rect 6432 871 6466 877
rect 6432 843 6466 871
rect 6432 803 6466 805
rect 6432 771 6466 803
rect 6432 701 6466 733
rect 6432 699 6466 701
rect 6432 633 6466 661
rect 6432 627 6466 633
rect 6432 565 6466 589
rect 6432 555 6466 565
rect 6432 497 6466 517
rect 6432 483 6466 497
rect 6432 429 6466 445
rect 6432 411 6466 429
rect 6432 361 6466 373
rect 6432 339 6466 361
rect 6432 293 6466 301
rect 6432 267 6466 293
rect 6528 1211 6562 1237
rect 6528 1203 6562 1211
rect 6528 1143 6562 1165
rect 6528 1131 6562 1143
rect 6528 1075 6562 1093
rect 6528 1059 6562 1075
rect 6528 1007 6562 1021
rect 6528 987 6562 1007
rect 6528 939 6562 949
rect 6528 915 6562 939
rect 6528 871 6562 877
rect 6528 843 6562 871
rect 6528 803 6562 805
rect 6528 771 6562 803
rect 6528 701 6562 733
rect 6528 699 6562 701
rect 6528 633 6562 661
rect 6528 627 6562 633
rect 6528 565 6562 589
rect 6528 555 6562 565
rect 6528 497 6562 517
rect 6528 483 6562 497
rect 6528 429 6562 445
rect 6528 411 6562 429
rect 6528 361 6562 373
rect 6528 339 6562 361
rect 6528 293 6562 301
rect 6528 267 6562 293
rect 6624 1211 6658 1237
rect 6624 1203 6658 1211
rect 6624 1143 6658 1165
rect 6624 1131 6658 1143
rect 6624 1075 6658 1093
rect 6624 1059 6658 1075
rect 6624 1007 6658 1021
rect 6624 987 6658 1007
rect 6624 939 6658 949
rect 6624 915 6658 939
rect 6624 871 6658 877
rect 6624 843 6658 871
rect 6624 803 6658 805
rect 6624 771 6658 803
rect 6624 701 6658 733
rect 6624 699 6658 701
rect 6624 633 6658 661
rect 6624 627 6658 633
rect 6624 565 6658 589
rect 6624 555 6658 565
rect 6624 497 6658 517
rect 6624 483 6658 497
rect 6624 429 6658 445
rect 6624 411 6658 429
rect 6624 361 6658 373
rect 6624 339 6658 361
rect 6624 293 6658 301
rect 6624 267 6658 293
rect 6720 1211 6754 1237
rect 6720 1203 6754 1211
rect 6720 1143 6754 1165
rect 6720 1131 6754 1143
rect 6720 1075 6754 1093
rect 6720 1059 6754 1075
rect 6720 1007 6754 1021
rect 6720 987 6754 1007
rect 6720 939 6754 949
rect 6720 915 6754 939
rect 6720 871 6754 877
rect 6720 843 6754 871
rect 6720 803 6754 805
rect 6720 771 6754 803
rect 6720 701 6754 733
rect 6720 699 6754 701
rect 6720 633 6754 661
rect 6720 627 6754 633
rect 6720 565 6754 589
rect 6720 555 6754 565
rect 6720 497 6754 517
rect 6720 483 6754 497
rect 6720 429 6754 445
rect 6720 411 6754 429
rect 6720 361 6754 373
rect 6720 339 6754 361
rect 6720 293 6754 301
rect 6720 267 6754 293
rect 6816 1211 6850 1237
rect 6816 1203 6850 1211
rect 6816 1143 6850 1165
rect 6816 1131 6850 1143
rect 6816 1075 6850 1093
rect 6816 1059 6850 1075
rect 6816 1007 6850 1021
rect 6816 987 6850 1007
rect 6816 939 6850 949
rect 6816 915 6850 939
rect 6816 871 6850 877
rect 6816 843 6850 871
rect 6816 803 6850 805
rect 6816 771 6850 803
rect 6816 701 6850 733
rect 6816 699 6850 701
rect 6816 633 6850 661
rect 6816 627 6850 633
rect 6816 565 6850 589
rect 6816 555 6850 565
rect 6816 497 6850 517
rect 6816 483 6850 497
rect 6816 429 6850 445
rect 6816 411 6850 429
rect 6816 361 6850 373
rect 6816 339 6850 361
rect 6816 293 6850 301
rect 6816 267 6850 293
rect 6912 1211 6946 1237
rect 6912 1203 6946 1211
rect 6912 1143 6946 1165
rect 6912 1131 6946 1143
rect 6912 1075 6946 1093
rect 6912 1059 6946 1075
rect 6912 1007 6946 1021
rect 6912 987 6946 1007
rect 6912 939 6946 949
rect 6912 915 6946 939
rect 6912 871 6946 877
rect 6912 843 6946 871
rect 6912 803 6946 805
rect 6912 771 6946 803
rect 6912 701 6946 733
rect 6912 699 6946 701
rect 6912 633 6946 661
rect 6912 627 6946 633
rect 6912 565 6946 589
rect 6912 555 6946 565
rect 6912 497 6946 517
rect 6912 483 6946 497
rect 6912 429 6946 445
rect 6912 411 6946 429
rect 6912 361 6946 373
rect 6912 339 6946 361
rect 6912 293 6946 301
rect 6912 267 6946 293
rect 7008 1211 7042 1237
rect 7008 1203 7042 1211
rect 7008 1143 7042 1165
rect 7008 1131 7042 1143
rect 7008 1075 7042 1093
rect 7008 1059 7042 1075
rect 7008 1007 7042 1021
rect 7008 987 7042 1007
rect 7008 939 7042 949
rect 7008 915 7042 939
rect 7008 871 7042 877
rect 7008 843 7042 871
rect 7008 803 7042 805
rect 7008 771 7042 803
rect 7008 701 7042 733
rect 7008 699 7042 701
rect 7008 633 7042 661
rect 7008 627 7042 633
rect 7008 565 7042 589
rect 7008 555 7042 565
rect 7008 497 7042 517
rect 7008 483 7042 497
rect 7008 429 7042 445
rect 7008 411 7042 429
rect 7008 361 7042 373
rect 7008 339 7042 361
rect 7008 293 7042 301
rect 7008 267 7042 293
rect 7104 1211 7138 1237
rect 7104 1203 7138 1211
rect 7104 1143 7138 1165
rect 7104 1131 7138 1143
rect 7104 1075 7138 1093
rect 7104 1059 7138 1075
rect 7104 1007 7138 1021
rect 7104 987 7138 1007
rect 7104 939 7138 949
rect 7104 915 7138 939
rect 7104 871 7138 877
rect 7104 843 7138 871
rect 7104 803 7138 805
rect 7104 771 7138 803
rect 7104 701 7138 733
rect 7104 699 7138 701
rect 7104 633 7138 661
rect 7104 627 7138 633
rect 7104 565 7138 589
rect 7104 555 7138 565
rect 7104 497 7138 517
rect 7104 483 7138 497
rect 7104 429 7138 445
rect 7104 411 7138 429
rect 7104 361 7138 373
rect 7104 339 7138 361
rect 7104 293 7138 301
rect 7104 267 7138 293
rect 7200 1211 7234 1237
rect 7200 1203 7234 1211
rect 7200 1143 7234 1165
rect 7200 1131 7234 1143
rect 7200 1075 7234 1093
rect 7200 1059 7234 1075
rect 7200 1007 7234 1021
rect 7200 987 7234 1007
rect 7200 939 7234 949
rect 7200 915 7234 939
rect 7200 871 7234 877
rect 7200 843 7234 871
rect 7200 803 7234 805
rect 7200 771 7234 803
rect 7200 701 7234 733
rect 7200 699 7234 701
rect 7200 633 7234 661
rect 7200 627 7234 633
rect 7200 565 7234 589
rect 7200 555 7234 565
rect 7200 497 7234 517
rect 7200 483 7234 497
rect 7200 429 7234 445
rect 7200 411 7234 429
rect 7200 361 7234 373
rect 7200 339 7234 361
rect 7200 293 7234 301
rect 7200 267 7234 293
rect 7296 1211 7330 1237
rect 7296 1203 7330 1211
rect 7296 1143 7330 1165
rect 7296 1131 7330 1143
rect 7296 1075 7330 1093
rect 7296 1059 7330 1075
rect 7296 1007 7330 1021
rect 7296 987 7330 1007
rect 7296 939 7330 949
rect 7296 915 7330 939
rect 7296 871 7330 877
rect 7296 843 7330 871
rect 7296 803 7330 805
rect 7296 771 7330 803
rect 7296 701 7330 733
rect 7296 699 7330 701
rect 7296 633 7330 661
rect 7296 627 7330 633
rect 7296 565 7330 589
rect 7296 555 7330 565
rect 7296 497 7330 517
rect 7296 483 7330 497
rect 7296 429 7330 445
rect 7296 411 7330 429
rect 7296 361 7330 373
rect 7296 339 7330 361
rect 7296 293 7330 301
rect 7296 267 7330 293
rect 5450 96 5484 130
rect 5744 80 5778 114
rect 6142 80 6176 114
rect 6816 70 6850 104
rect 4584 -24 4806 12
rect 8386 1402 8420 1436
rect 9808 1406 9842 1440
rect 7912 1211 7946 1237
rect 7912 1203 7946 1211
rect 7912 1143 7946 1165
rect 7912 1131 7946 1143
rect 7912 1075 7946 1093
rect 7912 1059 7946 1075
rect 7912 1007 7946 1021
rect 7912 987 7946 1007
rect 7912 939 7946 949
rect 7912 915 7946 939
rect 7912 871 7946 877
rect 7912 843 7946 871
rect 7912 803 7946 805
rect 7912 771 7946 803
rect 7912 701 7946 733
rect 7912 699 7946 701
rect 7912 633 7946 661
rect 7912 627 7946 633
rect 7912 565 7946 589
rect 7912 555 7946 565
rect 7912 497 7946 517
rect 7912 483 7946 497
rect 7912 429 7946 445
rect 7912 411 7946 429
rect 7912 361 7946 373
rect 7912 339 7946 361
rect 7912 293 7946 301
rect 7912 267 7946 293
rect 8008 1211 8042 1237
rect 8008 1203 8042 1211
rect 8008 1143 8042 1165
rect 8008 1131 8042 1143
rect 8008 1075 8042 1093
rect 8008 1059 8042 1075
rect 8008 1007 8042 1021
rect 8008 987 8042 1007
rect 8008 939 8042 949
rect 8008 915 8042 939
rect 8008 871 8042 877
rect 8008 843 8042 871
rect 8008 803 8042 805
rect 8008 771 8042 803
rect 8008 701 8042 733
rect 8008 699 8042 701
rect 8008 633 8042 661
rect 8008 627 8042 633
rect 8008 565 8042 589
rect 8008 555 8042 565
rect 8008 497 8042 517
rect 8008 483 8042 497
rect 8008 429 8042 445
rect 8008 411 8042 429
rect 8008 361 8042 373
rect 8008 339 8042 361
rect 8008 293 8042 301
rect 8008 267 8042 293
rect 8104 1211 8138 1237
rect 8104 1203 8138 1211
rect 8104 1143 8138 1165
rect 8104 1131 8138 1143
rect 8104 1075 8138 1093
rect 8104 1059 8138 1075
rect 8104 1007 8138 1021
rect 8104 987 8138 1007
rect 8104 939 8138 949
rect 8104 915 8138 939
rect 8104 871 8138 877
rect 8104 843 8138 871
rect 8104 803 8138 805
rect 8104 771 8138 803
rect 8104 701 8138 733
rect 8104 699 8138 701
rect 8104 633 8138 661
rect 8104 627 8138 633
rect 8104 565 8138 589
rect 8104 555 8138 565
rect 8104 497 8138 517
rect 8104 483 8138 497
rect 8104 429 8138 445
rect 8104 411 8138 429
rect 8104 361 8138 373
rect 8104 339 8138 361
rect 8104 293 8138 301
rect 8104 267 8138 293
rect 8200 1211 8234 1237
rect 8200 1203 8234 1211
rect 8200 1143 8234 1165
rect 8200 1131 8234 1143
rect 8200 1075 8234 1093
rect 8200 1059 8234 1075
rect 8200 1007 8234 1021
rect 8200 987 8234 1007
rect 8200 939 8234 949
rect 8200 915 8234 939
rect 8200 871 8234 877
rect 8200 843 8234 871
rect 8200 803 8234 805
rect 8200 771 8234 803
rect 8200 701 8234 733
rect 8200 699 8234 701
rect 8200 633 8234 661
rect 8200 627 8234 633
rect 8200 565 8234 589
rect 8200 555 8234 565
rect 8200 497 8234 517
rect 8200 483 8234 497
rect 8200 429 8234 445
rect 8200 411 8234 429
rect 8200 361 8234 373
rect 8200 339 8234 361
rect 8200 293 8234 301
rect 8200 267 8234 293
rect 8296 1211 8330 1237
rect 8296 1203 8330 1211
rect 8296 1143 8330 1165
rect 8296 1131 8330 1143
rect 8296 1075 8330 1093
rect 8296 1059 8330 1075
rect 8296 1007 8330 1021
rect 8296 987 8330 1007
rect 8296 939 8330 949
rect 8296 915 8330 939
rect 8296 871 8330 877
rect 8296 843 8330 871
rect 8296 803 8330 805
rect 8296 771 8330 803
rect 8296 701 8330 733
rect 8296 699 8330 701
rect 8296 633 8330 661
rect 8296 627 8330 633
rect 8296 565 8330 589
rect 8296 555 8330 565
rect 8296 497 8330 517
rect 8296 483 8330 497
rect 8296 429 8330 445
rect 8296 411 8330 429
rect 8296 361 8330 373
rect 8296 339 8330 361
rect 8296 293 8330 301
rect 8296 267 8330 293
rect 8392 1211 8426 1237
rect 8392 1203 8426 1211
rect 8392 1143 8426 1165
rect 8392 1131 8426 1143
rect 8392 1075 8426 1093
rect 8392 1059 8426 1075
rect 8392 1007 8426 1021
rect 8392 987 8426 1007
rect 8392 939 8426 949
rect 8392 915 8426 939
rect 8392 871 8426 877
rect 8392 843 8426 871
rect 8392 803 8426 805
rect 8392 771 8426 803
rect 8392 701 8426 733
rect 8392 699 8426 701
rect 8392 633 8426 661
rect 8392 627 8426 633
rect 8392 565 8426 589
rect 8392 555 8426 565
rect 8392 497 8426 517
rect 8392 483 8426 497
rect 8392 429 8426 445
rect 8392 411 8426 429
rect 8392 361 8426 373
rect 8392 339 8426 361
rect 8392 293 8426 301
rect 8392 267 8426 293
rect 8488 1211 8522 1237
rect 8488 1203 8522 1211
rect 8488 1143 8522 1165
rect 8488 1131 8522 1143
rect 8488 1075 8522 1093
rect 8488 1059 8522 1075
rect 8488 1007 8522 1021
rect 8488 987 8522 1007
rect 8488 939 8522 949
rect 8488 915 8522 939
rect 8488 871 8522 877
rect 8488 843 8522 871
rect 8488 803 8522 805
rect 8488 771 8522 803
rect 8488 701 8522 733
rect 8488 699 8522 701
rect 8488 633 8522 661
rect 8488 627 8522 633
rect 8488 565 8522 589
rect 8488 555 8522 565
rect 8488 497 8522 517
rect 8488 483 8522 497
rect 8488 429 8522 445
rect 8488 411 8522 429
rect 8488 361 8522 373
rect 8488 339 8522 361
rect 8488 293 8522 301
rect 8488 267 8522 293
rect 8584 1211 8618 1237
rect 8584 1203 8618 1211
rect 8584 1143 8618 1165
rect 8584 1131 8618 1143
rect 8584 1075 8618 1093
rect 8584 1059 8618 1075
rect 8584 1007 8618 1021
rect 8584 987 8618 1007
rect 8584 939 8618 949
rect 8584 915 8618 939
rect 8584 871 8618 877
rect 8584 843 8618 871
rect 8584 803 8618 805
rect 8584 771 8618 803
rect 8584 701 8618 733
rect 8584 699 8618 701
rect 8584 633 8618 661
rect 8584 627 8618 633
rect 8584 565 8618 589
rect 8584 555 8618 565
rect 8584 497 8618 517
rect 8584 483 8618 497
rect 8584 429 8618 445
rect 8584 411 8618 429
rect 8584 361 8618 373
rect 8584 339 8618 361
rect 8584 293 8618 301
rect 8584 267 8618 293
rect 8680 1211 8714 1237
rect 8680 1203 8714 1211
rect 8680 1143 8714 1165
rect 8680 1131 8714 1143
rect 8680 1075 8714 1093
rect 8680 1059 8714 1075
rect 8680 1007 8714 1021
rect 8680 987 8714 1007
rect 8680 939 8714 949
rect 8680 915 8714 939
rect 8680 871 8714 877
rect 8680 843 8714 871
rect 8680 803 8714 805
rect 8680 771 8714 803
rect 8680 701 8714 733
rect 8680 699 8714 701
rect 8680 633 8714 661
rect 8680 627 8714 633
rect 8680 565 8714 589
rect 8680 555 8714 565
rect 8680 497 8714 517
rect 8680 483 8714 497
rect 8680 429 8714 445
rect 8680 411 8714 429
rect 8680 361 8714 373
rect 8680 339 8714 361
rect 8680 293 8714 301
rect 8680 267 8714 293
rect 8776 1211 8810 1237
rect 8776 1203 8810 1211
rect 8776 1143 8810 1165
rect 8776 1131 8810 1143
rect 8776 1075 8810 1093
rect 8776 1059 8810 1075
rect 8776 1007 8810 1021
rect 8776 987 8810 1007
rect 8776 939 8810 949
rect 8776 915 8810 939
rect 8776 871 8810 877
rect 8776 843 8810 871
rect 8776 803 8810 805
rect 8776 771 8810 803
rect 8776 701 8810 733
rect 8776 699 8810 701
rect 8776 633 8810 661
rect 8776 627 8810 633
rect 8776 565 8810 589
rect 8776 555 8810 565
rect 8776 497 8810 517
rect 8776 483 8810 497
rect 8776 429 8810 445
rect 8776 411 8810 429
rect 8776 361 8810 373
rect 8776 339 8810 361
rect 8776 293 8810 301
rect 8776 267 8810 293
rect 8872 1211 8906 1237
rect 8872 1203 8906 1211
rect 8872 1143 8906 1165
rect 8872 1131 8906 1143
rect 8872 1075 8906 1093
rect 8872 1059 8906 1075
rect 8872 1007 8906 1021
rect 8872 987 8906 1007
rect 8872 939 8906 949
rect 8872 915 8906 939
rect 8872 871 8906 877
rect 8872 843 8906 871
rect 8872 803 8906 805
rect 8872 771 8906 803
rect 8872 701 8906 733
rect 8872 699 8906 701
rect 8872 633 8906 661
rect 8872 627 8906 633
rect 8872 565 8906 589
rect 8872 555 8906 565
rect 8872 497 8906 517
rect 8872 483 8906 497
rect 8872 429 8906 445
rect 8872 411 8906 429
rect 8872 361 8906 373
rect 8872 339 8906 361
rect 8872 293 8906 301
rect 8872 267 8906 293
rect 8968 1211 9002 1237
rect 8968 1203 9002 1211
rect 8968 1143 9002 1165
rect 8968 1131 9002 1143
rect 8968 1075 9002 1093
rect 8968 1059 9002 1075
rect 8968 1007 9002 1021
rect 8968 987 9002 1007
rect 8968 939 9002 949
rect 8968 915 9002 939
rect 8968 871 9002 877
rect 8968 843 9002 871
rect 8968 803 9002 805
rect 8968 771 9002 803
rect 8968 701 9002 733
rect 8968 699 9002 701
rect 8968 633 9002 661
rect 8968 627 9002 633
rect 8968 565 9002 589
rect 8968 555 9002 565
rect 8968 497 9002 517
rect 8968 483 9002 497
rect 8968 429 9002 445
rect 8968 411 9002 429
rect 8968 361 9002 373
rect 8968 339 9002 361
rect 8968 293 9002 301
rect 8968 267 9002 293
rect 9232 1209 9266 1235
rect 9232 1201 9266 1209
rect 9232 1141 9266 1163
rect 9232 1129 9266 1141
rect 9232 1073 9266 1091
rect 9232 1057 9266 1073
rect 9232 1005 9266 1019
rect 9232 985 9266 1005
rect 9232 937 9266 947
rect 9232 913 9266 937
rect 9232 869 9266 875
rect 9232 841 9266 869
rect 9232 801 9266 803
rect 9232 769 9266 801
rect 9232 699 9266 731
rect 9232 697 9266 699
rect 9232 631 9266 659
rect 9232 625 9266 631
rect 9232 563 9266 587
rect 9232 553 9266 563
rect 9232 495 9266 515
rect 9232 481 9266 495
rect 9232 427 9266 443
rect 9232 409 9266 427
rect 9232 359 9266 371
rect 9232 337 9266 359
rect 9232 291 9266 299
rect 9232 265 9266 291
rect 9328 1209 9362 1235
rect 9328 1201 9362 1209
rect 9328 1141 9362 1163
rect 9328 1129 9362 1141
rect 9328 1073 9362 1091
rect 9328 1057 9362 1073
rect 9328 1005 9362 1019
rect 9328 985 9362 1005
rect 9328 937 9362 947
rect 9328 913 9362 937
rect 9328 869 9362 875
rect 9328 841 9362 869
rect 9328 801 9362 803
rect 9328 769 9362 801
rect 9328 699 9362 731
rect 9328 697 9362 699
rect 9328 631 9362 659
rect 9328 625 9362 631
rect 9328 563 9362 587
rect 9328 553 9362 563
rect 9328 495 9362 515
rect 9328 481 9362 495
rect 9328 427 9362 443
rect 9328 409 9362 427
rect 9328 359 9362 371
rect 9328 337 9362 359
rect 9328 291 9362 299
rect 9328 265 9362 291
rect 9424 1209 9458 1235
rect 9424 1201 9458 1209
rect 9424 1141 9458 1163
rect 9424 1129 9458 1141
rect 9424 1073 9458 1091
rect 9424 1057 9458 1073
rect 9424 1005 9458 1019
rect 9424 985 9458 1005
rect 9424 937 9458 947
rect 9424 913 9458 937
rect 9424 869 9458 875
rect 9424 841 9458 869
rect 9424 801 9458 803
rect 9424 769 9458 801
rect 9424 699 9458 731
rect 9424 697 9458 699
rect 9424 631 9458 659
rect 9424 625 9458 631
rect 9424 563 9458 587
rect 9424 553 9458 563
rect 9424 495 9458 515
rect 9424 481 9458 495
rect 9424 427 9458 443
rect 9424 409 9458 427
rect 9424 359 9458 371
rect 9424 337 9458 359
rect 9424 291 9458 299
rect 9424 265 9458 291
rect 9520 1209 9554 1235
rect 9520 1201 9554 1209
rect 9520 1141 9554 1163
rect 9520 1129 9554 1141
rect 9520 1073 9554 1091
rect 9520 1057 9554 1073
rect 9520 1005 9554 1019
rect 9520 985 9554 1005
rect 9520 937 9554 947
rect 9520 913 9554 937
rect 9520 869 9554 875
rect 9520 841 9554 869
rect 9520 801 9554 803
rect 9520 769 9554 801
rect 9520 699 9554 731
rect 9520 697 9554 699
rect 9520 631 9554 659
rect 9520 625 9554 631
rect 9520 563 9554 587
rect 9520 553 9554 563
rect 9520 495 9554 515
rect 9520 481 9554 495
rect 9520 427 9554 443
rect 9520 409 9554 427
rect 9520 359 9554 371
rect 9520 337 9554 359
rect 9520 291 9554 299
rect 9520 265 9554 291
rect 9616 1209 9650 1235
rect 9616 1201 9650 1209
rect 9616 1141 9650 1163
rect 9616 1129 9650 1141
rect 9616 1073 9650 1091
rect 9616 1057 9650 1073
rect 9616 1005 9650 1019
rect 9616 985 9650 1005
rect 9616 937 9650 947
rect 9616 913 9650 937
rect 9616 869 9650 875
rect 9616 841 9650 869
rect 9616 801 9650 803
rect 9616 769 9650 801
rect 9616 699 9650 731
rect 9616 697 9650 699
rect 9616 631 9650 659
rect 9616 625 9650 631
rect 9616 563 9650 587
rect 9616 553 9650 563
rect 9616 495 9650 515
rect 9616 481 9650 495
rect 9616 427 9650 443
rect 9616 409 9650 427
rect 9616 359 9650 371
rect 9616 337 9650 359
rect 9616 291 9650 299
rect 9616 265 9650 291
rect 9712 1209 9746 1235
rect 9712 1201 9746 1209
rect 9712 1141 9746 1163
rect 9712 1129 9746 1141
rect 9712 1073 9746 1091
rect 9712 1057 9746 1073
rect 9712 1005 9746 1019
rect 9712 985 9746 1005
rect 9712 937 9746 947
rect 9712 913 9746 937
rect 9712 869 9746 875
rect 9712 841 9746 869
rect 9712 801 9746 803
rect 9712 769 9746 801
rect 9712 699 9746 731
rect 9712 697 9746 699
rect 9712 631 9746 659
rect 9712 625 9746 631
rect 9712 563 9746 587
rect 9712 553 9746 563
rect 9712 495 9746 515
rect 9712 481 9746 495
rect 9712 427 9746 443
rect 9712 409 9746 427
rect 9712 359 9746 371
rect 9712 337 9746 359
rect 9712 291 9746 299
rect 9712 265 9746 291
rect 9808 1209 9842 1235
rect 9808 1201 9842 1209
rect 9808 1141 9842 1163
rect 9808 1129 9842 1141
rect 9808 1073 9842 1091
rect 9808 1057 9842 1073
rect 9808 1005 9842 1019
rect 9808 985 9842 1005
rect 9808 937 9842 947
rect 9808 913 9842 937
rect 9808 869 9842 875
rect 9808 841 9842 869
rect 9808 801 9842 803
rect 9808 769 9842 801
rect 9808 699 9842 731
rect 9808 697 9842 699
rect 9808 631 9842 659
rect 9808 625 9842 631
rect 9808 563 9842 587
rect 9808 553 9842 563
rect 9808 495 9842 515
rect 9808 481 9842 495
rect 9808 427 9842 443
rect 9808 409 9842 427
rect 9808 359 9842 371
rect 9808 337 9842 359
rect 9808 291 9842 299
rect 9808 265 9842 291
rect 9904 1209 9938 1235
rect 9904 1201 9938 1209
rect 9904 1141 9938 1163
rect 9904 1129 9938 1141
rect 9904 1073 9938 1091
rect 9904 1057 9938 1073
rect 9904 1005 9938 1019
rect 9904 985 9938 1005
rect 9904 937 9938 947
rect 9904 913 9938 937
rect 9904 869 9938 875
rect 9904 841 9938 869
rect 9904 801 9938 803
rect 9904 769 9938 801
rect 9904 699 9938 731
rect 9904 697 9938 699
rect 9904 631 9938 659
rect 9904 625 9938 631
rect 9904 563 9938 587
rect 9904 553 9938 563
rect 9904 495 9938 515
rect 9904 481 9938 495
rect 9904 427 9938 443
rect 9904 409 9938 427
rect 9904 359 9938 371
rect 9904 337 9938 359
rect 9904 291 9938 299
rect 9904 265 9938 291
rect 10000 1209 10034 1235
rect 10000 1201 10034 1209
rect 10000 1141 10034 1163
rect 10000 1129 10034 1141
rect 10000 1073 10034 1091
rect 10000 1057 10034 1073
rect 10000 1005 10034 1019
rect 10000 985 10034 1005
rect 10000 937 10034 947
rect 10000 913 10034 937
rect 10000 869 10034 875
rect 10000 841 10034 869
rect 10000 801 10034 803
rect 10000 769 10034 801
rect 10000 699 10034 731
rect 10000 697 10034 699
rect 10000 631 10034 659
rect 10000 625 10034 631
rect 10000 563 10034 587
rect 10000 553 10034 563
rect 10000 495 10034 515
rect 10000 481 10034 495
rect 10000 427 10034 443
rect 10000 409 10034 427
rect 10000 359 10034 371
rect 10000 337 10034 359
rect 10000 291 10034 299
rect 10000 265 10034 291
rect 10096 1209 10130 1235
rect 10096 1201 10130 1209
rect 10096 1141 10130 1163
rect 10096 1129 10130 1141
rect 10096 1073 10130 1091
rect 10096 1057 10130 1073
rect 10096 1005 10130 1019
rect 10096 985 10130 1005
rect 10096 937 10130 947
rect 10096 913 10130 937
rect 10096 869 10130 875
rect 10096 841 10130 869
rect 10096 801 10130 803
rect 10096 769 10130 801
rect 10096 699 10130 731
rect 10096 697 10130 699
rect 10096 631 10130 659
rect 10096 625 10130 631
rect 10096 563 10130 587
rect 10096 553 10130 563
rect 10096 495 10130 515
rect 10096 481 10130 495
rect 10096 427 10130 443
rect 10096 409 10130 427
rect 10096 359 10130 371
rect 10096 337 10130 359
rect 10096 291 10130 299
rect 10096 265 10130 291
rect 10192 1209 10226 1235
rect 10192 1201 10226 1209
rect 10192 1141 10226 1163
rect 10192 1129 10226 1141
rect 10192 1073 10226 1091
rect 10192 1057 10226 1073
rect 10192 1005 10226 1019
rect 10192 985 10226 1005
rect 10192 937 10226 947
rect 10192 913 10226 937
rect 10192 869 10226 875
rect 10192 841 10226 869
rect 10192 801 10226 803
rect 10192 769 10226 801
rect 10192 699 10226 731
rect 10192 697 10226 699
rect 10192 631 10226 659
rect 10192 625 10226 631
rect 10192 563 10226 587
rect 10192 553 10226 563
rect 10192 495 10226 515
rect 10192 481 10226 495
rect 10192 427 10226 443
rect 10192 409 10226 427
rect 10192 359 10226 371
rect 10192 337 10226 359
rect 10192 291 10226 299
rect 10192 265 10226 291
rect 10288 1209 10322 1235
rect 10288 1201 10322 1209
rect 10288 1141 10322 1163
rect 10288 1129 10322 1141
rect 10288 1073 10322 1091
rect 10288 1057 10322 1073
rect 10288 1005 10322 1019
rect 10288 985 10322 1005
rect 10288 937 10322 947
rect 10288 913 10322 937
rect 10288 869 10322 875
rect 10288 841 10322 869
rect 10288 801 10322 803
rect 10288 769 10322 801
rect 10288 699 10322 731
rect 10288 697 10322 699
rect 10288 631 10322 659
rect 10288 625 10322 631
rect 10288 563 10322 587
rect 10288 553 10322 563
rect 10288 495 10322 515
rect 10288 481 10322 495
rect 10288 427 10322 443
rect 10288 409 10322 427
rect 10288 359 10322 371
rect 10288 337 10322 359
rect 10288 291 10322 299
rect 10288 265 10322 291
rect 10384 1209 10418 1235
rect 10384 1201 10418 1209
rect 10384 1141 10418 1163
rect 10384 1129 10418 1141
rect 10384 1073 10418 1091
rect 10384 1057 10418 1073
rect 10384 1005 10418 1019
rect 10384 985 10418 1005
rect 10384 937 10418 947
rect 10384 913 10418 937
rect 10384 869 10418 875
rect 10384 841 10418 869
rect 10384 801 10418 803
rect 10384 769 10418 801
rect 10384 699 10418 731
rect 10384 697 10418 699
rect 10384 631 10418 659
rect 10384 625 10418 631
rect 10384 563 10418 587
rect 10384 553 10418 563
rect 10384 495 10418 515
rect 10384 481 10418 495
rect 10384 427 10418 443
rect 10384 409 10418 427
rect 10384 359 10418 371
rect 10384 337 10418 359
rect 10384 291 10418 299
rect 10384 265 10418 291
rect 8480 96 8514 130
rect 8774 80 8808 114
rect 9230 78 9264 112
rect 9904 68 9938 102
rect 7632 -16 7854 18
rect 15466 1458 15500 1492
rect 11474 1400 11508 1434
rect 12964 1380 12998 1414
rect 11000 1209 11034 1235
rect 11000 1201 11034 1209
rect 11000 1141 11034 1163
rect 11000 1129 11034 1141
rect 11000 1073 11034 1091
rect 11000 1057 11034 1073
rect 11000 1005 11034 1019
rect 11000 985 11034 1005
rect 11000 937 11034 947
rect 11000 913 11034 937
rect 11000 869 11034 875
rect 11000 841 11034 869
rect 11000 801 11034 803
rect 11000 769 11034 801
rect 11000 699 11034 731
rect 11000 697 11034 699
rect 11000 631 11034 659
rect 11000 625 11034 631
rect 11000 563 11034 587
rect 11000 553 11034 563
rect 11000 495 11034 515
rect 11000 481 11034 495
rect 11000 427 11034 443
rect 11000 409 11034 427
rect 11000 359 11034 371
rect 11000 337 11034 359
rect 11000 291 11034 299
rect 11000 265 11034 291
rect 11096 1209 11130 1235
rect 11096 1201 11130 1209
rect 11096 1141 11130 1163
rect 11096 1129 11130 1141
rect 11096 1073 11130 1091
rect 11096 1057 11130 1073
rect 11096 1005 11130 1019
rect 11096 985 11130 1005
rect 11096 937 11130 947
rect 11096 913 11130 937
rect 11096 869 11130 875
rect 11096 841 11130 869
rect 11096 801 11130 803
rect 11096 769 11130 801
rect 11096 699 11130 731
rect 11096 697 11130 699
rect 11096 631 11130 659
rect 11096 625 11130 631
rect 11096 563 11130 587
rect 11096 553 11130 563
rect 11096 495 11130 515
rect 11096 481 11130 495
rect 11096 427 11130 443
rect 11096 409 11130 427
rect 11096 359 11130 371
rect 11096 337 11130 359
rect 11096 291 11130 299
rect 11096 265 11130 291
rect 11192 1209 11226 1235
rect 11192 1201 11226 1209
rect 11192 1141 11226 1163
rect 11192 1129 11226 1141
rect 11192 1073 11226 1091
rect 11192 1057 11226 1073
rect 11192 1005 11226 1019
rect 11192 985 11226 1005
rect 11192 937 11226 947
rect 11192 913 11226 937
rect 11192 869 11226 875
rect 11192 841 11226 869
rect 11192 801 11226 803
rect 11192 769 11226 801
rect 11192 699 11226 731
rect 11192 697 11226 699
rect 11192 631 11226 659
rect 11192 625 11226 631
rect 11192 563 11226 587
rect 11192 553 11226 563
rect 11192 495 11226 515
rect 11192 481 11226 495
rect 11192 427 11226 443
rect 11192 409 11226 427
rect 11192 359 11226 371
rect 11192 337 11226 359
rect 11192 291 11226 299
rect 11192 265 11226 291
rect 11288 1209 11322 1235
rect 11288 1201 11322 1209
rect 11288 1141 11322 1163
rect 11288 1129 11322 1141
rect 11288 1073 11322 1091
rect 11288 1057 11322 1073
rect 11288 1005 11322 1019
rect 11288 985 11322 1005
rect 11288 937 11322 947
rect 11288 913 11322 937
rect 11288 869 11322 875
rect 11288 841 11322 869
rect 11288 801 11322 803
rect 11288 769 11322 801
rect 11288 699 11322 731
rect 11288 697 11322 699
rect 11288 631 11322 659
rect 11288 625 11322 631
rect 11288 563 11322 587
rect 11288 553 11322 563
rect 11288 495 11322 515
rect 11288 481 11322 495
rect 11288 427 11322 443
rect 11288 409 11322 427
rect 11288 359 11322 371
rect 11288 337 11322 359
rect 11288 291 11322 299
rect 11288 265 11322 291
rect 11384 1209 11418 1235
rect 11384 1201 11418 1209
rect 11384 1141 11418 1163
rect 11384 1129 11418 1141
rect 11384 1073 11418 1091
rect 11384 1057 11418 1073
rect 11384 1005 11418 1019
rect 11384 985 11418 1005
rect 11384 937 11418 947
rect 11384 913 11418 937
rect 11384 869 11418 875
rect 11384 841 11418 869
rect 11384 801 11418 803
rect 11384 769 11418 801
rect 11384 699 11418 731
rect 11384 697 11418 699
rect 11384 631 11418 659
rect 11384 625 11418 631
rect 11384 563 11418 587
rect 11384 553 11418 563
rect 11384 495 11418 515
rect 11384 481 11418 495
rect 11384 427 11418 443
rect 11384 409 11418 427
rect 11384 359 11418 371
rect 11384 337 11418 359
rect 11384 291 11418 299
rect 11384 265 11418 291
rect 11480 1209 11514 1235
rect 11480 1201 11514 1209
rect 11480 1141 11514 1163
rect 11480 1129 11514 1141
rect 11480 1073 11514 1091
rect 11480 1057 11514 1073
rect 11480 1005 11514 1019
rect 11480 985 11514 1005
rect 11480 937 11514 947
rect 11480 913 11514 937
rect 11480 869 11514 875
rect 11480 841 11514 869
rect 11480 801 11514 803
rect 11480 769 11514 801
rect 11480 699 11514 731
rect 11480 697 11514 699
rect 11480 631 11514 659
rect 11480 625 11514 631
rect 11480 563 11514 587
rect 11480 553 11514 563
rect 11480 495 11514 515
rect 11480 481 11514 495
rect 11480 427 11514 443
rect 11480 409 11514 427
rect 11480 359 11514 371
rect 11480 337 11514 359
rect 11480 291 11514 299
rect 11480 265 11514 291
rect 11576 1209 11610 1235
rect 11576 1201 11610 1209
rect 11576 1141 11610 1163
rect 11576 1129 11610 1141
rect 11576 1073 11610 1091
rect 11576 1057 11610 1073
rect 11576 1005 11610 1019
rect 11576 985 11610 1005
rect 11576 937 11610 947
rect 11576 913 11610 937
rect 11576 869 11610 875
rect 11576 841 11610 869
rect 11576 801 11610 803
rect 11576 769 11610 801
rect 11576 699 11610 731
rect 11576 697 11610 699
rect 11576 631 11610 659
rect 11576 625 11610 631
rect 11576 563 11610 587
rect 11576 553 11610 563
rect 11576 495 11610 515
rect 11576 481 11610 495
rect 11576 427 11610 443
rect 11576 409 11610 427
rect 11576 359 11610 371
rect 11576 337 11610 359
rect 11576 291 11610 299
rect 11576 265 11610 291
rect 11672 1209 11706 1235
rect 11672 1201 11706 1209
rect 11672 1141 11706 1163
rect 11672 1129 11706 1141
rect 11672 1073 11706 1091
rect 11672 1057 11706 1073
rect 11672 1005 11706 1019
rect 11672 985 11706 1005
rect 11672 937 11706 947
rect 11672 913 11706 937
rect 11672 869 11706 875
rect 11672 841 11706 869
rect 11672 801 11706 803
rect 11672 769 11706 801
rect 11672 699 11706 731
rect 11672 697 11706 699
rect 11672 631 11706 659
rect 11672 625 11706 631
rect 11672 563 11706 587
rect 11672 553 11706 563
rect 11672 495 11706 515
rect 11672 481 11706 495
rect 11672 427 11706 443
rect 11672 409 11706 427
rect 11672 359 11706 371
rect 11672 337 11706 359
rect 11672 291 11706 299
rect 11672 265 11706 291
rect 11768 1209 11802 1235
rect 11768 1201 11802 1209
rect 11768 1141 11802 1163
rect 11768 1129 11802 1141
rect 11768 1073 11802 1091
rect 11768 1057 11802 1073
rect 11768 1005 11802 1019
rect 11768 985 11802 1005
rect 11768 937 11802 947
rect 11768 913 11802 937
rect 11768 869 11802 875
rect 11768 841 11802 869
rect 11768 801 11802 803
rect 11768 769 11802 801
rect 11768 699 11802 731
rect 11768 697 11802 699
rect 11768 631 11802 659
rect 11768 625 11802 631
rect 11768 563 11802 587
rect 11768 553 11802 563
rect 11768 495 11802 515
rect 11768 481 11802 495
rect 11768 427 11802 443
rect 11768 409 11802 427
rect 11768 359 11802 371
rect 11768 337 11802 359
rect 11768 291 11802 299
rect 11768 265 11802 291
rect 11864 1209 11898 1235
rect 11864 1201 11898 1209
rect 11864 1141 11898 1163
rect 11864 1129 11898 1141
rect 11864 1073 11898 1091
rect 11864 1057 11898 1073
rect 11864 1005 11898 1019
rect 11864 985 11898 1005
rect 11864 937 11898 947
rect 11864 913 11898 937
rect 11864 869 11898 875
rect 11864 841 11898 869
rect 11864 801 11898 803
rect 11864 769 11898 801
rect 11864 699 11898 731
rect 11864 697 11898 699
rect 11864 631 11898 659
rect 11864 625 11898 631
rect 11864 563 11898 587
rect 11864 553 11898 563
rect 11864 495 11898 515
rect 11864 481 11898 495
rect 11864 427 11898 443
rect 11864 409 11898 427
rect 11864 359 11898 371
rect 11864 337 11898 359
rect 11864 291 11898 299
rect 11864 265 11898 291
rect 11960 1209 11994 1235
rect 11960 1201 11994 1209
rect 11960 1141 11994 1163
rect 11960 1129 11994 1141
rect 11960 1073 11994 1091
rect 11960 1057 11994 1073
rect 11960 1005 11994 1019
rect 11960 985 11994 1005
rect 11960 937 11994 947
rect 11960 913 11994 937
rect 11960 869 11994 875
rect 11960 841 11994 869
rect 11960 801 11994 803
rect 11960 769 11994 801
rect 11960 699 11994 731
rect 11960 697 11994 699
rect 11960 631 11994 659
rect 11960 625 11994 631
rect 11960 563 11994 587
rect 11960 553 11994 563
rect 11960 495 11994 515
rect 11960 481 11994 495
rect 11960 427 11994 443
rect 11960 409 11994 427
rect 11960 359 11994 371
rect 11960 337 11994 359
rect 11960 291 11994 299
rect 11960 265 11994 291
rect 12056 1209 12090 1235
rect 12056 1201 12090 1209
rect 12056 1141 12090 1163
rect 12056 1129 12090 1141
rect 12056 1073 12090 1091
rect 12056 1057 12090 1073
rect 12056 1005 12090 1019
rect 12056 985 12090 1005
rect 12056 937 12090 947
rect 12056 913 12090 937
rect 12056 869 12090 875
rect 12056 841 12090 869
rect 12056 801 12090 803
rect 12056 769 12090 801
rect 12056 699 12090 731
rect 12056 697 12090 699
rect 12056 631 12090 659
rect 12056 625 12090 631
rect 12056 563 12090 587
rect 12056 553 12090 563
rect 12056 495 12090 515
rect 12056 481 12090 495
rect 12056 427 12090 443
rect 12056 409 12090 427
rect 12056 359 12090 371
rect 12056 337 12090 359
rect 12056 291 12090 299
rect 12056 265 12090 291
rect 12388 1183 12422 1209
rect 12388 1175 12422 1183
rect 12388 1115 12422 1137
rect 12388 1103 12422 1115
rect 12388 1047 12422 1065
rect 12388 1031 12422 1047
rect 12388 979 12422 993
rect 12388 959 12422 979
rect 12388 911 12422 921
rect 12388 887 12422 911
rect 12388 843 12422 849
rect 12388 815 12422 843
rect 12388 775 12422 777
rect 12388 743 12422 775
rect 12388 673 12422 705
rect 12388 671 12422 673
rect 12388 605 12422 633
rect 12388 599 12422 605
rect 12388 537 12422 561
rect 12388 527 12422 537
rect 12388 469 12422 489
rect 12388 455 12422 469
rect 12388 401 12422 417
rect 12388 383 12422 401
rect 12388 333 12422 345
rect 12388 311 12422 333
rect 12388 265 12422 273
rect 12388 239 12422 265
rect 12484 1183 12518 1209
rect 12484 1175 12518 1183
rect 12484 1115 12518 1137
rect 12484 1103 12518 1115
rect 12484 1047 12518 1065
rect 12484 1031 12518 1047
rect 12484 979 12518 993
rect 12484 959 12518 979
rect 12484 911 12518 921
rect 12484 887 12518 911
rect 12484 843 12518 849
rect 12484 815 12518 843
rect 12484 775 12518 777
rect 12484 743 12518 775
rect 12484 673 12518 705
rect 12484 671 12518 673
rect 12484 605 12518 633
rect 12484 599 12518 605
rect 12484 537 12518 561
rect 12484 527 12518 537
rect 12484 469 12518 489
rect 12484 455 12518 469
rect 12484 401 12518 417
rect 12484 383 12518 401
rect 12484 333 12518 345
rect 12484 311 12518 333
rect 12484 265 12518 273
rect 12484 239 12518 265
rect 12580 1183 12614 1209
rect 12580 1175 12614 1183
rect 12580 1115 12614 1137
rect 12580 1103 12614 1115
rect 12580 1047 12614 1065
rect 12580 1031 12614 1047
rect 12580 979 12614 993
rect 12580 959 12614 979
rect 12580 911 12614 921
rect 12580 887 12614 911
rect 12580 843 12614 849
rect 12580 815 12614 843
rect 12580 775 12614 777
rect 12580 743 12614 775
rect 12580 673 12614 705
rect 12580 671 12614 673
rect 12580 605 12614 633
rect 12580 599 12614 605
rect 12580 537 12614 561
rect 12580 527 12614 537
rect 12580 469 12614 489
rect 12580 455 12614 469
rect 12580 401 12614 417
rect 12580 383 12614 401
rect 12580 333 12614 345
rect 12580 311 12614 333
rect 12580 265 12614 273
rect 12580 239 12614 265
rect 12676 1183 12710 1209
rect 12676 1175 12710 1183
rect 12676 1115 12710 1137
rect 12676 1103 12710 1115
rect 12676 1047 12710 1065
rect 12676 1031 12710 1047
rect 12676 979 12710 993
rect 12676 959 12710 979
rect 12676 911 12710 921
rect 12676 887 12710 911
rect 12676 843 12710 849
rect 12676 815 12710 843
rect 12676 775 12710 777
rect 12676 743 12710 775
rect 12676 673 12710 705
rect 12676 671 12710 673
rect 12676 605 12710 633
rect 12676 599 12710 605
rect 12676 537 12710 561
rect 12676 527 12710 537
rect 12676 469 12710 489
rect 12676 455 12710 469
rect 12676 401 12710 417
rect 12676 383 12710 401
rect 12676 333 12710 345
rect 12676 311 12710 333
rect 12676 265 12710 273
rect 12676 239 12710 265
rect 12772 1183 12806 1209
rect 12772 1175 12806 1183
rect 12772 1115 12806 1137
rect 12772 1103 12806 1115
rect 12772 1047 12806 1065
rect 12772 1031 12806 1047
rect 12772 979 12806 993
rect 12772 959 12806 979
rect 12772 911 12806 921
rect 12772 887 12806 911
rect 12772 843 12806 849
rect 12772 815 12806 843
rect 12772 775 12806 777
rect 12772 743 12806 775
rect 12772 673 12806 705
rect 12772 671 12806 673
rect 12772 605 12806 633
rect 12772 599 12806 605
rect 12772 537 12806 561
rect 12772 527 12806 537
rect 12772 469 12806 489
rect 12772 455 12806 469
rect 12772 401 12806 417
rect 12772 383 12806 401
rect 12772 333 12806 345
rect 12772 311 12806 333
rect 12772 265 12806 273
rect 12772 239 12806 265
rect 12868 1183 12902 1209
rect 12868 1175 12902 1183
rect 12868 1115 12902 1137
rect 12868 1103 12902 1115
rect 12868 1047 12902 1065
rect 12868 1031 12902 1047
rect 12868 979 12902 993
rect 12868 959 12902 979
rect 12868 911 12902 921
rect 12868 887 12902 911
rect 12868 843 12902 849
rect 12868 815 12902 843
rect 12868 775 12902 777
rect 12868 743 12902 775
rect 12868 673 12902 705
rect 12868 671 12902 673
rect 12868 605 12902 633
rect 12868 599 12902 605
rect 12868 537 12902 561
rect 12868 527 12902 537
rect 12868 469 12902 489
rect 12868 455 12902 469
rect 12868 401 12902 417
rect 12868 383 12902 401
rect 12868 333 12902 345
rect 12868 311 12902 333
rect 12868 265 12902 273
rect 12868 239 12902 265
rect 12964 1183 12998 1209
rect 12964 1175 12998 1183
rect 12964 1115 12998 1137
rect 12964 1103 12998 1115
rect 12964 1047 12998 1065
rect 12964 1031 12998 1047
rect 12964 979 12998 993
rect 12964 959 12998 979
rect 12964 911 12998 921
rect 12964 887 12998 911
rect 12964 843 12998 849
rect 12964 815 12998 843
rect 12964 775 12998 777
rect 12964 743 12998 775
rect 12964 673 12998 705
rect 12964 671 12998 673
rect 12964 605 12998 633
rect 12964 599 12998 605
rect 12964 537 12998 561
rect 12964 527 12998 537
rect 12964 469 12998 489
rect 12964 455 12998 469
rect 12964 401 12998 417
rect 12964 383 12998 401
rect 12964 333 12998 345
rect 12964 311 12998 333
rect 12964 265 12998 273
rect 12964 239 12998 265
rect 13060 1183 13094 1209
rect 13060 1175 13094 1183
rect 13060 1115 13094 1137
rect 13060 1103 13094 1115
rect 13060 1047 13094 1065
rect 13060 1031 13094 1047
rect 13060 979 13094 993
rect 13060 959 13094 979
rect 13060 911 13094 921
rect 13060 887 13094 911
rect 13060 843 13094 849
rect 13060 815 13094 843
rect 13060 775 13094 777
rect 13060 743 13094 775
rect 13060 673 13094 705
rect 13060 671 13094 673
rect 13060 605 13094 633
rect 13060 599 13094 605
rect 13060 537 13094 561
rect 13060 527 13094 537
rect 13060 469 13094 489
rect 13060 455 13094 469
rect 13060 401 13094 417
rect 13060 383 13094 401
rect 13060 333 13094 345
rect 13060 311 13094 333
rect 13060 265 13094 273
rect 13060 239 13094 265
rect 13156 1183 13190 1209
rect 13156 1175 13190 1183
rect 13156 1115 13190 1137
rect 13156 1103 13190 1115
rect 13156 1047 13190 1065
rect 13156 1031 13190 1047
rect 13156 979 13190 993
rect 13156 959 13190 979
rect 13156 911 13190 921
rect 13156 887 13190 911
rect 13156 843 13190 849
rect 13156 815 13190 843
rect 13156 775 13190 777
rect 13156 743 13190 775
rect 13156 673 13190 705
rect 13156 671 13190 673
rect 13156 605 13190 633
rect 13156 599 13190 605
rect 13156 537 13190 561
rect 13156 527 13190 537
rect 13156 469 13190 489
rect 13156 455 13190 469
rect 13156 401 13190 417
rect 13156 383 13190 401
rect 13156 333 13190 345
rect 13156 311 13190 333
rect 13156 265 13190 273
rect 13156 239 13190 265
rect 13252 1183 13286 1209
rect 13252 1175 13286 1183
rect 13252 1115 13286 1137
rect 13252 1103 13286 1115
rect 13252 1047 13286 1065
rect 13252 1031 13286 1047
rect 13252 979 13286 993
rect 13252 959 13286 979
rect 13252 911 13286 921
rect 13252 887 13286 911
rect 13252 843 13286 849
rect 13252 815 13286 843
rect 13252 775 13286 777
rect 13252 743 13286 775
rect 13252 673 13286 705
rect 13252 671 13286 673
rect 13252 605 13286 633
rect 13252 599 13286 605
rect 13252 537 13286 561
rect 13252 527 13286 537
rect 13252 469 13286 489
rect 13252 455 13286 469
rect 13252 401 13286 417
rect 13252 383 13286 401
rect 13252 333 13286 345
rect 13252 311 13286 333
rect 13252 265 13286 273
rect 13252 239 13286 265
rect 13348 1183 13382 1209
rect 13348 1175 13382 1183
rect 13348 1115 13382 1137
rect 13348 1103 13382 1115
rect 13348 1047 13382 1065
rect 13348 1031 13382 1047
rect 13348 979 13382 993
rect 13348 959 13382 979
rect 13348 911 13382 921
rect 13348 887 13382 911
rect 13348 843 13382 849
rect 13348 815 13382 843
rect 13348 775 13382 777
rect 13348 743 13382 775
rect 13348 673 13382 705
rect 13348 671 13382 673
rect 13348 605 13382 633
rect 13348 599 13382 605
rect 13348 537 13382 561
rect 13348 527 13382 537
rect 13348 469 13382 489
rect 13348 455 13382 469
rect 13348 401 13382 417
rect 13348 383 13382 401
rect 13348 333 13382 345
rect 13348 311 13382 333
rect 13348 265 13382 273
rect 13348 239 13382 265
rect 13444 1183 13478 1209
rect 13444 1175 13478 1183
rect 13444 1115 13478 1137
rect 13444 1103 13478 1115
rect 13444 1047 13478 1065
rect 13444 1031 13478 1047
rect 13444 979 13478 993
rect 13444 959 13478 979
rect 13444 911 13478 921
rect 13444 887 13478 911
rect 13444 843 13478 849
rect 13444 815 13478 843
rect 13444 775 13478 777
rect 13444 743 13478 775
rect 13444 673 13478 705
rect 13444 671 13478 673
rect 13444 605 13478 633
rect 13444 599 13478 605
rect 13444 537 13478 561
rect 13444 527 13478 537
rect 13444 469 13478 489
rect 13444 455 13478 469
rect 13444 401 13478 417
rect 13444 383 13478 401
rect 13444 333 13478 345
rect 13444 311 13478 333
rect 13444 265 13478 273
rect 13444 239 13478 265
rect 13540 1183 13574 1209
rect 13540 1175 13574 1183
rect 13540 1115 13574 1137
rect 13540 1103 13574 1115
rect 13540 1047 13574 1065
rect 13540 1031 13574 1047
rect 13540 979 13574 993
rect 13540 959 13574 979
rect 13540 911 13574 921
rect 13540 887 13574 911
rect 13540 843 13574 849
rect 13540 815 13574 843
rect 13540 775 13574 777
rect 13540 743 13574 775
rect 13540 673 13574 705
rect 13540 671 13574 673
rect 13540 605 13574 633
rect 13540 599 13574 605
rect 13540 537 13574 561
rect 13540 527 13574 537
rect 13540 469 13574 489
rect 13540 455 13574 469
rect 13540 401 13574 417
rect 13540 383 13574 401
rect 13540 333 13574 345
rect 13540 311 13574 333
rect 13540 265 13574 273
rect 13540 239 13574 265
rect 11568 94 11602 128
rect 11862 78 11896 112
rect 12386 52 12420 86
rect 13060 42 13094 76
rect 10562 -24 10796 12
rect 14630 1374 14664 1408
rect 15422 1336 15456 1370
rect 14156 1183 14190 1209
rect 14156 1175 14190 1183
rect 14156 1115 14190 1137
rect 14156 1103 14190 1115
rect 14156 1047 14190 1065
rect 14156 1031 14190 1047
rect 14156 979 14190 993
rect 14156 959 14190 979
rect 14156 911 14190 921
rect 14156 887 14190 911
rect 14156 843 14190 849
rect 14156 815 14190 843
rect 14156 775 14190 777
rect 14156 743 14190 775
rect 14156 673 14190 705
rect 14156 671 14190 673
rect 14156 605 14190 633
rect 14156 599 14190 605
rect 14156 537 14190 561
rect 14156 527 14190 537
rect 14156 469 14190 489
rect 14156 455 14190 469
rect 14156 401 14190 417
rect 14156 383 14190 401
rect 14156 333 14190 345
rect 14156 311 14190 333
rect 14156 265 14190 273
rect 14156 239 14190 265
rect 14252 1183 14286 1209
rect 14252 1175 14286 1183
rect 14252 1115 14286 1137
rect 14252 1103 14286 1115
rect 14252 1047 14286 1065
rect 14252 1031 14286 1047
rect 14252 979 14286 993
rect 14252 959 14286 979
rect 14252 911 14286 921
rect 14252 887 14286 911
rect 14252 843 14286 849
rect 14252 815 14286 843
rect 14252 775 14286 777
rect 14252 743 14286 775
rect 14252 673 14286 705
rect 14252 671 14286 673
rect 14252 605 14286 633
rect 14252 599 14286 605
rect 14252 537 14286 561
rect 14252 527 14286 537
rect 14252 469 14286 489
rect 14252 455 14286 469
rect 14252 401 14286 417
rect 14252 383 14286 401
rect 14252 333 14286 345
rect 14252 311 14286 333
rect 14252 265 14286 273
rect 14252 239 14286 265
rect 14348 1183 14382 1209
rect 14348 1175 14382 1183
rect 14348 1115 14382 1137
rect 14348 1103 14382 1115
rect 14348 1047 14382 1065
rect 14348 1031 14382 1047
rect 14348 979 14382 993
rect 14348 959 14382 979
rect 14348 911 14382 921
rect 14348 887 14382 911
rect 14348 843 14382 849
rect 14348 815 14382 843
rect 14348 775 14382 777
rect 14348 743 14382 775
rect 14348 673 14382 705
rect 14348 671 14382 673
rect 14348 605 14382 633
rect 14348 599 14382 605
rect 14348 537 14382 561
rect 14348 527 14382 537
rect 14348 469 14382 489
rect 14348 455 14382 469
rect 14348 401 14382 417
rect 14348 383 14382 401
rect 14348 333 14382 345
rect 14348 311 14382 333
rect 14348 265 14382 273
rect 14348 239 14382 265
rect 14444 1183 14478 1209
rect 14444 1175 14478 1183
rect 14444 1115 14478 1137
rect 14444 1103 14478 1115
rect 14444 1047 14478 1065
rect 14444 1031 14478 1047
rect 14444 979 14478 993
rect 14444 959 14478 979
rect 14444 911 14478 921
rect 14444 887 14478 911
rect 14444 843 14478 849
rect 14444 815 14478 843
rect 14444 775 14478 777
rect 14444 743 14478 775
rect 14444 673 14478 705
rect 14444 671 14478 673
rect 14444 605 14478 633
rect 14444 599 14478 605
rect 14444 537 14478 561
rect 14444 527 14478 537
rect 14444 469 14478 489
rect 14444 455 14478 469
rect 14444 401 14478 417
rect 14444 383 14478 401
rect 14444 333 14478 345
rect 14444 311 14478 333
rect 14444 265 14478 273
rect 14444 239 14478 265
rect 14540 1183 14574 1209
rect 14540 1175 14574 1183
rect 14540 1115 14574 1137
rect 14540 1103 14574 1115
rect 14540 1047 14574 1065
rect 14540 1031 14574 1047
rect 14540 979 14574 993
rect 14540 959 14574 979
rect 14540 911 14574 921
rect 14540 887 14574 911
rect 14540 843 14574 849
rect 14540 815 14574 843
rect 14540 775 14574 777
rect 14540 743 14574 775
rect 14540 673 14574 705
rect 14540 671 14574 673
rect 14540 605 14574 633
rect 14540 599 14574 605
rect 14540 537 14574 561
rect 14540 527 14574 537
rect 14540 469 14574 489
rect 14540 455 14574 469
rect 14540 401 14574 417
rect 14540 383 14574 401
rect 14540 333 14574 345
rect 14540 311 14574 333
rect 14540 265 14574 273
rect 14540 239 14574 265
rect 14636 1183 14670 1209
rect 14636 1175 14670 1183
rect 14636 1115 14670 1137
rect 14636 1103 14670 1115
rect 14636 1047 14670 1065
rect 14636 1031 14670 1047
rect 14636 979 14670 993
rect 14636 959 14670 979
rect 14636 911 14670 921
rect 14636 887 14670 911
rect 14636 843 14670 849
rect 14636 815 14670 843
rect 14636 775 14670 777
rect 14636 743 14670 775
rect 14636 673 14670 705
rect 14636 671 14670 673
rect 14636 605 14670 633
rect 14636 599 14670 605
rect 14636 537 14670 561
rect 14636 527 14670 537
rect 14636 469 14670 489
rect 14636 455 14670 469
rect 14636 401 14670 417
rect 14636 383 14670 401
rect 14636 333 14670 345
rect 14636 311 14670 333
rect 14636 265 14670 273
rect 14636 239 14670 265
rect 14732 1183 14766 1209
rect 14732 1175 14766 1183
rect 14732 1115 14766 1137
rect 14732 1103 14766 1115
rect 14732 1047 14766 1065
rect 14732 1031 14766 1047
rect 14732 979 14766 993
rect 14732 959 14766 979
rect 14732 911 14766 921
rect 14732 887 14766 911
rect 14732 843 14766 849
rect 14732 815 14766 843
rect 14732 775 14766 777
rect 14732 743 14766 775
rect 14732 673 14766 705
rect 14732 671 14766 673
rect 14732 605 14766 633
rect 14732 599 14766 605
rect 14732 537 14766 561
rect 14732 527 14766 537
rect 14732 469 14766 489
rect 14732 455 14766 469
rect 14732 401 14766 417
rect 14732 383 14766 401
rect 14732 333 14766 345
rect 14732 311 14766 333
rect 14732 265 14766 273
rect 14732 239 14766 265
rect 14828 1183 14862 1209
rect 14828 1175 14862 1183
rect 14828 1115 14862 1137
rect 14828 1103 14862 1115
rect 14828 1047 14862 1065
rect 14828 1031 14862 1047
rect 14828 979 14862 993
rect 14828 959 14862 979
rect 14828 911 14862 921
rect 14828 887 14862 911
rect 14828 843 14862 849
rect 14828 815 14862 843
rect 14828 775 14862 777
rect 14828 743 14862 775
rect 14828 673 14862 705
rect 14828 671 14862 673
rect 14828 605 14862 633
rect 14828 599 14862 605
rect 14828 537 14862 561
rect 14828 527 14862 537
rect 14828 469 14862 489
rect 14828 455 14862 469
rect 14828 401 14862 417
rect 14828 383 14862 401
rect 14828 333 14862 345
rect 14828 311 14862 333
rect 14828 265 14862 273
rect 14828 239 14862 265
rect 14924 1183 14958 1209
rect 14924 1175 14958 1183
rect 14924 1115 14958 1137
rect 14924 1103 14958 1115
rect 14924 1047 14958 1065
rect 14924 1031 14958 1047
rect 14924 979 14958 993
rect 14924 959 14958 979
rect 14924 911 14958 921
rect 14924 887 14958 911
rect 14924 843 14958 849
rect 14924 815 14958 843
rect 14924 775 14958 777
rect 14924 743 14958 775
rect 14924 673 14958 705
rect 14924 671 14958 673
rect 14924 605 14958 633
rect 14924 599 14958 605
rect 14924 537 14958 561
rect 14924 527 14958 537
rect 14924 469 14958 489
rect 14924 455 14958 469
rect 14924 401 14958 417
rect 14924 383 14958 401
rect 14924 333 14958 345
rect 14924 311 14958 333
rect 14924 265 14958 273
rect 14924 239 14958 265
rect 15020 1183 15054 1209
rect 15020 1175 15054 1183
rect 15020 1115 15054 1137
rect 15020 1103 15054 1115
rect 15020 1047 15054 1065
rect 15020 1031 15054 1047
rect 15020 979 15054 993
rect 15020 959 15054 979
rect 15020 911 15054 921
rect 15020 887 15054 911
rect 15020 843 15054 849
rect 15020 815 15054 843
rect 15020 775 15054 777
rect 15020 743 15054 775
rect 15020 673 15054 705
rect 15020 671 15054 673
rect 15020 605 15054 633
rect 15020 599 15054 605
rect 15020 537 15054 561
rect 15020 527 15054 537
rect 15020 469 15054 489
rect 15020 455 15054 469
rect 15020 401 15054 417
rect 15020 383 15054 401
rect 15020 333 15054 345
rect 15020 311 15054 333
rect 15020 265 15054 273
rect 15020 239 15054 265
rect 15116 1183 15150 1209
rect 15116 1175 15150 1183
rect 15116 1115 15150 1137
rect 15116 1103 15150 1115
rect 15116 1047 15150 1065
rect 15116 1031 15150 1047
rect 15116 979 15150 993
rect 15116 959 15150 979
rect 15116 911 15150 921
rect 15116 887 15150 911
rect 15116 843 15150 849
rect 15116 815 15150 843
rect 15116 775 15150 777
rect 15116 743 15150 775
rect 15116 673 15150 705
rect 15116 671 15150 673
rect 15116 605 15150 633
rect 15116 599 15150 605
rect 15116 537 15150 561
rect 15116 527 15150 537
rect 15116 469 15150 489
rect 15116 455 15150 469
rect 15116 401 15150 417
rect 15116 383 15150 401
rect 15116 333 15150 345
rect 15116 311 15150 333
rect 15116 265 15150 273
rect 15116 239 15150 265
rect 15212 1183 15246 1209
rect 15212 1175 15246 1183
rect 15212 1115 15246 1137
rect 15212 1103 15246 1115
rect 15212 1047 15246 1065
rect 15212 1031 15246 1047
rect 15212 979 15246 993
rect 15212 959 15246 979
rect 15212 911 15246 921
rect 15212 887 15246 911
rect 15212 843 15246 849
rect 15212 815 15246 843
rect 15212 775 15246 777
rect 15212 743 15246 775
rect 15212 673 15246 705
rect 15212 671 15246 673
rect 15212 605 15246 633
rect 15212 599 15246 605
rect 15212 537 15246 561
rect 15212 527 15246 537
rect 15212 469 15246 489
rect 15212 455 15246 469
rect 15212 401 15246 417
rect 15212 383 15246 401
rect 15212 333 15246 345
rect 15212 311 15246 333
rect 15212 265 15246 273
rect 15212 239 15246 265
rect 15422 1227 15456 1257
rect 15422 1223 15456 1227
rect 15422 1159 15456 1185
rect 15422 1151 15456 1159
rect 15422 1091 15456 1113
rect 15422 1079 15456 1091
rect 15422 1023 15456 1041
rect 15422 1007 15456 1023
rect 15422 955 15456 969
rect 15422 935 15456 955
rect 15422 887 15456 897
rect 15422 863 15456 887
rect 15422 819 15456 825
rect 15422 791 15456 819
rect 15422 751 15456 753
rect 15422 719 15456 751
rect 15422 649 15456 681
rect 15422 647 15456 649
rect 15422 581 15456 609
rect 15422 575 15456 581
rect 15422 513 15456 537
rect 15422 503 15456 513
rect 15422 445 15456 465
rect 15422 431 15456 445
rect 15422 377 15456 393
rect 15422 359 15456 377
rect 15422 309 15456 321
rect 15422 287 15456 309
rect 15422 241 15456 249
rect 15422 215 15456 241
rect 15422 173 15456 177
rect 15422 143 15456 173
rect 14724 68 14758 102
rect 15510 1227 15544 1257
rect 15510 1223 15544 1227
rect 15510 1159 15544 1185
rect 15510 1151 15544 1159
rect 15510 1091 15544 1113
rect 15510 1079 15544 1091
rect 15510 1023 15544 1041
rect 15510 1007 15544 1023
rect 15510 955 15544 969
rect 15510 935 15544 955
rect 15510 887 15544 897
rect 15510 863 15544 887
rect 15510 819 15544 825
rect 15510 791 15544 819
rect 15510 751 15544 753
rect 15510 719 15544 751
rect 15510 649 15544 681
rect 15510 647 15544 649
rect 15510 581 15544 609
rect 15510 575 15544 581
rect 15510 513 15544 537
rect 15510 503 15544 513
rect 15510 445 15544 465
rect 15510 431 15544 445
rect 15510 377 15544 393
rect 15510 359 15544 377
rect 15510 309 15544 321
rect 15510 287 15544 309
rect 15510 241 15544 249
rect 15510 215 15544 241
rect 15510 173 15544 177
rect 15510 143 15544 173
rect 15018 52 15052 86
rect 15510 18 15544 52
rect 13856 -50 14090 -14
rect 346 -1216 596 -1038
rect 15498 -1197 15676 -1019
rect 2269 -1643 2447 -1465
rect 4269 -1643 4447 -1465
rect 6269 -1643 6447 -1465
rect 8493 -1660 8671 -1482
rect 10269 -1643 10447 -1465
rect 12269 -1643 12447 -1465
rect 14269 -1643 14447 -1465
<< metal1 >>
rect -392 9061 -112 9074
rect -392 8817 -374 9061
rect -130 8817 -112 9061
rect -392 8804 -112 8817
rect 1608 9061 1888 9074
rect 1608 8817 1626 9061
rect 1870 8817 1888 9061
rect 1608 8804 1888 8817
rect 3608 9061 3888 9074
rect 3608 8817 3626 9061
rect 3870 8817 3888 9061
rect 3608 8804 3888 8817
rect 5608 9061 5888 9074
rect 5608 8817 5626 9061
rect 5870 8817 5888 9061
rect 5608 8804 5888 8817
rect 7608 9061 7888 9074
rect 7608 8817 7626 9061
rect 7870 8817 7888 9061
rect 7608 8804 7888 8817
rect 9608 9061 9888 9074
rect 9608 8817 9626 9061
rect 9870 8817 9888 9061
rect 9608 8804 9888 8817
rect 11608 9061 11888 9074
rect 11608 8817 11626 9061
rect 11870 8817 11888 9061
rect 11608 8804 11888 8817
rect 13608 9061 13888 9074
rect 13608 8817 13626 9061
rect 13870 8817 13888 9061
rect 15404 9066 15682 9090
rect 15404 8886 15421 9066
rect 15665 8886 15682 9066
rect 15404 8879 15454 8886
rect 15632 8879 15682 8886
rect 15404 8862 15682 8879
rect 13608 8804 13888 8817
rect -1360 8166 -762 8182
rect -1360 7858 -1343 8166
rect -779 7858 -762 8166
rect -1360 7842 -762 7858
rect 15394 8159 15832 8178
rect 15394 7851 15427 8159
rect 15799 7851 15832 8159
rect 15394 7832 15832 7851
rect -558 6998 12598 7210
rect -1658 5921 -1612 5936
rect -1658 5887 -1652 5921
rect -1618 5887 -1612 5921
rect -1658 5849 -1612 5887
rect -1658 5815 -1652 5849
rect -1618 5815 -1612 5849
rect -1658 5777 -1612 5815
rect -1658 5743 -1652 5777
rect -1618 5743 -1612 5777
rect -1658 5705 -1612 5743
rect -1658 5671 -1652 5705
rect -1618 5671 -1612 5705
rect -1658 5633 -1612 5671
rect -1658 5599 -1652 5633
rect -1618 5599 -1612 5633
rect -1658 5561 -1612 5599
rect -1658 5527 -1652 5561
rect -1618 5527 -1612 5561
rect -1658 5489 -1612 5527
rect -1658 5455 -1652 5489
rect -1618 5455 -1612 5489
rect -1658 5417 -1612 5455
rect -1658 5383 -1652 5417
rect -1618 5383 -1612 5417
rect -1658 5345 -1612 5383
rect -1658 5311 -1652 5345
rect -1618 5311 -1612 5345
rect -1658 5273 -1612 5311
rect -1658 5239 -1652 5273
rect -1618 5239 -1612 5273
rect -1658 5201 -1612 5239
rect -1658 5167 -1652 5201
rect -1618 5167 -1612 5201
rect -1658 5129 -1612 5167
rect -1658 5095 -1652 5129
rect -1618 5095 -1612 5129
rect -1658 5057 -1612 5095
rect -1658 5023 -1652 5057
rect -1618 5023 -1612 5057
rect -1658 4985 -1612 5023
rect -1658 4951 -1652 4985
rect -1618 4951 -1612 4985
rect -1658 4936 -1612 4951
rect -1560 5921 -1514 5936
rect -1560 5887 -1554 5921
rect -1520 5887 -1514 5921
rect -1560 5849 -1514 5887
rect -1560 5815 -1554 5849
rect -1520 5815 -1514 5849
rect -1560 5777 -1514 5815
rect -1560 5743 -1554 5777
rect -1520 5743 -1514 5777
rect -1560 5705 -1514 5743
rect -1560 5671 -1554 5705
rect -1520 5671 -1514 5705
rect -1560 5633 -1514 5671
rect -1560 5599 -1554 5633
rect -1520 5599 -1514 5633
rect -1560 5561 -1514 5599
rect -1560 5527 -1554 5561
rect -1520 5527 -1514 5561
rect -1560 5489 -1514 5527
rect -1560 5455 -1554 5489
rect -1520 5455 -1514 5489
rect -1560 5417 -1514 5455
rect -1560 5383 -1554 5417
rect -1520 5383 -1514 5417
rect -1560 5345 -1514 5383
rect -1560 5311 -1554 5345
rect -1520 5311 -1514 5345
rect -1560 5273 -1514 5311
rect -1560 5239 -1554 5273
rect -1520 5239 -1514 5273
rect -1560 5201 -1514 5239
rect -1560 5167 -1554 5201
rect -1520 5167 -1514 5201
rect -1560 5129 -1514 5167
rect -1560 5095 -1554 5129
rect -1520 5095 -1514 5129
rect -1560 5057 -1514 5095
rect -1560 5023 -1554 5057
rect -1520 5023 -1514 5057
rect -1560 4985 -1514 5023
rect -1560 4951 -1554 4985
rect -1520 4951 -1514 4985
rect -1560 4936 -1514 4951
rect -1462 5921 -1416 5936
rect -1462 5887 -1456 5921
rect -1422 5887 -1416 5921
rect -1462 5849 -1416 5887
rect -1462 5815 -1456 5849
rect -1422 5815 -1416 5849
rect -1462 5777 -1416 5815
rect -1462 5743 -1456 5777
rect -1422 5743 -1416 5777
rect -1462 5705 -1416 5743
rect -1462 5671 -1456 5705
rect -1422 5671 -1416 5705
rect -1462 5633 -1416 5671
rect -1462 5599 -1456 5633
rect -1422 5599 -1416 5633
rect -1462 5561 -1416 5599
rect -1462 5527 -1456 5561
rect -1422 5527 -1416 5561
rect -1462 5489 -1416 5527
rect -1462 5455 -1456 5489
rect -1422 5455 -1416 5489
rect -1462 5417 -1416 5455
rect -1462 5383 -1456 5417
rect -1422 5383 -1416 5417
rect -1462 5345 -1416 5383
rect -1462 5311 -1456 5345
rect -1422 5311 -1416 5345
rect -1462 5273 -1416 5311
rect -1462 5239 -1456 5273
rect -1422 5239 -1416 5273
rect -1462 5201 -1416 5239
rect -1462 5167 -1456 5201
rect -1422 5167 -1416 5201
rect -1462 5129 -1416 5167
rect -1462 5095 -1456 5129
rect -1422 5095 -1416 5129
rect -1462 5057 -1416 5095
rect -1462 5023 -1456 5057
rect -1422 5023 -1416 5057
rect -1462 4985 -1416 5023
rect -1462 4951 -1456 4985
rect -1422 4951 -1416 4985
rect -1462 4936 -1416 4951
rect -1364 5921 -1318 5936
rect -1364 5887 -1358 5921
rect -1324 5887 -1318 5921
rect -1364 5849 -1318 5887
rect -1364 5815 -1358 5849
rect -1324 5815 -1318 5849
rect -1364 5777 -1318 5815
rect -1364 5743 -1358 5777
rect -1324 5743 -1318 5777
rect -1364 5705 -1318 5743
rect -1364 5671 -1358 5705
rect -1324 5671 -1318 5705
rect -1364 5633 -1318 5671
rect -1364 5599 -1358 5633
rect -1324 5599 -1318 5633
rect -1364 5561 -1318 5599
rect -1364 5527 -1358 5561
rect -1324 5527 -1318 5561
rect -1364 5489 -1318 5527
rect -1364 5455 -1358 5489
rect -1324 5455 -1318 5489
rect -1364 5417 -1318 5455
rect -1364 5383 -1358 5417
rect -1324 5383 -1318 5417
rect -1364 5345 -1318 5383
rect -1364 5311 -1358 5345
rect -1324 5311 -1318 5345
rect -1364 5273 -1318 5311
rect -1364 5239 -1358 5273
rect -1324 5239 -1318 5273
rect -1364 5201 -1318 5239
rect -1364 5167 -1358 5201
rect -1324 5167 -1318 5201
rect -1364 5129 -1318 5167
rect -1364 5095 -1358 5129
rect -1324 5095 -1318 5129
rect -1364 5057 -1318 5095
rect -1364 5023 -1358 5057
rect -1324 5023 -1318 5057
rect -1364 4985 -1318 5023
rect -1364 4951 -1358 4985
rect -1324 4951 -1318 4985
rect -1364 4936 -1318 4951
rect -1266 5921 -1220 5936
rect -1266 5887 -1260 5921
rect -1226 5887 -1220 5921
rect -1266 5849 -1220 5887
rect -1266 5815 -1260 5849
rect -1226 5815 -1220 5849
rect -1266 5777 -1220 5815
rect -1266 5743 -1260 5777
rect -1226 5743 -1220 5777
rect -1266 5705 -1220 5743
rect -1266 5671 -1260 5705
rect -1226 5671 -1220 5705
rect -1266 5633 -1220 5671
rect -1266 5599 -1260 5633
rect -1226 5599 -1220 5633
rect -1266 5561 -1220 5599
rect -1266 5527 -1260 5561
rect -1226 5527 -1220 5561
rect -1266 5489 -1220 5527
rect -1266 5455 -1260 5489
rect -1226 5455 -1220 5489
rect -1266 5417 -1220 5455
rect -1266 5383 -1260 5417
rect -1226 5383 -1220 5417
rect -1266 5345 -1220 5383
rect -1266 5311 -1260 5345
rect -1226 5311 -1220 5345
rect -1266 5273 -1220 5311
rect -1266 5239 -1260 5273
rect -1226 5239 -1220 5273
rect -1266 5201 -1220 5239
rect -1266 5167 -1260 5201
rect -1226 5167 -1220 5201
rect -1266 5129 -1220 5167
rect -1266 5095 -1260 5129
rect -1226 5095 -1220 5129
rect -1266 5057 -1220 5095
rect -1266 5023 -1260 5057
rect -1226 5023 -1220 5057
rect -1266 4985 -1220 5023
rect -1266 4951 -1260 4985
rect -1226 4951 -1220 4985
rect -1266 4936 -1220 4951
rect -1168 5921 -1122 5936
rect -1168 5887 -1162 5921
rect -1128 5887 -1122 5921
rect -1168 5849 -1122 5887
rect -1168 5815 -1162 5849
rect -1128 5815 -1122 5849
rect -1168 5777 -1122 5815
rect -1168 5743 -1162 5777
rect -1128 5743 -1122 5777
rect -1168 5705 -1122 5743
rect -1168 5671 -1162 5705
rect -1128 5671 -1122 5705
rect -1168 5633 -1122 5671
rect -1168 5599 -1162 5633
rect -1128 5599 -1122 5633
rect -1168 5561 -1122 5599
rect -1168 5527 -1162 5561
rect -1128 5527 -1122 5561
rect -1168 5489 -1122 5527
rect -1168 5455 -1162 5489
rect -1128 5455 -1122 5489
rect -1168 5417 -1122 5455
rect -1168 5383 -1162 5417
rect -1128 5383 -1122 5417
rect -1168 5345 -1122 5383
rect -1168 5311 -1162 5345
rect -1128 5311 -1122 5345
rect -1168 5273 -1122 5311
rect -1168 5239 -1162 5273
rect -1128 5239 -1122 5273
rect -1168 5201 -1122 5239
rect -1168 5167 -1162 5201
rect -1128 5167 -1122 5201
rect -1168 5129 -1122 5167
rect -1168 5095 -1162 5129
rect -1128 5095 -1122 5129
rect -1168 5057 -1122 5095
rect -1168 5023 -1162 5057
rect -1128 5023 -1122 5057
rect -1168 4985 -1122 5023
rect -1168 4951 -1162 4985
rect -1128 4951 -1122 4985
rect -1168 4936 -1122 4951
rect -1070 5921 -1024 5936
rect -1070 5887 -1064 5921
rect -1030 5887 -1024 5921
rect -1070 5849 -1024 5887
rect -1070 5815 -1064 5849
rect -1030 5815 -1024 5849
rect -1070 5777 -1024 5815
rect -1070 5743 -1064 5777
rect -1030 5743 -1024 5777
rect -1070 5705 -1024 5743
rect -1070 5671 -1064 5705
rect -1030 5671 -1024 5705
rect -1070 5633 -1024 5671
rect -1070 5599 -1064 5633
rect -1030 5599 -1024 5633
rect -1070 5561 -1024 5599
rect -1070 5527 -1064 5561
rect -1030 5527 -1024 5561
rect -1070 5489 -1024 5527
rect -1070 5455 -1064 5489
rect -1030 5455 -1024 5489
rect -1070 5417 -1024 5455
rect -1070 5383 -1064 5417
rect -1030 5383 -1024 5417
rect -1070 5345 -1024 5383
rect -1070 5311 -1064 5345
rect -1030 5311 -1024 5345
rect -1070 5273 -1024 5311
rect -1070 5239 -1064 5273
rect -1030 5239 -1024 5273
rect -1070 5201 -1024 5239
rect -1070 5167 -1064 5201
rect -1030 5167 -1024 5201
rect -1070 5129 -1024 5167
rect -1070 5095 -1064 5129
rect -1030 5095 -1024 5129
rect -1070 5057 -1024 5095
rect -1070 5023 -1064 5057
rect -1030 5023 -1024 5057
rect -1070 4985 -1024 5023
rect -1070 4951 -1064 4985
rect -1030 4951 -1024 4985
rect -1070 4936 -1024 4951
rect -972 5921 -926 5936
rect -972 5887 -966 5921
rect -932 5887 -926 5921
rect -972 5849 -926 5887
rect -972 5815 -966 5849
rect -932 5815 -926 5849
rect -972 5777 -926 5815
rect -972 5743 -966 5777
rect -932 5743 -926 5777
rect -972 5705 -926 5743
rect -972 5671 -966 5705
rect -932 5671 -926 5705
rect -972 5633 -926 5671
rect -972 5599 -966 5633
rect -932 5599 -926 5633
rect -972 5561 -926 5599
rect -972 5527 -966 5561
rect -932 5527 -926 5561
rect -972 5489 -926 5527
rect -972 5455 -966 5489
rect -932 5455 -926 5489
rect -972 5417 -926 5455
rect -972 5383 -966 5417
rect -932 5383 -926 5417
rect -972 5345 -926 5383
rect -972 5311 -966 5345
rect -932 5311 -926 5345
rect -972 5273 -926 5311
rect -972 5239 -966 5273
rect -932 5239 -926 5273
rect -972 5201 -926 5239
rect -972 5167 -966 5201
rect -932 5167 -926 5201
rect -972 5129 -926 5167
rect -972 5095 -966 5129
rect -932 5095 -926 5129
rect -972 5057 -926 5095
rect -972 5023 -966 5057
rect -932 5023 -926 5057
rect -972 4985 -926 5023
rect -972 4951 -966 4985
rect -932 4951 -926 4985
rect -972 4936 -926 4951
rect -874 5921 -828 5936
rect -874 5887 -868 5921
rect -834 5887 -828 5921
rect -874 5849 -828 5887
rect -874 5815 -868 5849
rect -834 5815 -828 5849
rect -874 5777 -828 5815
rect -874 5743 -868 5777
rect -834 5743 -828 5777
rect -874 5705 -828 5743
rect -874 5671 -868 5705
rect -834 5671 -828 5705
rect -874 5633 -828 5671
rect -874 5599 -868 5633
rect -834 5599 -828 5633
rect -874 5561 -828 5599
rect -874 5527 -868 5561
rect -834 5527 -828 5561
rect -874 5489 -828 5527
rect -874 5455 -868 5489
rect -834 5455 -828 5489
rect -874 5417 -828 5455
rect -874 5383 -868 5417
rect -834 5383 -828 5417
rect -874 5345 -828 5383
rect -874 5311 -868 5345
rect -834 5311 -828 5345
rect -874 5273 -828 5311
rect -874 5239 -868 5273
rect -834 5239 -828 5273
rect -874 5201 -828 5239
rect -874 5167 -868 5201
rect -834 5167 -828 5201
rect -874 5129 -828 5167
rect -874 5095 -868 5129
rect -834 5095 -828 5129
rect -874 5057 -828 5095
rect -874 5023 -868 5057
rect -834 5023 -828 5057
rect -874 4985 -828 5023
rect -874 4951 -868 4985
rect -834 4951 -828 4985
rect -874 4936 -828 4951
rect -21020 4813 -20676 4826
rect -23016 4632 -23006 4812
rect -22698 4632 -22688 4812
rect -21020 4633 -21002 4813
rect -20694 4633 -20676 4813
rect -21020 4620 -20676 4633
rect -19020 4811 -18680 4826
rect -19020 4631 -19004 4811
rect -18696 4631 -18680 4811
rect -16400 4824 -16064 4834
rect -16400 4644 -16386 4824
rect -16078 4644 -16064 4824
rect -16400 4634 -16064 4644
rect -14402 4825 -14054 4838
rect -14402 4645 -14382 4825
rect -14074 4645 -14054 4825
rect -14402 4632 -14054 4645
rect -12402 4827 -12058 4838
rect -12402 4647 -12384 4827
rect -12076 4647 -12058 4827
rect -12402 4636 -12058 4647
rect -10052 4822 -9712 4836
rect -10052 4642 -10036 4822
rect -9728 4642 -9712 4822
rect -19020 4616 -18680 4631
rect -10052 4628 -9712 4642
rect -8052 4820 -7714 4836
rect -8052 4640 -8037 4820
rect -7729 4640 -7714 4820
rect -8052 4624 -7714 4640
rect -6052 4820 -5712 4836
rect -6052 4640 -6036 4820
rect -5728 4640 -5712 4820
rect -6052 4624 -5712 4640
rect -1126 4792 -1022 4794
rect -558 4792 -402 6998
rect 274 6807 336 6998
rect 274 6773 288 6807
rect 322 6773 336 6807
rect 274 6762 336 6773
rect 722 6906 2486 6912
rect 722 6896 2488 6906
rect 722 6892 1694 6896
rect 722 6858 764 6892
rect 798 6858 1694 6892
rect 722 6792 1694 6858
rect 1888 6792 2488 6896
rect 2758 6809 2960 6814
rect 722 6788 2488 6792
rect 722 6754 2440 6788
rect 2474 6754 2488 6788
rect 2716 6803 2893 6809
rect 2716 6769 2728 6803
rect 2762 6769 2893 6803
rect 2716 6763 2893 6769
rect 722 6748 2488 6754
rect 2758 6757 2893 6763
rect 2945 6757 2960 6809
rect 2758 6752 2960 6757
rect 3230 6791 3292 6998
rect 3230 6757 3244 6791
rect 3278 6757 3292 6791
rect 2428 6744 2488 6748
rect 3230 6742 3292 6757
rect 3682 6880 5446 6892
rect 3682 6876 4552 6880
rect 3682 6842 3720 6876
rect 3754 6842 4552 6876
rect 3682 6776 4552 6842
rect 4746 6776 5446 6880
rect 5908 6803 5990 6806
rect 5908 6800 5923 6803
rect 5706 6793 5923 6800
rect 3682 6772 5446 6776
rect 3682 6738 5396 6772
rect 5430 6738 5446 6772
rect 5672 6787 5923 6793
rect 5672 6753 5684 6787
rect 5718 6753 5923 6787
rect 5672 6751 5923 6753
rect 5975 6751 5990 6803
rect 5672 6748 5990 6751
rect 6260 6791 6322 6998
rect 6260 6757 6274 6791
rect 6308 6757 6322 6791
rect 5672 6747 5950 6748
rect 5706 6742 5950 6747
rect 6260 6744 6322 6757
rect 6712 6878 8476 6892
rect 6712 6876 7486 6878
rect 6712 6842 6750 6876
rect 6784 6842 7486 6876
rect 6712 6774 7486 6842
rect 7680 6774 8476 6878
rect 8740 6799 8972 6804
rect 8740 6793 8905 6799
rect 6712 6772 8476 6774
rect 3682 6728 5446 6738
rect 6712 6738 8426 6772
rect 8460 6738 8476 6772
rect 8702 6787 8905 6793
rect 8702 6753 8714 6787
rect 8748 6753 8905 6787
rect 8702 6747 8905 6753
rect 8957 6747 8972 6799
rect 8740 6742 8972 6747
rect 9348 6789 9410 6998
rect 9348 6755 9362 6789
rect 9396 6755 9410 6789
rect 9348 6742 9410 6755
rect 9798 6878 11576 6892
rect 9798 6874 10568 6878
rect 9798 6840 9838 6874
rect 9872 6840 10568 6874
rect 9798 6774 10568 6840
rect 10762 6774 11576 6878
rect 11814 6801 12122 6806
rect 11814 6791 12055 6801
rect 9798 6770 11576 6774
rect 6712 6728 8476 6738
rect 9798 6736 11514 6770
rect 11548 6736 11576 6770
rect 11790 6785 12055 6791
rect 11790 6751 11802 6785
rect 11836 6751 12055 6785
rect 11790 6749 12055 6751
rect 12107 6749 12122 6801
rect 11790 6745 12122 6749
rect 11814 6744 12122 6745
rect 12504 6763 12566 6998
rect 9798 6726 11576 6736
rect 12504 6729 12518 6763
rect 12552 6729 12566 6763
rect 12504 6718 12566 6729
rect 12964 6852 14728 6866
rect 12964 6848 13724 6852
rect 12964 6814 12994 6848
rect 13028 6814 13724 6848
rect 12964 6748 13724 6814
rect 13918 6748 14728 6852
rect 12964 6744 14728 6748
rect 12964 6710 14670 6744
rect 14704 6710 14728 6744
rect 14844 6769 14978 6774
rect 14844 6717 14855 6769
rect 14907 6765 14978 6769
rect 14907 6759 15004 6765
rect 14907 6725 14958 6759
rect 14992 6725 15004 6759
rect 14907 6719 15004 6725
rect 14907 6717 14978 6719
rect 14844 6712 14978 6717
rect 12964 6702 14728 6710
rect 14658 6700 14718 6702
rect 188 6591 234 6606
rect 188 6557 194 6591
rect 228 6557 234 6591
rect 188 6519 234 6557
rect 188 6485 194 6519
rect 228 6485 234 6519
rect 188 6447 234 6485
rect 188 6413 194 6447
rect 228 6413 234 6447
rect 188 6375 234 6413
rect 188 6341 194 6375
rect 228 6341 234 6375
rect 188 6303 234 6341
rect 188 6269 194 6303
rect 228 6269 234 6303
rect 188 6231 234 6269
rect 188 6197 194 6231
rect 228 6197 234 6231
rect 188 6159 234 6197
rect 188 6125 194 6159
rect 228 6125 234 6159
rect 188 6087 234 6125
rect 188 6053 194 6087
rect 228 6053 234 6087
rect 188 6015 234 6053
rect 188 5981 194 6015
rect 228 5981 234 6015
rect 188 5943 234 5981
rect 188 5909 194 5943
rect 228 5909 234 5943
rect 188 5871 234 5909
rect 188 5837 194 5871
rect 228 5837 234 5871
rect 188 5799 234 5837
rect 188 5765 194 5799
rect 228 5765 234 5799
rect 188 5727 234 5765
rect 188 5693 194 5727
rect 228 5693 234 5727
rect 188 5655 234 5693
rect 188 5621 194 5655
rect 228 5621 234 5655
rect 188 5606 234 5621
rect 284 6591 330 6606
rect 284 6557 290 6591
rect 324 6557 330 6591
rect 284 6519 330 6557
rect 284 6485 290 6519
rect 324 6485 330 6519
rect 284 6447 330 6485
rect 284 6413 290 6447
rect 324 6413 330 6447
rect 284 6375 330 6413
rect 284 6341 290 6375
rect 324 6341 330 6375
rect 284 6303 330 6341
rect 284 6269 290 6303
rect 324 6269 330 6303
rect 284 6231 330 6269
rect 284 6197 290 6231
rect 324 6197 330 6231
rect 284 6159 330 6197
rect 284 6125 290 6159
rect 324 6125 330 6159
rect 284 6087 330 6125
rect 284 6053 290 6087
rect 324 6053 330 6087
rect 284 6015 330 6053
rect 284 5981 290 6015
rect 324 5981 330 6015
rect 284 5943 330 5981
rect 284 5909 290 5943
rect 324 5909 330 5943
rect 284 5871 330 5909
rect 284 5837 290 5871
rect 324 5837 330 5871
rect 284 5799 330 5837
rect 284 5765 290 5799
rect 324 5765 330 5799
rect 284 5727 330 5765
rect 284 5693 290 5727
rect 324 5693 330 5727
rect 284 5655 330 5693
rect 284 5621 290 5655
rect 324 5621 330 5655
rect 284 5606 330 5621
rect 380 6591 426 6606
rect 380 6557 386 6591
rect 420 6557 426 6591
rect 380 6519 426 6557
rect 380 6485 386 6519
rect 420 6485 426 6519
rect 380 6447 426 6485
rect 380 6413 386 6447
rect 420 6413 426 6447
rect 380 6375 426 6413
rect 380 6341 386 6375
rect 420 6341 426 6375
rect 380 6303 426 6341
rect 380 6269 386 6303
rect 420 6269 426 6303
rect 380 6231 426 6269
rect 380 6197 386 6231
rect 420 6197 426 6231
rect 380 6159 426 6197
rect 380 6125 386 6159
rect 420 6125 426 6159
rect 380 6087 426 6125
rect 380 6053 386 6087
rect 420 6053 426 6087
rect 380 6015 426 6053
rect 380 5981 386 6015
rect 420 5981 426 6015
rect 380 5943 426 5981
rect 380 5909 386 5943
rect 420 5909 426 5943
rect 380 5871 426 5909
rect 380 5837 386 5871
rect 420 5837 426 5871
rect 380 5799 426 5837
rect 380 5765 386 5799
rect 420 5765 426 5799
rect 380 5727 426 5765
rect 380 5693 386 5727
rect 420 5693 426 5727
rect 380 5655 426 5693
rect 380 5621 386 5655
rect 420 5621 426 5655
rect 380 5606 426 5621
rect 476 6591 522 6606
rect 476 6557 482 6591
rect 516 6557 522 6591
rect 476 6519 522 6557
rect 476 6485 482 6519
rect 516 6485 522 6519
rect 476 6447 522 6485
rect 476 6413 482 6447
rect 516 6413 522 6447
rect 476 6375 522 6413
rect 476 6341 482 6375
rect 516 6341 522 6375
rect 476 6303 522 6341
rect 476 6269 482 6303
rect 516 6269 522 6303
rect 476 6231 522 6269
rect 476 6197 482 6231
rect 516 6197 522 6231
rect 476 6159 522 6197
rect 476 6125 482 6159
rect 516 6125 522 6159
rect 476 6087 522 6125
rect 476 6053 482 6087
rect 516 6053 522 6087
rect 476 6015 522 6053
rect 476 5981 482 6015
rect 516 5981 522 6015
rect 476 5943 522 5981
rect 476 5909 482 5943
rect 516 5909 522 5943
rect 476 5871 522 5909
rect 476 5837 482 5871
rect 516 5837 522 5871
rect 476 5799 522 5837
rect 476 5765 482 5799
rect 516 5765 522 5799
rect 476 5727 522 5765
rect 476 5693 482 5727
rect 516 5693 522 5727
rect 476 5655 522 5693
rect 476 5621 482 5655
rect 516 5621 522 5655
rect 476 5606 522 5621
rect 572 6591 618 6606
rect 572 6557 578 6591
rect 612 6557 618 6591
rect 572 6519 618 6557
rect 572 6485 578 6519
rect 612 6485 618 6519
rect 572 6447 618 6485
rect 572 6413 578 6447
rect 612 6413 618 6447
rect 572 6375 618 6413
rect 572 6341 578 6375
rect 612 6341 618 6375
rect 572 6303 618 6341
rect 572 6269 578 6303
rect 612 6269 618 6303
rect 572 6231 618 6269
rect 572 6197 578 6231
rect 612 6197 618 6231
rect 572 6159 618 6197
rect 572 6125 578 6159
rect 612 6125 618 6159
rect 572 6087 618 6125
rect 572 6053 578 6087
rect 612 6053 618 6087
rect 572 6015 618 6053
rect 572 5981 578 6015
rect 612 5981 618 6015
rect 572 5943 618 5981
rect 572 5909 578 5943
rect 612 5909 618 5943
rect 572 5871 618 5909
rect 572 5837 578 5871
rect 612 5837 618 5871
rect 572 5799 618 5837
rect 572 5765 578 5799
rect 612 5765 618 5799
rect 572 5727 618 5765
rect 572 5693 578 5727
rect 612 5693 618 5727
rect 572 5655 618 5693
rect 572 5621 578 5655
rect 612 5621 618 5655
rect 572 5606 618 5621
rect 668 6591 714 6606
rect 668 6557 674 6591
rect 708 6557 714 6591
rect 668 6519 714 6557
rect 668 6485 674 6519
rect 708 6485 714 6519
rect 668 6447 714 6485
rect 668 6413 674 6447
rect 708 6413 714 6447
rect 668 6375 714 6413
rect 668 6341 674 6375
rect 708 6341 714 6375
rect 668 6303 714 6341
rect 668 6269 674 6303
rect 708 6269 714 6303
rect 668 6231 714 6269
rect 668 6197 674 6231
rect 708 6197 714 6231
rect 668 6159 714 6197
rect 668 6125 674 6159
rect 708 6125 714 6159
rect 668 6087 714 6125
rect 668 6053 674 6087
rect 708 6053 714 6087
rect 668 6015 714 6053
rect 668 5981 674 6015
rect 708 5981 714 6015
rect 668 5943 714 5981
rect 668 5909 674 5943
rect 708 5909 714 5943
rect 668 5871 714 5909
rect 668 5837 674 5871
rect 708 5837 714 5871
rect 668 5799 714 5837
rect 668 5765 674 5799
rect 708 5765 714 5799
rect 668 5727 714 5765
rect 668 5693 674 5727
rect 708 5693 714 5727
rect 668 5655 714 5693
rect 668 5621 674 5655
rect 708 5621 714 5655
rect 668 5606 714 5621
rect 764 6591 810 6606
rect 764 6557 770 6591
rect 804 6557 810 6591
rect 764 6519 810 6557
rect 764 6485 770 6519
rect 804 6485 810 6519
rect 764 6447 810 6485
rect 764 6413 770 6447
rect 804 6413 810 6447
rect 764 6375 810 6413
rect 764 6341 770 6375
rect 804 6341 810 6375
rect 764 6303 810 6341
rect 764 6269 770 6303
rect 804 6269 810 6303
rect 764 6231 810 6269
rect 764 6197 770 6231
rect 804 6197 810 6231
rect 764 6159 810 6197
rect 764 6125 770 6159
rect 804 6125 810 6159
rect 764 6087 810 6125
rect 764 6053 770 6087
rect 804 6053 810 6087
rect 764 6015 810 6053
rect 764 5981 770 6015
rect 804 5981 810 6015
rect 764 5943 810 5981
rect 764 5909 770 5943
rect 804 5909 810 5943
rect 764 5871 810 5909
rect 764 5837 770 5871
rect 804 5837 810 5871
rect 764 5799 810 5837
rect 764 5765 770 5799
rect 804 5765 810 5799
rect 764 5727 810 5765
rect 764 5693 770 5727
rect 804 5693 810 5727
rect 764 5655 810 5693
rect 764 5621 770 5655
rect 804 5621 810 5655
rect 764 5606 810 5621
rect 860 6591 906 6606
rect 860 6557 866 6591
rect 900 6557 906 6591
rect 860 6519 906 6557
rect 860 6485 866 6519
rect 900 6485 906 6519
rect 860 6447 906 6485
rect 860 6413 866 6447
rect 900 6413 906 6447
rect 860 6375 906 6413
rect 860 6341 866 6375
rect 900 6341 906 6375
rect 860 6303 906 6341
rect 860 6269 866 6303
rect 900 6269 906 6303
rect 860 6231 906 6269
rect 860 6197 866 6231
rect 900 6197 906 6231
rect 860 6159 906 6197
rect 860 6125 866 6159
rect 900 6125 906 6159
rect 860 6087 906 6125
rect 860 6053 866 6087
rect 900 6053 906 6087
rect 860 6015 906 6053
rect 860 5981 866 6015
rect 900 5981 906 6015
rect 860 5943 906 5981
rect 860 5909 866 5943
rect 900 5909 906 5943
rect 860 5871 906 5909
rect 860 5837 866 5871
rect 900 5837 906 5871
rect 860 5799 906 5837
rect 860 5765 866 5799
rect 900 5765 906 5799
rect 860 5727 906 5765
rect 860 5693 866 5727
rect 900 5693 906 5727
rect 860 5655 906 5693
rect 860 5621 866 5655
rect 900 5621 906 5655
rect 860 5606 906 5621
rect 956 6591 1002 6606
rect 956 6557 962 6591
rect 996 6557 1002 6591
rect 956 6519 1002 6557
rect 956 6485 962 6519
rect 996 6485 1002 6519
rect 956 6447 1002 6485
rect 956 6413 962 6447
rect 996 6413 1002 6447
rect 956 6375 1002 6413
rect 956 6341 962 6375
rect 996 6341 1002 6375
rect 956 6303 1002 6341
rect 956 6269 962 6303
rect 996 6269 1002 6303
rect 956 6231 1002 6269
rect 956 6197 962 6231
rect 996 6197 1002 6231
rect 956 6159 1002 6197
rect 956 6125 962 6159
rect 996 6125 1002 6159
rect 956 6087 1002 6125
rect 956 6053 962 6087
rect 996 6053 1002 6087
rect 956 6015 1002 6053
rect 956 5981 962 6015
rect 996 5981 1002 6015
rect 956 5943 1002 5981
rect 956 5909 962 5943
rect 996 5909 1002 5943
rect 956 5871 1002 5909
rect 956 5837 962 5871
rect 996 5837 1002 5871
rect 956 5799 1002 5837
rect 956 5765 962 5799
rect 996 5765 1002 5799
rect 956 5727 1002 5765
rect 956 5693 962 5727
rect 996 5693 1002 5727
rect 956 5655 1002 5693
rect 956 5621 962 5655
rect 996 5621 1002 5655
rect 956 5606 1002 5621
rect 1052 6591 1098 6606
rect 1052 6557 1058 6591
rect 1092 6557 1098 6591
rect 1052 6519 1098 6557
rect 1052 6485 1058 6519
rect 1092 6485 1098 6519
rect 1052 6447 1098 6485
rect 1052 6413 1058 6447
rect 1092 6413 1098 6447
rect 1052 6375 1098 6413
rect 1052 6341 1058 6375
rect 1092 6341 1098 6375
rect 1052 6303 1098 6341
rect 1052 6269 1058 6303
rect 1092 6269 1098 6303
rect 1052 6231 1098 6269
rect 1052 6197 1058 6231
rect 1092 6197 1098 6231
rect 1052 6159 1098 6197
rect 1052 6125 1058 6159
rect 1092 6125 1098 6159
rect 1052 6087 1098 6125
rect 1052 6053 1058 6087
rect 1092 6053 1098 6087
rect 1052 6015 1098 6053
rect 1052 5981 1058 6015
rect 1092 5981 1098 6015
rect 1052 5943 1098 5981
rect 1052 5909 1058 5943
rect 1092 5909 1098 5943
rect 1052 5871 1098 5909
rect 1052 5837 1058 5871
rect 1092 5837 1098 5871
rect 1052 5799 1098 5837
rect 1052 5765 1058 5799
rect 1092 5765 1098 5799
rect 1052 5727 1098 5765
rect 1052 5693 1058 5727
rect 1092 5693 1098 5727
rect 1052 5655 1098 5693
rect 1052 5621 1058 5655
rect 1092 5621 1098 5655
rect 1052 5606 1098 5621
rect 1148 6591 1194 6606
rect 1148 6557 1154 6591
rect 1188 6557 1194 6591
rect 1148 6519 1194 6557
rect 1148 6485 1154 6519
rect 1188 6485 1194 6519
rect 1148 6447 1194 6485
rect 1148 6413 1154 6447
rect 1188 6413 1194 6447
rect 1148 6375 1194 6413
rect 1148 6341 1154 6375
rect 1188 6341 1194 6375
rect 1148 6303 1194 6341
rect 1148 6269 1154 6303
rect 1188 6269 1194 6303
rect 1148 6231 1194 6269
rect 1148 6197 1154 6231
rect 1188 6197 1194 6231
rect 1148 6159 1194 6197
rect 1148 6125 1154 6159
rect 1188 6125 1194 6159
rect 1148 6087 1194 6125
rect 1148 6053 1154 6087
rect 1188 6053 1194 6087
rect 1148 6015 1194 6053
rect 1148 5981 1154 6015
rect 1188 5981 1194 6015
rect 1148 5943 1194 5981
rect 1148 5909 1154 5943
rect 1188 5909 1194 5943
rect 1148 5871 1194 5909
rect 1148 5837 1154 5871
rect 1188 5837 1194 5871
rect 1148 5799 1194 5837
rect 1148 5765 1154 5799
rect 1188 5765 1194 5799
rect 1148 5727 1194 5765
rect 1148 5693 1154 5727
rect 1188 5693 1194 5727
rect 1148 5655 1194 5693
rect 1148 5621 1154 5655
rect 1188 5621 1194 5655
rect 1148 5606 1194 5621
rect 1244 6591 1290 6606
rect 1244 6557 1250 6591
rect 1284 6557 1290 6591
rect 1244 6519 1290 6557
rect 1244 6485 1250 6519
rect 1284 6485 1290 6519
rect 1244 6447 1290 6485
rect 1244 6413 1250 6447
rect 1284 6413 1290 6447
rect 1244 6375 1290 6413
rect 1244 6341 1250 6375
rect 1284 6341 1290 6375
rect 1244 6303 1290 6341
rect 1244 6269 1250 6303
rect 1284 6269 1290 6303
rect 1244 6231 1290 6269
rect 1244 6197 1250 6231
rect 1284 6197 1290 6231
rect 1244 6159 1290 6197
rect 1244 6125 1250 6159
rect 1284 6125 1290 6159
rect 1244 6087 1290 6125
rect 1244 6053 1250 6087
rect 1284 6053 1290 6087
rect 1244 6015 1290 6053
rect 1244 5981 1250 6015
rect 1284 5981 1290 6015
rect 1244 5943 1290 5981
rect 1244 5909 1250 5943
rect 1284 5909 1290 5943
rect 1244 5871 1290 5909
rect 1244 5837 1250 5871
rect 1284 5837 1290 5871
rect 1244 5799 1290 5837
rect 1244 5765 1250 5799
rect 1284 5765 1290 5799
rect 1244 5727 1290 5765
rect 1244 5693 1250 5727
rect 1284 5693 1290 5727
rect 1244 5655 1290 5693
rect 1244 5621 1250 5655
rect 1284 5621 1290 5655
rect 1244 5606 1290 5621
rect 1340 6591 1386 6606
rect 1340 6557 1346 6591
rect 1380 6557 1386 6591
rect 1340 6519 1386 6557
rect 1340 6485 1346 6519
rect 1380 6485 1386 6519
rect 1340 6447 1386 6485
rect 1340 6413 1346 6447
rect 1380 6413 1386 6447
rect 1340 6375 1386 6413
rect 1340 6341 1346 6375
rect 1380 6341 1386 6375
rect 1340 6303 1386 6341
rect 1340 6269 1346 6303
rect 1380 6269 1386 6303
rect 1340 6231 1386 6269
rect 1340 6197 1346 6231
rect 1380 6197 1386 6231
rect 1340 6159 1386 6197
rect 1340 6125 1346 6159
rect 1380 6125 1386 6159
rect 1340 6087 1386 6125
rect 1340 6053 1346 6087
rect 1380 6053 1386 6087
rect 1340 6015 1386 6053
rect 1340 5981 1346 6015
rect 1380 5981 1386 6015
rect 1340 5943 1386 5981
rect 1340 5909 1346 5943
rect 1380 5909 1386 5943
rect 1340 5871 1386 5909
rect 1340 5837 1346 5871
rect 1380 5837 1386 5871
rect 1340 5799 1386 5837
rect 1340 5765 1346 5799
rect 1380 5765 1386 5799
rect 1340 5727 1386 5765
rect 1340 5693 1346 5727
rect 1380 5693 1386 5727
rect 1340 5655 1386 5693
rect 1340 5621 1346 5655
rect 1380 5621 1386 5655
rect 1340 5606 1386 5621
rect 1954 6587 2000 6602
rect 1954 6553 1960 6587
rect 1994 6553 2000 6587
rect 1954 6515 2000 6553
rect 1954 6481 1960 6515
rect 1994 6481 2000 6515
rect 1954 6443 2000 6481
rect 1954 6409 1960 6443
rect 1994 6409 2000 6443
rect 1954 6371 2000 6409
rect 1954 6337 1960 6371
rect 1994 6337 2000 6371
rect 1954 6299 2000 6337
rect 1954 6265 1960 6299
rect 1994 6265 2000 6299
rect 1954 6227 2000 6265
rect 1954 6193 1960 6227
rect 1994 6193 2000 6227
rect 1954 6155 2000 6193
rect 1954 6121 1960 6155
rect 1994 6121 2000 6155
rect 1954 6083 2000 6121
rect 1954 6049 1960 6083
rect 1994 6049 2000 6083
rect 1954 6011 2000 6049
rect 1954 5977 1960 6011
rect 1994 5977 2000 6011
rect 1954 5939 2000 5977
rect 1954 5905 1960 5939
rect 1994 5905 2000 5939
rect 1954 5867 2000 5905
rect 1954 5833 1960 5867
rect 1994 5833 2000 5867
rect 1954 5795 2000 5833
rect 1954 5761 1960 5795
rect 1994 5761 2000 5795
rect 1954 5723 2000 5761
rect 1954 5689 1960 5723
rect 1994 5689 2000 5723
rect 1954 5651 2000 5689
rect 1954 5617 1960 5651
rect 1994 5617 2000 5651
rect 1954 5602 2000 5617
rect 2050 6587 2096 6602
rect 2050 6553 2056 6587
rect 2090 6553 2096 6587
rect 2050 6515 2096 6553
rect 2050 6481 2056 6515
rect 2090 6481 2096 6515
rect 2050 6443 2096 6481
rect 2050 6409 2056 6443
rect 2090 6409 2096 6443
rect 2050 6371 2096 6409
rect 2050 6337 2056 6371
rect 2090 6337 2096 6371
rect 2050 6299 2096 6337
rect 2050 6265 2056 6299
rect 2090 6265 2096 6299
rect 2050 6227 2096 6265
rect 2050 6193 2056 6227
rect 2090 6193 2096 6227
rect 2050 6155 2096 6193
rect 2050 6121 2056 6155
rect 2090 6121 2096 6155
rect 2050 6083 2096 6121
rect 2050 6049 2056 6083
rect 2090 6049 2096 6083
rect 2050 6011 2096 6049
rect 2050 5977 2056 6011
rect 2090 5977 2096 6011
rect 2050 5939 2096 5977
rect 2050 5905 2056 5939
rect 2090 5905 2096 5939
rect 2050 5867 2096 5905
rect 2050 5833 2056 5867
rect 2090 5833 2096 5867
rect 2050 5795 2096 5833
rect 2050 5761 2056 5795
rect 2090 5761 2096 5795
rect 2050 5723 2096 5761
rect 2050 5689 2056 5723
rect 2090 5689 2096 5723
rect 2050 5651 2096 5689
rect 2050 5617 2056 5651
rect 2090 5617 2096 5651
rect 2050 5602 2096 5617
rect 2146 6587 2192 6602
rect 2146 6553 2152 6587
rect 2186 6553 2192 6587
rect 2146 6515 2192 6553
rect 2146 6481 2152 6515
rect 2186 6481 2192 6515
rect 2146 6443 2192 6481
rect 2146 6409 2152 6443
rect 2186 6409 2192 6443
rect 2146 6371 2192 6409
rect 2146 6337 2152 6371
rect 2186 6337 2192 6371
rect 2146 6299 2192 6337
rect 2146 6265 2152 6299
rect 2186 6265 2192 6299
rect 2146 6227 2192 6265
rect 2146 6193 2152 6227
rect 2186 6193 2192 6227
rect 2146 6155 2192 6193
rect 2146 6121 2152 6155
rect 2186 6121 2192 6155
rect 2146 6083 2192 6121
rect 2146 6049 2152 6083
rect 2186 6049 2192 6083
rect 2146 6011 2192 6049
rect 2146 5977 2152 6011
rect 2186 5977 2192 6011
rect 2146 5939 2192 5977
rect 2146 5905 2152 5939
rect 2186 5905 2192 5939
rect 2146 5867 2192 5905
rect 2146 5833 2152 5867
rect 2186 5833 2192 5867
rect 2146 5795 2192 5833
rect 2146 5761 2152 5795
rect 2186 5761 2192 5795
rect 2146 5723 2192 5761
rect 2146 5689 2152 5723
rect 2186 5689 2192 5723
rect 2146 5651 2192 5689
rect 2146 5617 2152 5651
rect 2186 5617 2192 5651
rect 2146 5602 2192 5617
rect 2242 6587 2288 6602
rect 2242 6553 2248 6587
rect 2282 6553 2288 6587
rect 2242 6515 2288 6553
rect 2242 6481 2248 6515
rect 2282 6481 2288 6515
rect 2242 6443 2288 6481
rect 2242 6409 2248 6443
rect 2282 6409 2288 6443
rect 2242 6371 2288 6409
rect 2242 6337 2248 6371
rect 2282 6337 2288 6371
rect 2242 6299 2288 6337
rect 2242 6265 2248 6299
rect 2282 6265 2288 6299
rect 2242 6227 2288 6265
rect 2242 6193 2248 6227
rect 2282 6193 2288 6227
rect 2242 6155 2288 6193
rect 2242 6121 2248 6155
rect 2282 6121 2288 6155
rect 2242 6083 2288 6121
rect 2242 6049 2248 6083
rect 2282 6049 2288 6083
rect 2242 6011 2288 6049
rect 2242 5977 2248 6011
rect 2282 5977 2288 6011
rect 2242 5939 2288 5977
rect 2242 5905 2248 5939
rect 2282 5905 2288 5939
rect 2242 5867 2288 5905
rect 2242 5833 2248 5867
rect 2282 5833 2288 5867
rect 2242 5795 2288 5833
rect 2242 5761 2248 5795
rect 2282 5761 2288 5795
rect 2242 5723 2288 5761
rect 2242 5689 2248 5723
rect 2282 5689 2288 5723
rect 2242 5651 2288 5689
rect 2242 5617 2248 5651
rect 2282 5617 2288 5651
rect 2242 5602 2288 5617
rect 2338 6587 2384 6602
rect 2338 6553 2344 6587
rect 2378 6553 2384 6587
rect 2338 6515 2384 6553
rect 2338 6481 2344 6515
rect 2378 6481 2384 6515
rect 2338 6443 2384 6481
rect 2338 6409 2344 6443
rect 2378 6409 2384 6443
rect 2338 6371 2384 6409
rect 2338 6337 2344 6371
rect 2378 6337 2384 6371
rect 2338 6299 2384 6337
rect 2338 6265 2344 6299
rect 2378 6265 2384 6299
rect 2338 6227 2384 6265
rect 2338 6193 2344 6227
rect 2378 6193 2384 6227
rect 2338 6155 2384 6193
rect 2338 6121 2344 6155
rect 2378 6121 2384 6155
rect 2338 6083 2384 6121
rect 2338 6049 2344 6083
rect 2378 6049 2384 6083
rect 2338 6011 2384 6049
rect 2338 5977 2344 6011
rect 2378 5977 2384 6011
rect 2338 5939 2384 5977
rect 2338 5905 2344 5939
rect 2378 5905 2384 5939
rect 2338 5867 2384 5905
rect 2338 5833 2344 5867
rect 2378 5833 2384 5867
rect 2338 5795 2384 5833
rect 2338 5761 2344 5795
rect 2378 5761 2384 5795
rect 2338 5723 2384 5761
rect 2338 5689 2344 5723
rect 2378 5689 2384 5723
rect 2338 5651 2384 5689
rect 2338 5617 2344 5651
rect 2378 5617 2384 5651
rect 2338 5602 2384 5617
rect 2434 6587 2480 6602
rect 2434 6553 2440 6587
rect 2474 6553 2480 6587
rect 2434 6515 2480 6553
rect 2434 6481 2440 6515
rect 2474 6481 2480 6515
rect 2434 6443 2480 6481
rect 2434 6409 2440 6443
rect 2474 6409 2480 6443
rect 2434 6371 2480 6409
rect 2434 6337 2440 6371
rect 2474 6337 2480 6371
rect 2434 6299 2480 6337
rect 2434 6265 2440 6299
rect 2474 6265 2480 6299
rect 2434 6227 2480 6265
rect 2434 6193 2440 6227
rect 2474 6193 2480 6227
rect 2434 6155 2480 6193
rect 2434 6121 2440 6155
rect 2474 6121 2480 6155
rect 2434 6083 2480 6121
rect 2434 6049 2440 6083
rect 2474 6049 2480 6083
rect 2434 6011 2480 6049
rect 2434 5977 2440 6011
rect 2474 5977 2480 6011
rect 2434 5939 2480 5977
rect 2434 5905 2440 5939
rect 2474 5905 2480 5939
rect 2434 5867 2480 5905
rect 2434 5833 2440 5867
rect 2474 5833 2480 5867
rect 2434 5795 2480 5833
rect 2434 5761 2440 5795
rect 2474 5761 2480 5795
rect 2434 5723 2480 5761
rect 2434 5689 2440 5723
rect 2474 5689 2480 5723
rect 2434 5651 2480 5689
rect 2434 5617 2440 5651
rect 2474 5617 2480 5651
rect 2434 5602 2480 5617
rect 2530 6587 2576 6602
rect 2530 6553 2536 6587
rect 2570 6553 2576 6587
rect 2530 6515 2576 6553
rect 2530 6481 2536 6515
rect 2570 6481 2576 6515
rect 2530 6443 2576 6481
rect 2530 6409 2536 6443
rect 2570 6409 2576 6443
rect 2530 6371 2576 6409
rect 2530 6337 2536 6371
rect 2570 6337 2576 6371
rect 2530 6299 2576 6337
rect 2530 6265 2536 6299
rect 2570 6265 2576 6299
rect 2530 6227 2576 6265
rect 2530 6193 2536 6227
rect 2570 6193 2576 6227
rect 2530 6155 2576 6193
rect 2530 6121 2536 6155
rect 2570 6121 2576 6155
rect 2530 6083 2576 6121
rect 2530 6049 2536 6083
rect 2570 6049 2576 6083
rect 2530 6011 2576 6049
rect 2530 5977 2536 6011
rect 2570 5977 2576 6011
rect 2530 5939 2576 5977
rect 2530 5905 2536 5939
rect 2570 5905 2576 5939
rect 2530 5867 2576 5905
rect 2530 5833 2536 5867
rect 2570 5833 2576 5867
rect 2530 5795 2576 5833
rect 2530 5761 2536 5795
rect 2570 5761 2576 5795
rect 2530 5723 2576 5761
rect 2530 5689 2536 5723
rect 2570 5689 2576 5723
rect 2530 5651 2576 5689
rect 2530 5617 2536 5651
rect 2570 5617 2576 5651
rect 2530 5602 2576 5617
rect 2626 6587 2672 6602
rect 2626 6553 2632 6587
rect 2666 6553 2672 6587
rect 2626 6515 2672 6553
rect 2626 6481 2632 6515
rect 2666 6481 2672 6515
rect 2626 6443 2672 6481
rect 2626 6409 2632 6443
rect 2666 6409 2672 6443
rect 2626 6371 2672 6409
rect 2626 6337 2632 6371
rect 2666 6337 2672 6371
rect 2626 6299 2672 6337
rect 2626 6265 2632 6299
rect 2666 6265 2672 6299
rect 2626 6227 2672 6265
rect 2626 6193 2632 6227
rect 2666 6193 2672 6227
rect 2626 6155 2672 6193
rect 2626 6121 2632 6155
rect 2666 6121 2672 6155
rect 2626 6083 2672 6121
rect 2626 6049 2632 6083
rect 2666 6049 2672 6083
rect 2626 6011 2672 6049
rect 2626 5977 2632 6011
rect 2666 5977 2672 6011
rect 2626 5939 2672 5977
rect 2626 5905 2632 5939
rect 2666 5905 2672 5939
rect 2626 5867 2672 5905
rect 2626 5833 2632 5867
rect 2666 5833 2672 5867
rect 2626 5795 2672 5833
rect 2626 5761 2632 5795
rect 2666 5761 2672 5795
rect 2626 5723 2672 5761
rect 2626 5689 2632 5723
rect 2666 5689 2672 5723
rect 2626 5651 2672 5689
rect 2626 5617 2632 5651
rect 2666 5617 2672 5651
rect 2626 5602 2672 5617
rect 2722 6587 2768 6602
rect 2722 6553 2728 6587
rect 2762 6553 2768 6587
rect 2722 6515 2768 6553
rect 2722 6481 2728 6515
rect 2762 6481 2768 6515
rect 2722 6443 2768 6481
rect 2722 6409 2728 6443
rect 2762 6409 2768 6443
rect 2722 6371 2768 6409
rect 2722 6337 2728 6371
rect 2762 6337 2768 6371
rect 2722 6299 2768 6337
rect 2722 6265 2728 6299
rect 2762 6265 2768 6299
rect 2722 6227 2768 6265
rect 2722 6193 2728 6227
rect 2762 6193 2768 6227
rect 2722 6155 2768 6193
rect 2722 6121 2728 6155
rect 2762 6121 2768 6155
rect 2722 6083 2768 6121
rect 2722 6049 2728 6083
rect 2762 6049 2768 6083
rect 2722 6011 2768 6049
rect 2722 5977 2728 6011
rect 2762 5977 2768 6011
rect 2722 5939 2768 5977
rect 2722 5905 2728 5939
rect 2762 5905 2768 5939
rect 2722 5867 2768 5905
rect 2722 5833 2728 5867
rect 2762 5833 2768 5867
rect 2722 5795 2768 5833
rect 2722 5761 2728 5795
rect 2762 5761 2768 5795
rect 2722 5723 2768 5761
rect 2722 5689 2728 5723
rect 2762 5689 2768 5723
rect 2722 5651 2768 5689
rect 2722 5617 2728 5651
rect 2762 5617 2768 5651
rect 2722 5602 2768 5617
rect 3144 6575 3190 6590
rect 3144 6541 3150 6575
rect 3184 6541 3190 6575
rect 3144 6503 3190 6541
rect 3144 6469 3150 6503
rect 3184 6469 3190 6503
rect 3144 6431 3190 6469
rect 3144 6397 3150 6431
rect 3184 6397 3190 6431
rect 3144 6359 3190 6397
rect 3144 6325 3150 6359
rect 3184 6325 3190 6359
rect 3144 6287 3190 6325
rect 3144 6253 3150 6287
rect 3184 6253 3190 6287
rect 3144 6215 3190 6253
rect 3144 6181 3150 6215
rect 3184 6181 3190 6215
rect 3144 6143 3190 6181
rect 3144 6109 3150 6143
rect 3184 6109 3190 6143
rect 3144 6071 3190 6109
rect 3144 6037 3150 6071
rect 3184 6037 3190 6071
rect 3144 5999 3190 6037
rect 3144 5965 3150 5999
rect 3184 5965 3190 5999
rect 3144 5927 3190 5965
rect 3144 5893 3150 5927
rect 3184 5893 3190 5927
rect 3144 5855 3190 5893
rect 3144 5821 3150 5855
rect 3184 5821 3190 5855
rect 3144 5783 3190 5821
rect 3144 5749 3150 5783
rect 3184 5749 3190 5783
rect 3144 5711 3190 5749
rect 3144 5677 3150 5711
rect 3184 5677 3190 5711
rect 3144 5639 3190 5677
rect 3144 5605 3150 5639
rect 3184 5605 3190 5639
rect 3144 5590 3190 5605
rect 3240 6575 3286 6590
rect 3240 6541 3246 6575
rect 3280 6541 3286 6575
rect 3240 6503 3286 6541
rect 3240 6469 3246 6503
rect 3280 6469 3286 6503
rect 3240 6431 3286 6469
rect 3240 6397 3246 6431
rect 3280 6397 3286 6431
rect 3240 6359 3286 6397
rect 3240 6325 3246 6359
rect 3280 6325 3286 6359
rect 3240 6287 3286 6325
rect 3240 6253 3246 6287
rect 3280 6253 3286 6287
rect 3240 6215 3286 6253
rect 3240 6181 3246 6215
rect 3280 6181 3286 6215
rect 3240 6143 3286 6181
rect 3240 6109 3246 6143
rect 3280 6109 3286 6143
rect 3240 6071 3286 6109
rect 3240 6037 3246 6071
rect 3280 6037 3286 6071
rect 3240 5999 3286 6037
rect 3240 5965 3246 5999
rect 3280 5965 3286 5999
rect 3240 5927 3286 5965
rect 3240 5893 3246 5927
rect 3280 5893 3286 5927
rect 3240 5855 3286 5893
rect 3240 5821 3246 5855
rect 3280 5821 3286 5855
rect 3240 5783 3286 5821
rect 3240 5749 3246 5783
rect 3280 5749 3286 5783
rect 3240 5711 3286 5749
rect 3240 5677 3246 5711
rect 3280 5677 3286 5711
rect 3240 5639 3286 5677
rect 3240 5605 3246 5639
rect 3280 5605 3286 5639
rect 3240 5590 3286 5605
rect 3336 6575 3382 6590
rect 3336 6541 3342 6575
rect 3376 6541 3382 6575
rect 3336 6503 3382 6541
rect 3336 6469 3342 6503
rect 3376 6469 3382 6503
rect 3336 6431 3382 6469
rect 3336 6397 3342 6431
rect 3376 6397 3382 6431
rect 3336 6359 3382 6397
rect 3336 6325 3342 6359
rect 3376 6325 3382 6359
rect 3336 6287 3382 6325
rect 3336 6253 3342 6287
rect 3376 6253 3382 6287
rect 3336 6215 3382 6253
rect 3336 6181 3342 6215
rect 3376 6181 3382 6215
rect 3336 6143 3382 6181
rect 3336 6109 3342 6143
rect 3376 6109 3382 6143
rect 3336 6071 3382 6109
rect 3336 6037 3342 6071
rect 3376 6037 3382 6071
rect 3336 5999 3382 6037
rect 3336 5965 3342 5999
rect 3376 5965 3382 5999
rect 3336 5927 3382 5965
rect 3336 5893 3342 5927
rect 3376 5893 3382 5927
rect 3336 5855 3382 5893
rect 3336 5821 3342 5855
rect 3376 5821 3382 5855
rect 3336 5783 3382 5821
rect 3336 5749 3342 5783
rect 3376 5749 3382 5783
rect 3336 5711 3382 5749
rect 3336 5677 3342 5711
rect 3376 5677 3382 5711
rect 3336 5639 3382 5677
rect 3336 5605 3342 5639
rect 3376 5605 3382 5639
rect 3336 5590 3382 5605
rect 3432 6575 3478 6590
rect 3432 6541 3438 6575
rect 3472 6541 3478 6575
rect 3432 6503 3478 6541
rect 3432 6469 3438 6503
rect 3472 6469 3478 6503
rect 3432 6431 3478 6469
rect 3432 6397 3438 6431
rect 3472 6397 3478 6431
rect 3432 6359 3478 6397
rect 3432 6325 3438 6359
rect 3472 6325 3478 6359
rect 3432 6287 3478 6325
rect 3432 6253 3438 6287
rect 3472 6253 3478 6287
rect 3432 6215 3478 6253
rect 3432 6181 3438 6215
rect 3472 6181 3478 6215
rect 3432 6143 3478 6181
rect 3432 6109 3438 6143
rect 3472 6109 3478 6143
rect 3432 6071 3478 6109
rect 3432 6037 3438 6071
rect 3472 6037 3478 6071
rect 3432 5999 3478 6037
rect 3432 5965 3438 5999
rect 3472 5965 3478 5999
rect 3432 5927 3478 5965
rect 3432 5893 3438 5927
rect 3472 5893 3478 5927
rect 3432 5855 3478 5893
rect 3432 5821 3438 5855
rect 3472 5821 3478 5855
rect 3432 5783 3478 5821
rect 3432 5749 3438 5783
rect 3472 5749 3478 5783
rect 3432 5711 3478 5749
rect 3432 5677 3438 5711
rect 3472 5677 3478 5711
rect 3432 5639 3478 5677
rect 3432 5605 3438 5639
rect 3472 5605 3478 5639
rect 3432 5590 3478 5605
rect 3528 6575 3574 6590
rect 3528 6541 3534 6575
rect 3568 6541 3574 6575
rect 3528 6503 3574 6541
rect 3528 6469 3534 6503
rect 3568 6469 3574 6503
rect 3528 6431 3574 6469
rect 3528 6397 3534 6431
rect 3568 6397 3574 6431
rect 3528 6359 3574 6397
rect 3528 6325 3534 6359
rect 3568 6325 3574 6359
rect 3528 6287 3574 6325
rect 3528 6253 3534 6287
rect 3568 6253 3574 6287
rect 3528 6215 3574 6253
rect 3528 6181 3534 6215
rect 3568 6181 3574 6215
rect 3528 6143 3574 6181
rect 3528 6109 3534 6143
rect 3568 6109 3574 6143
rect 3528 6071 3574 6109
rect 3528 6037 3534 6071
rect 3568 6037 3574 6071
rect 3528 5999 3574 6037
rect 3528 5965 3534 5999
rect 3568 5965 3574 5999
rect 3528 5927 3574 5965
rect 3528 5893 3534 5927
rect 3568 5893 3574 5927
rect 3528 5855 3574 5893
rect 3528 5821 3534 5855
rect 3568 5821 3574 5855
rect 3528 5783 3574 5821
rect 3528 5749 3534 5783
rect 3568 5749 3574 5783
rect 3528 5711 3574 5749
rect 3528 5677 3534 5711
rect 3568 5677 3574 5711
rect 3528 5639 3574 5677
rect 3528 5605 3534 5639
rect 3568 5605 3574 5639
rect 3528 5590 3574 5605
rect 3624 6575 3670 6590
rect 3624 6541 3630 6575
rect 3664 6541 3670 6575
rect 3624 6503 3670 6541
rect 3624 6469 3630 6503
rect 3664 6469 3670 6503
rect 3624 6431 3670 6469
rect 3624 6397 3630 6431
rect 3664 6397 3670 6431
rect 3624 6359 3670 6397
rect 3624 6325 3630 6359
rect 3664 6325 3670 6359
rect 3624 6287 3670 6325
rect 3624 6253 3630 6287
rect 3664 6253 3670 6287
rect 3624 6215 3670 6253
rect 3624 6181 3630 6215
rect 3664 6181 3670 6215
rect 3624 6143 3670 6181
rect 3624 6109 3630 6143
rect 3664 6109 3670 6143
rect 3624 6071 3670 6109
rect 3624 6037 3630 6071
rect 3664 6037 3670 6071
rect 3624 5999 3670 6037
rect 3624 5965 3630 5999
rect 3664 5965 3670 5999
rect 3624 5927 3670 5965
rect 3624 5893 3630 5927
rect 3664 5893 3670 5927
rect 3624 5855 3670 5893
rect 3624 5821 3630 5855
rect 3664 5821 3670 5855
rect 3624 5783 3670 5821
rect 3624 5749 3630 5783
rect 3664 5749 3670 5783
rect 3624 5711 3670 5749
rect 3624 5677 3630 5711
rect 3664 5677 3670 5711
rect 3624 5639 3670 5677
rect 3624 5605 3630 5639
rect 3664 5605 3670 5639
rect 3624 5590 3670 5605
rect 3720 6575 3766 6590
rect 3720 6541 3726 6575
rect 3760 6541 3766 6575
rect 3720 6503 3766 6541
rect 3720 6469 3726 6503
rect 3760 6469 3766 6503
rect 3720 6431 3766 6469
rect 3720 6397 3726 6431
rect 3760 6397 3766 6431
rect 3720 6359 3766 6397
rect 3720 6325 3726 6359
rect 3760 6325 3766 6359
rect 3720 6287 3766 6325
rect 3720 6253 3726 6287
rect 3760 6253 3766 6287
rect 3720 6215 3766 6253
rect 3720 6181 3726 6215
rect 3760 6181 3766 6215
rect 3720 6143 3766 6181
rect 3720 6109 3726 6143
rect 3760 6109 3766 6143
rect 3720 6071 3766 6109
rect 3720 6037 3726 6071
rect 3760 6037 3766 6071
rect 3720 5999 3766 6037
rect 3720 5965 3726 5999
rect 3760 5965 3766 5999
rect 3720 5927 3766 5965
rect 3720 5893 3726 5927
rect 3760 5893 3766 5927
rect 3720 5855 3766 5893
rect 3720 5821 3726 5855
rect 3760 5821 3766 5855
rect 3720 5783 3766 5821
rect 3720 5749 3726 5783
rect 3760 5749 3766 5783
rect 3720 5711 3766 5749
rect 3720 5677 3726 5711
rect 3760 5677 3766 5711
rect 3720 5639 3766 5677
rect 3720 5605 3726 5639
rect 3760 5605 3766 5639
rect 3720 5590 3766 5605
rect 3816 6575 3862 6590
rect 3816 6541 3822 6575
rect 3856 6541 3862 6575
rect 3816 6503 3862 6541
rect 3816 6469 3822 6503
rect 3856 6469 3862 6503
rect 3816 6431 3862 6469
rect 3816 6397 3822 6431
rect 3856 6397 3862 6431
rect 3816 6359 3862 6397
rect 3816 6325 3822 6359
rect 3856 6325 3862 6359
rect 3816 6287 3862 6325
rect 3816 6253 3822 6287
rect 3856 6253 3862 6287
rect 3816 6215 3862 6253
rect 3816 6181 3822 6215
rect 3856 6181 3862 6215
rect 3816 6143 3862 6181
rect 3816 6109 3822 6143
rect 3856 6109 3862 6143
rect 3816 6071 3862 6109
rect 3816 6037 3822 6071
rect 3856 6037 3862 6071
rect 3816 5999 3862 6037
rect 3816 5965 3822 5999
rect 3856 5965 3862 5999
rect 3816 5927 3862 5965
rect 3816 5893 3822 5927
rect 3856 5893 3862 5927
rect 3816 5855 3862 5893
rect 3816 5821 3822 5855
rect 3856 5821 3862 5855
rect 3816 5783 3862 5821
rect 3816 5749 3822 5783
rect 3856 5749 3862 5783
rect 3816 5711 3862 5749
rect 3816 5677 3822 5711
rect 3856 5677 3862 5711
rect 3816 5639 3862 5677
rect 3816 5605 3822 5639
rect 3856 5605 3862 5639
rect 3816 5590 3862 5605
rect 3912 6575 3958 6590
rect 3912 6541 3918 6575
rect 3952 6541 3958 6575
rect 3912 6503 3958 6541
rect 3912 6469 3918 6503
rect 3952 6469 3958 6503
rect 3912 6431 3958 6469
rect 3912 6397 3918 6431
rect 3952 6397 3958 6431
rect 3912 6359 3958 6397
rect 3912 6325 3918 6359
rect 3952 6325 3958 6359
rect 3912 6287 3958 6325
rect 3912 6253 3918 6287
rect 3952 6253 3958 6287
rect 3912 6215 3958 6253
rect 3912 6181 3918 6215
rect 3952 6181 3958 6215
rect 3912 6143 3958 6181
rect 3912 6109 3918 6143
rect 3952 6109 3958 6143
rect 3912 6071 3958 6109
rect 3912 6037 3918 6071
rect 3952 6037 3958 6071
rect 3912 5999 3958 6037
rect 3912 5965 3918 5999
rect 3952 5965 3958 5999
rect 3912 5927 3958 5965
rect 3912 5893 3918 5927
rect 3952 5893 3958 5927
rect 3912 5855 3958 5893
rect 3912 5821 3918 5855
rect 3952 5821 3958 5855
rect 3912 5783 3958 5821
rect 3912 5749 3918 5783
rect 3952 5749 3958 5783
rect 3912 5711 3958 5749
rect 3912 5677 3918 5711
rect 3952 5677 3958 5711
rect 3912 5639 3958 5677
rect 3912 5605 3918 5639
rect 3952 5605 3958 5639
rect 3912 5590 3958 5605
rect 4008 6575 4054 6590
rect 4008 6541 4014 6575
rect 4048 6541 4054 6575
rect 4008 6503 4054 6541
rect 4008 6469 4014 6503
rect 4048 6469 4054 6503
rect 4008 6431 4054 6469
rect 4008 6397 4014 6431
rect 4048 6397 4054 6431
rect 4008 6359 4054 6397
rect 4008 6325 4014 6359
rect 4048 6325 4054 6359
rect 4008 6287 4054 6325
rect 4008 6253 4014 6287
rect 4048 6253 4054 6287
rect 4008 6215 4054 6253
rect 4008 6181 4014 6215
rect 4048 6181 4054 6215
rect 4008 6143 4054 6181
rect 4008 6109 4014 6143
rect 4048 6109 4054 6143
rect 4008 6071 4054 6109
rect 4008 6037 4014 6071
rect 4048 6037 4054 6071
rect 4008 5999 4054 6037
rect 4008 5965 4014 5999
rect 4048 5965 4054 5999
rect 4008 5927 4054 5965
rect 4008 5893 4014 5927
rect 4048 5893 4054 5927
rect 4008 5855 4054 5893
rect 4008 5821 4014 5855
rect 4048 5821 4054 5855
rect 4008 5783 4054 5821
rect 4008 5749 4014 5783
rect 4048 5749 4054 5783
rect 4008 5711 4054 5749
rect 4008 5677 4014 5711
rect 4048 5677 4054 5711
rect 4008 5639 4054 5677
rect 4008 5605 4014 5639
rect 4048 5605 4054 5639
rect 4008 5590 4054 5605
rect 4104 6575 4150 6590
rect 4104 6541 4110 6575
rect 4144 6541 4150 6575
rect 4104 6503 4150 6541
rect 4104 6469 4110 6503
rect 4144 6469 4150 6503
rect 4104 6431 4150 6469
rect 4104 6397 4110 6431
rect 4144 6397 4150 6431
rect 4104 6359 4150 6397
rect 4104 6325 4110 6359
rect 4144 6325 4150 6359
rect 4104 6287 4150 6325
rect 4104 6253 4110 6287
rect 4144 6253 4150 6287
rect 4104 6215 4150 6253
rect 4104 6181 4110 6215
rect 4144 6181 4150 6215
rect 4104 6143 4150 6181
rect 4104 6109 4110 6143
rect 4144 6109 4150 6143
rect 4104 6071 4150 6109
rect 4104 6037 4110 6071
rect 4144 6037 4150 6071
rect 4104 5999 4150 6037
rect 4104 5965 4110 5999
rect 4144 5965 4150 5999
rect 4104 5927 4150 5965
rect 4104 5893 4110 5927
rect 4144 5893 4150 5927
rect 4104 5855 4150 5893
rect 4104 5821 4110 5855
rect 4144 5821 4150 5855
rect 4104 5783 4150 5821
rect 4104 5749 4110 5783
rect 4144 5749 4150 5783
rect 4104 5711 4150 5749
rect 4104 5677 4110 5711
rect 4144 5677 4150 5711
rect 4104 5639 4150 5677
rect 4104 5605 4110 5639
rect 4144 5605 4150 5639
rect 4104 5590 4150 5605
rect 4200 6575 4246 6590
rect 4200 6541 4206 6575
rect 4240 6541 4246 6575
rect 4200 6503 4246 6541
rect 4200 6469 4206 6503
rect 4240 6469 4246 6503
rect 4200 6431 4246 6469
rect 4200 6397 4206 6431
rect 4240 6397 4246 6431
rect 4200 6359 4246 6397
rect 4200 6325 4206 6359
rect 4240 6325 4246 6359
rect 4200 6287 4246 6325
rect 4200 6253 4206 6287
rect 4240 6253 4246 6287
rect 4200 6215 4246 6253
rect 4200 6181 4206 6215
rect 4240 6181 4246 6215
rect 4200 6143 4246 6181
rect 4200 6109 4206 6143
rect 4240 6109 4246 6143
rect 4200 6071 4246 6109
rect 4200 6037 4206 6071
rect 4240 6037 4246 6071
rect 4200 5999 4246 6037
rect 4200 5965 4206 5999
rect 4240 5965 4246 5999
rect 4200 5927 4246 5965
rect 4200 5893 4206 5927
rect 4240 5893 4246 5927
rect 4200 5855 4246 5893
rect 4200 5821 4206 5855
rect 4240 5821 4246 5855
rect 4200 5783 4246 5821
rect 4200 5749 4206 5783
rect 4240 5749 4246 5783
rect 4200 5711 4246 5749
rect 4200 5677 4206 5711
rect 4240 5677 4246 5711
rect 4200 5639 4246 5677
rect 4200 5605 4206 5639
rect 4240 5605 4246 5639
rect 4200 5590 4246 5605
rect 4296 6575 4342 6590
rect 4296 6541 4302 6575
rect 4336 6541 4342 6575
rect 4296 6503 4342 6541
rect 4296 6469 4302 6503
rect 4336 6469 4342 6503
rect 4296 6431 4342 6469
rect 4296 6397 4302 6431
rect 4336 6397 4342 6431
rect 4296 6359 4342 6397
rect 4296 6325 4302 6359
rect 4336 6325 4342 6359
rect 4296 6287 4342 6325
rect 4296 6253 4302 6287
rect 4336 6253 4342 6287
rect 4296 6215 4342 6253
rect 4296 6181 4302 6215
rect 4336 6181 4342 6215
rect 4296 6143 4342 6181
rect 4296 6109 4302 6143
rect 4336 6109 4342 6143
rect 4296 6071 4342 6109
rect 4296 6037 4302 6071
rect 4336 6037 4342 6071
rect 4296 5999 4342 6037
rect 4296 5965 4302 5999
rect 4336 5965 4342 5999
rect 4296 5927 4342 5965
rect 4296 5893 4302 5927
rect 4336 5893 4342 5927
rect 4296 5855 4342 5893
rect 4296 5821 4302 5855
rect 4336 5821 4342 5855
rect 4296 5783 4342 5821
rect 4296 5749 4302 5783
rect 4336 5749 4342 5783
rect 4296 5711 4342 5749
rect 4296 5677 4302 5711
rect 4336 5677 4342 5711
rect 4296 5639 4342 5677
rect 4296 5605 4302 5639
rect 4336 5605 4342 5639
rect 4296 5590 4342 5605
rect 4910 6571 4956 6586
rect 4910 6537 4916 6571
rect 4950 6537 4956 6571
rect 4910 6499 4956 6537
rect 4910 6465 4916 6499
rect 4950 6465 4956 6499
rect 4910 6427 4956 6465
rect 4910 6393 4916 6427
rect 4950 6393 4956 6427
rect 4910 6355 4956 6393
rect 4910 6321 4916 6355
rect 4950 6321 4956 6355
rect 4910 6283 4956 6321
rect 4910 6249 4916 6283
rect 4950 6249 4956 6283
rect 4910 6211 4956 6249
rect 4910 6177 4916 6211
rect 4950 6177 4956 6211
rect 4910 6139 4956 6177
rect 4910 6105 4916 6139
rect 4950 6105 4956 6139
rect 4910 6067 4956 6105
rect 4910 6033 4916 6067
rect 4950 6033 4956 6067
rect 4910 5995 4956 6033
rect 4910 5961 4916 5995
rect 4950 5961 4956 5995
rect 4910 5923 4956 5961
rect 4910 5889 4916 5923
rect 4950 5889 4956 5923
rect 4910 5851 4956 5889
rect 4910 5817 4916 5851
rect 4950 5817 4956 5851
rect 4910 5779 4956 5817
rect 4910 5745 4916 5779
rect 4950 5745 4956 5779
rect 4910 5707 4956 5745
rect 4910 5673 4916 5707
rect 4950 5673 4956 5707
rect 4910 5635 4956 5673
rect 4910 5601 4916 5635
rect 4950 5601 4956 5635
rect 4910 5586 4956 5601
rect 5006 6571 5052 6586
rect 5006 6537 5012 6571
rect 5046 6537 5052 6571
rect 5006 6499 5052 6537
rect 5006 6465 5012 6499
rect 5046 6465 5052 6499
rect 5006 6427 5052 6465
rect 5006 6393 5012 6427
rect 5046 6393 5052 6427
rect 5006 6355 5052 6393
rect 5006 6321 5012 6355
rect 5046 6321 5052 6355
rect 5006 6283 5052 6321
rect 5006 6249 5012 6283
rect 5046 6249 5052 6283
rect 5006 6211 5052 6249
rect 5006 6177 5012 6211
rect 5046 6177 5052 6211
rect 5006 6139 5052 6177
rect 5006 6105 5012 6139
rect 5046 6105 5052 6139
rect 5006 6067 5052 6105
rect 5006 6033 5012 6067
rect 5046 6033 5052 6067
rect 5006 5995 5052 6033
rect 5006 5961 5012 5995
rect 5046 5961 5052 5995
rect 5006 5923 5052 5961
rect 5006 5889 5012 5923
rect 5046 5889 5052 5923
rect 5006 5851 5052 5889
rect 5006 5817 5012 5851
rect 5046 5817 5052 5851
rect 5006 5779 5052 5817
rect 5006 5745 5012 5779
rect 5046 5745 5052 5779
rect 5006 5707 5052 5745
rect 5006 5673 5012 5707
rect 5046 5673 5052 5707
rect 5006 5635 5052 5673
rect 5006 5601 5012 5635
rect 5046 5601 5052 5635
rect 5006 5586 5052 5601
rect 5102 6571 5148 6586
rect 5102 6537 5108 6571
rect 5142 6537 5148 6571
rect 5102 6499 5148 6537
rect 5102 6465 5108 6499
rect 5142 6465 5148 6499
rect 5102 6427 5148 6465
rect 5102 6393 5108 6427
rect 5142 6393 5148 6427
rect 5102 6355 5148 6393
rect 5102 6321 5108 6355
rect 5142 6321 5148 6355
rect 5102 6283 5148 6321
rect 5102 6249 5108 6283
rect 5142 6249 5148 6283
rect 5102 6211 5148 6249
rect 5102 6177 5108 6211
rect 5142 6177 5148 6211
rect 5102 6139 5148 6177
rect 5102 6105 5108 6139
rect 5142 6105 5148 6139
rect 5102 6067 5148 6105
rect 5102 6033 5108 6067
rect 5142 6033 5148 6067
rect 5102 5995 5148 6033
rect 5102 5961 5108 5995
rect 5142 5961 5148 5995
rect 5102 5923 5148 5961
rect 5102 5889 5108 5923
rect 5142 5889 5148 5923
rect 5102 5851 5148 5889
rect 5102 5817 5108 5851
rect 5142 5817 5148 5851
rect 5102 5779 5148 5817
rect 5102 5745 5108 5779
rect 5142 5745 5148 5779
rect 5102 5707 5148 5745
rect 5102 5673 5108 5707
rect 5142 5673 5148 5707
rect 5102 5635 5148 5673
rect 5102 5601 5108 5635
rect 5142 5601 5148 5635
rect 5102 5586 5148 5601
rect 5198 6571 5244 6586
rect 5198 6537 5204 6571
rect 5238 6537 5244 6571
rect 5198 6499 5244 6537
rect 5198 6465 5204 6499
rect 5238 6465 5244 6499
rect 5198 6427 5244 6465
rect 5198 6393 5204 6427
rect 5238 6393 5244 6427
rect 5198 6355 5244 6393
rect 5198 6321 5204 6355
rect 5238 6321 5244 6355
rect 5198 6283 5244 6321
rect 5198 6249 5204 6283
rect 5238 6249 5244 6283
rect 5198 6211 5244 6249
rect 5198 6177 5204 6211
rect 5238 6177 5244 6211
rect 5198 6139 5244 6177
rect 5198 6105 5204 6139
rect 5238 6105 5244 6139
rect 5198 6067 5244 6105
rect 5198 6033 5204 6067
rect 5238 6033 5244 6067
rect 5198 5995 5244 6033
rect 5198 5961 5204 5995
rect 5238 5961 5244 5995
rect 5198 5923 5244 5961
rect 5198 5889 5204 5923
rect 5238 5889 5244 5923
rect 5198 5851 5244 5889
rect 5198 5817 5204 5851
rect 5238 5817 5244 5851
rect 5198 5779 5244 5817
rect 5198 5745 5204 5779
rect 5238 5745 5244 5779
rect 5198 5707 5244 5745
rect 5198 5673 5204 5707
rect 5238 5673 5244 5707
rect 5198 5635 5244 5673
rect 5198 5601 5204 5635
rect 5238 5601 5244 5635
rect 5198 5586 5244 5601
rect 5294 6571 5340 6586
rect 5294 6537 5300 6571
rect 5334 6537 5340 6571
rect 5294 6499 5340 6537
rect 5294 6465 5300 6499
rect 5334 6465 5340 6499
rect 5294 6427 5340 6465
rect 5294 6393 5300 6427
rect 5334 6393 5340 6427
rect 5294 6355 5340 6393
rect 5294 6321 5300 6355
rect 5334 6321 5340 6355
rect 5294 6283 5340 6321
rect 5294 6249 5300 6283
rect 5334 6249 5340 6283
rect 5294 6211 5340 6249
rect 5294 6177 5300 6211
rect 5334 6177 5340 6211
rect 5294 6139 5340 6177
rect 5294 6105 5300 6139
rect 5334 6105 5340 6139
rect 5294 6067 5340 6105
rect 5294 6033 5300 6067
rect 5334 6033 5340 6067
rect 5294 5995 5340 6033
rect 5294 5961 5300 5995
rect 5334 5961 5340 5995
rect 5294 5923 5340 5961
rect 5294 5889 5300 5923
rect 5334 5889 5340 5923
rect 5294 5851 5340 5889
rect 5294 5817 5300 5851
rect 5334 5817 5340 5851
rect 5294 5779 5340 5817
rect 5294 5745 5300 5779
rect 5334 5745 5340 5779
rect 5294 5707 5340 5745
rect 5294 5673 5300 5707
rect 5334 5673 5340 5707
rect 5294 5635 5340 5673
rect 5294 5601 5300 5635
rect 5334 5601 5340 5635
rect 5294 5586 5340 5601
rect 5390 6571 5436 6586
rect 5390 6537 5396 6571
rect 5430 6537 5436 6571
rect 5390 6499 5436 6537
rect 5390 6465 5396 6499
rect 5430 6465 5436 6499
rect 5390 6427 5436 6465
rect 5390 6393 5396 6427
rect 5430 6393 5436 6427
rect 5390 6355 5436 6393
rect 5390 6321 5396 6355
rect 5430 6321 5436 6355
rect 5390 6283 5436 6321
rect 5390 6249 5396 6283
rect 5430 6249 5436 6283
rect 5390 6211 5436 6249
rect 5390 6177 5396 6211
rect 5430 6177 5436 6211
rect 5390 6139 5436 6177
rect 5390 6105 5396 6139
rect 5430 6105 5436 6139
rect 5390 6067 5436 6105
rect 5390 6033 5396 6067
rect 5430 6033 5436 6067
rect 5390 5995 5436 6033
rect 5390 5961 5396 5995
rect 5430 5961 5436 5995
rect 5390 5923 5436 5961
rect 5390 5889 5396 5923
rect 5430 5889 5436 5923
rect 5390 5851 5436 5889
rect 5390 5817 5396 5851
rect 5430 5817 5436 5851
rect 5390 5779 5436 5817
rect 5390 5745 5396 5779
rect 5430 5745 5436 5779
rect 5390 5707 5436 5745
rect 5390 5673 5396 5707
rect 5430 5673 5436 5707
rect 5390 5635 5436 5673
rect 5390 5601 5396 5635
rect 5430 5601 5436 5635
rect 5390 5586 5436 5601
rect 5486 6571 5532 6586
rect 5486 6537 5492 6571
rect 5526 6537 5532 6571
rect 5486 6499 5532 6537
rect 5486 6465 5492 6499
rect 5526 6465 5532 6499
rect 5486 6427 5532 6465
rect 5486 6393 5492 6427
rect 5526 6393 5532 6427
rect 5486 6355 5532 6393
rect 5486 6321 5492 6355
rect 5526 6321 5532 6355
rect 5486 6283 5532 6321
rect 5486 6249 5492 6283
rect 5526 6249 5532 6283
rect 5486 6211 5532 6249
rect 5486 6177 5492 6211
rect 5526 6177 5532 6211
rect 5486 6139 5532 6177
rect 5486 6105 5492 6139
rect 5526 6105 5532 6139
rect 5486 6067 5532 6105
rect 5486 6033 5492 6067
rect 5526 6033 5532 6067
rect 5486 5995 5532 6033
rect 5486 5961 5492 5995
rect 5526 5961 5532 5995
rect 5486 5923 5532 5961
rect 5486 5889 5492 5923
rect 5526 5889 5532 5923
rect 5486 5851 5532 5889
rect 5486 5817 5492 5851
rect 5526 5817 5532 5851
rect 5486 5779 5532 5817
rect 5486 5745 5492 5779
rect 5526 5745 5532 5779
rect 5486 5707 5532 5745
rect 5486 5673 5492 5707
rect 5526 5673 5532 5707
rect 5486 5635 5532 5673
rect 5486 5601 5492 5635
rect 5526 5601 5532 5635
rect 5486 5586 5532 5601
rect 5582 6571 5628 6586
rect 5582 6537 5588 6571
rect 5622 6537 5628 6571
rect 5582 6499 5628 6537
rect 5582 6465 5588 6499
rect 5622 6465 5628 6499
rect 5582 6427 5628 6465
rect 5582 6393 5588 6427
rect 5622 6393 5628 6427
rect 5582 6355 5628 6393
rect 5582 6321 5588 6355
rect 5622 6321 5628 6355
rect 5582 6283 5628 6321
rect 5582 6249 5588 6283
rect 5622 6249 5628 6283
rect 5582 6211 5628 6249
rect 5582 6177 5588 6211
rect 5622 6177 5628 6211
rect 5582 6139 5628 6177
rect 5582 6105 5588 6139
rect 5622 6105 5628 6139
rect 5582 6067 5628 6105
rect 5582 6033 5588 6067
rect 5622 6033 5628 6067
rect 5582 5995 5628 6033
rect 5582 5961 5588 5995
rect 5622 5961 5628 5995
rect 5582 5923 5628 5961
rect 5582 5889 5588 5923
rect 5622 5889 5628 5923
rect 5582 5851 5628 5889
rect 5582 5817 5588 5851
rect 5622 5817 5628 5851
rect 5582 5779 5628 5817
rect 5582 5745 5588 5779
rect 5622 5745 5628 5779
rect 5582 5707 5628 5745
rect 5582 5673 5588 5707
rect 5622 5673 5628 5707
rect 5582 5635 5628 5673
rect 5582 5601 5588 5635
rect 5622 5601 5628 5635
rect 5582 5586 5628 5601
rect 5678 6571 5724 6586
rect 5678 6537 5684 6571
rect 5718 6537 5724 6571
rect 5678 6499 5724 6537
rect 5678 6465 5684 6499
rect 5718 6465 5724 6499
rect 5678 6427 5724 6465
rect 5678 6393 5684 6427
rect 5718 6393 5724 6427
rect 5678 6355 5724 6393
rect 5678 6321 5684 6355
rect 5718 6321 5724 6355
rect 5678 6283 5724 6321
rect 5678 6249 5684 6283
rect 5718 6249 5724 6283
rect 5678 6211 5724 6249
rect 5678 6177 5684 6211
rect 5718 6177 5724 6211
rect 5678 6139 5724 6177
rect 5678 6105 5684 6139
rect 5718 6105 5724 6139
rect 5678 6067 5724 6105
rect 5678 6033 5684 6067
rect 5718 6033 5724 6067
rect 5678 5995 5724 6033
rect 5678 5961 5684 5995
rect 5718 5961 5724 5995
rect 5678 5923 5724 5961
rect 5678 5889 5684 5923
rect 5718 5889 5724 5923
rect 5678 5851 5724 5889
rect 5678 5817 5684 5851
rect 5718 5817 5724 5851
rect 5678 5779 5724 5817
rect 5678 5745 5684 5779
rect 5718 5745 5724 5779
rect 5678 5707 5724 5745
rect 5678 5673 5684 5707
rect 5718 5673 5724 5707
rect 5678 5635 5724 5673
rect 5678 5601 5684 5635
rect 5718 5601 5724 5635
rect 5678 5586 5724 5601
rect 6174 6575 6220 6590
rect 6174 6541 6180 6575
rect 6214 6541 6220 6575
rect 6174 6503 6220 6541
rect 6174 6469 6180 6503
rect 6214 6469 6220 6503
rect 6174 6431 6220 6469
rect 6174 6397 6180 6431
rect 6214 6397 6220 6431
rect 6174 6359 6220 6397
rect 6174 6325 6180 6359
rect 6214 6325 6220 6359
rect 6174 6287 6220 6325
rect 6174 6253 6180 6287
rect 6214 6253 6220 6287
rect 6174 6215 6220 6253
rect 6174 6181 6180 6215
rect 6214 6181 6220 6215
rect 6174 6143 6220 6181
rect 6174 6109 6180 6143
rect 6214 6109 6220 6143
rect 6174 6071 6220 6109
rect 6174 6037 6180 6071
rect 6214 6037 6220 6071
rect 6174 5999 6220 6037
rect 6174 5965 6180 5999
rect 6214 5965 6220 5999
rect 6174 5927 6220 5965
rect 6174 5893 6180 5927
rect 6214 5893 6220 5927
rect 6174 5855 6220 5893
rect 6174 5821 6180 5855
rect 6214 5821 6220 5855
rect 6174 5783 6220 5821
rect 6174 5749 6180 5783
rect 6214 5749 6220 5783
rect 6174 5711 6220 5749
rect 6174 5677 6180 5711
rect 6214 5677 6220 5711
rect 6174 5639 6220 5677
rect 6174 5605 6180 5639
rect 6214 5605 6220 5639
rect 6174 5590 6220 5605
rect 6270 6575 6316 6590
rect 6270 6541 6276 6575
rect 6310 6541 6316 6575
rect 6270 6503 6316 6541
rect 6270 6469 6276 6503
rect 6310 6469 6316 6503
rect 6270 6431 6316 6469
rect 6270 6397 6276 6431
rect 6310 6397 6316 6431
rect 6270 6359 6316 6397
rect 6270 6325 6276 6359
rect 6310 6325 6316 6359
rect 6270 6287 6316 6325
rect 6270 6253 6276 6287
rect 6310 6253 6316 6287
rect 6270 6215 6316 6253
rect 6270 6181 6276 6215
rect 6310 6181 6316 6215
rect 6270 6143 6316 6181
rect 6270 6109 6276 6143
rect 6310 6109 6316 6143
rect 6270 6071 6316 6109
rect 6270 6037 6276 6071
rect 6310 6037 6316 6071
rect 6270 5999 6316 6037
rect 6270 5965 6276 5999
rect 6310 5965 6316 5999
rect 6270 5927 6316 5965
rect 6270 5893 6276 5927
rect 6310 5893 6316 5927
rect 6270 5855 6316 5893
rect 6270 5821 6276 5855
rect 6310 5821 6316 5855
rect 6270 5783 6316 5821
rect 6270 5749 6276 5783
rect 6310 5749 6316 5783
rect 6270 5711 6316 5749
rect 6270 5677 6276 5711
rect 6310 5677 6316 5711
rect 6270 5639 6316 5677
rect 6270 5605 6276 5639
rect 6310 5605 6316 5639
rect 6270 5590 6316 5605
rect 6366 6575 6412 6590
rect 6366 6541 6372 6575
rect 6406 6541 6412 6575
rect 6366 6503 6412 6541
rect 6366 6469 6372 6503
rect 6406 6469 6412 6503
rect 6366 6431 6412 6469
rect 6366 6397 6372 6431
rect 6406 6397 6412 6431
rect 6366 6359 6412 6397
rect 6366 6325 6372 6359
rect 6406 6325 6412 6359
rect 6366 6287 6412 6325
rect 6366 6253 6372 6287
rect 6406 6253 6412 6287
rect 6366 6215 6412 6253
rect 6366 6181 6372 6215
rect 6406 6181 6412 6215
rect 6366 6143 6412 6181
rect 6366 6109 6372 6143
rect 6406 6109 6412 6143
rect 6366 6071 6412 6109
rect 6366 6037 6372 6071
rect 6406 6037 6412 6071
rect 6366 5999 6412 6037
rect 6366 5965 6372 5999
rect 6406 5965 6412 5999
rect 6366 5927 6412 5965
rect 6366 5893 6372 5927
rect 6406 5893 6412 5927
rect 6366 5855 6412 5893
rect 6366 5821 6372 5855
rect 6406 5821 6412 5855
rect 6366 5783 6412 5821
rect 6366 5749 6372 5783
rect 6406 5749 6412 5783
rect 6366 5711 6412 5749
rect 6366 5677 6372 5711
rect 6406 5677 6412 5711
rect 6366 5639 6412 5677
rect 6366 5605 6372 5639
rect 6406 5605 6412 5639
rect 6366 5590 6412 5605
rect 6462 6575 6508 6590
rect 6462 6541 6468 6575
rect 6502 6541 6508 6575
rect 6462 6503 6508 6541
rect 6462 6469 6468 6503
rect 6502 6469 6508 6503
rect 6462 6431 6508 6469
rect 6462 6397 6468 6431
rect 6502 6397 6508 6431
rect 6462 6359 6508 6397
rect 6462 6325 6468 6359
rect 6502 6325 6508 6359
rect 6462 6287 6508 6325
rect 6462 6253 6468 6287
rect 6502 6253 6508 6287
rect 6462 6215 6508 6253
rect 6462 6181 6468 6215
rect 6502 6181 6508 6215
rect 6462 6143 6508 6181
rect 6462 6109 6468 6143
rect 6502 6109 6508 6143
rect 6462 6071 6508 6109
rect 6462 6037 6468 6071
rect 6502 6037 6508 6071
rect 6462 5999 6508 6037
rect 6462 5965 6468 5999
rect 6502 5965 6508 5999
rect 6462 5927 6508 5965
rect 6462 5893 6468 5927
rect 6502 5893 6508 5927
rect 6462 5855 6508 5893
rect 6462 5821 6468 5855
rect 6502 5821 6508 5855
rect 6462 5783 6508 5821
rect 6462 5749 6468 5783
rect 6502 5749 6508 5783
rect 6462 5711 6508 5749
rect 6462 5677 6468 5711
rect 6502 5677 6508 5711
rect 6462 5639 6508 5677
rect 6462 5605 6468 5639
rect 6502 5605 6508 5639
rect 6462 5590 6508 5605
rect 6558 6575 6604 6590
rect 6558 6541 6564 6575
rect 6598 6541 6604 6575
rect 6558 6503 6604 6541
rect 6558 6469 6564 6503
rect 6598 6469 6604 6503
rect 6558 6431 6604 6469
rect 6558 6397 6564 6431
rect 6598 6397 6604 6431
rect 6558 6359 6604 6397
rect 6558 6325 6564 6359
rect 6598 6325 6604 6359
rect 6558 6287 6604 6325
rect 6558 6253 6564 6287
rect 6598 6253 6604 6287
rect 6558 6215 6604 6253
rect 6558 6181 6564 6215
rect 6598 6181 6604 6215
rect 6558 6143 6604 6181
rect 6558 6109 6564 6143
rect 6598 6109 6604 6143
rect 6558 6071 6604 6109
rect 6558 6037 6564 6071
rect 6598 6037 6604 6071
rect 6558 5999 6604 6037
rect 6558 5965 6564 5999
rect 6598 5965 6604 5999
rect 6558 5927 6604 5965
rect 6558 5893 6564 5927
rect 6598 5893 6604 5927
rect 6558 5855 6604 5893
rect 6558 5821 6564 5855
rect 6598 5821 6604 5855
rect 6558 5783 6604 5821
rect 6558 5749 6564 5783
rect 6598 5749 6604 5783
rect 6558 5711 6604 5749
rect 6558 5677 6564 5711
rect 6598 5677 6604 5711
rect 6558 5639 6604 5677
rect 6558 5605 6564 5639
rect 6598 5605 6604 5639
rect 6558 5590 6604 5605
rect 6654 6575 6700 6590
rect 6654 6541 6660 6575
rect 6694 6541 6700 6575
rect 6654 6503 6700 6541
rect 6654 6469 6660 6503
rect 6694 6469 6700 6503
rect 6654 6431 6700 6469
rect 6654 6397 6660 6431
rect 6694 6397 6700 6431
rect 6654 6359 6700 6397
rect 6654 6325 6660 6359
rect 6694 6325 6700 6359
rect 6654 6287 6700 6325
rect 6654 6253 6660 6287
rect 6694 6253 6700 6287
rect 6654 6215 6700 6253
rect 6654 6181 6660 6215
rect 6694 6181 6700 6215
rect 6654 6143 6700 6181
rect 6654 6109 6660 6143
rect 6694 6109 6700 6143
rect 6654 6071 6700 6109
rect 6654 6037 6660 6071
rect 6694 6037 6700 6071
rect 6654 5999 6700 6037
rect 6654 5965 6660 5999
rect 6694 5965 6700 5999
rect 6654 5927 6700 5965
rect 6654 5893 6660 5927
rect 6694 5893 6700 5927
rect 6654 5855 6700 5893
rect 6654 5821 6660 5855
rect 6694 5821 6700 5855
rect 6654 5783 6700 5821
rect 6654 5749 6660 5783
rect 6694 5749 6700 5783
rect 6654 5711 6700 5749
rect 6654 5677 6660 5711
rect 6694 5677 6700 5711
rect 6654 5639 6700 5677
rect 6654 5605 6660 5639
rect 6694 5605 6700 5639
rect 6654 5590 6700 5605
rect 6750 6575 6796 6590
rect 6750 6541 6756 6575
rect 6790 6541 6796 6575
rect 6750 6503 6796 6541
rect 6750 6469 6756 6503
rect 6790 6469 6796 6503
rect 6750 6431 6796 6469
rect 6750 6397 6756 6431
rect 6790 6397 6796 6431
rect 6750 6359 6796 6397
rect 6750 6325 6756 6359
rect 6790 6325 6796 6359
rect 6750 6287 6796 6325
rect 6750 6253 6756 6287
rect 6790 6253 6796 6287
rect 6750 6215 6796 6253
rect 6750 6181 6756 6215
rect 6790 6181 6796 6215
rect 6750 6143 6796 6181
rect 6750 6109 6756 6143
rect 6790 6109 6796 6143
rect 6750 6071 6796 6109
rect 6750 6037 6756 6071
rect 6790 6037 6796 6071
rect 6750 5999 6796 6037
rect 6750 5965 6756 5999
rect 6790 5965 6796 5999
rect 6750 5927 6796 5965
rect 6750 5893 6756 5927
rect 6790 5893 6796 5927
rect 6750 5855 6796 5893
rect 6750 5821 6756 5855
rect 6790 5821 6796 5855
rect 6750 5783 6796 5821
rect 6750 5749 6756 5783
rect 6790 5749 6796 5783
rect 6750 5711 6796 5749
rect 6750 5677 6756 5711
rect 6790 5677 6796 5711
rect 6750 5639 6796 5677
rect 6750 5605 6756 5639
rect 6790 5605 6796 5639
rect 6750 5590 6796 5605
rect 6846 6575 6892 6590
rect 6846 6541 6852 6575
rect 6886 6541 6892 6575
rect 6846 6503 6892 6541
rect 6846 6469 6852 6503
rect 6886 6469 6892 6503
rect 6846 6431 6892 6469
rect 6846 6397 6852 6431
rect 6886 6397 6892 6431
rect 6846 6359 6892 6397
rect 6846 6325 6852 6359
rect 6886 6325 6892 6359
rect 6846 6287 6892 6325
rect 6846 6253 6852 6287
rect 6886 6253 6892 6287
rect 6846 6215 6892 6253
rect 6846 6181 6852 6215
rect 6886 6181 6892 6215
rect 6846 6143 6892 6181
rect 6846 6109 6852 6143
rect 6886 6109 6892 6143
rect 6846 6071 6892 6109
rect 6846 6037 6852 6071
rect 6886 6037 6892 6071
rect 6846 5999 6892 6037
rect 6846 5965 6852 5999
rect 6886 5965 6892 5999
rect 6846 5927 6892 5965
rect 6846 5893 6852 5927
rect 6886 5893 6892 5927
rect 6846 5855 6892 5893
rect 6846 5821 6852 5855
rect 6886 5821 6892 5855
rect 6846 5783 6892 5821
rect 6846 5749 6852 5783
rect 6886 5749 6892 5783
rect 6846 5711 6892 5749
rect 6846 5677 6852 5711
rect 6886 5677 6892 5711
rect 6846 5639 6892 5677
rect 6846 5605 6852 5639
rect 6886 5605 6892 5639
rect 6846 5590 6892 5605
rect 6942 6575 6988 6590
rect 6942 6541 6948 6575
rect 6982 6541 6988 6575
rect 6942 6503 6988 6541
rect 6942 6469 6948 6503
rect 6982 6469 6988 6503
rect 6942 6431 6988 6469
rect 6942 6397 6948 6431
rect 6982 6397 6988 6431
rect 6942 6359 6988 6397
rect 6942 6325 6948 6359
rect 6982 6325 6988 6359
rect 6942 6287 6988 6325
rect 6942 6253 6948 6287
rect 6982 6253 6988 6287
rect 6942 6215 6988 6253
rect 6942 6181 6948 6215
rect 6982 6181 6988 6215
rect 6942 6143 6988 6181
rect 6942 6109 6948 6143
rect 6982 6109 6988 6143
rect 6942 6071 6988 6109
rect 6942 6037 6948 6071
rect 6982 6037 6988 6071
rect 6942 5999 6988 6037
rect 6942 5965 6948 5999
rect 6982 5965 6988 5999
rect 6942 5927 6988 5965
rect 6942 5893 6948 5927
rect 6982 5893 6988 5927
rect 6942 5855 6988 5893
rect 6942 5821 6948 5855
rect 6982 5821 6988 5855
rect 6942 5783 6988 5821
rect 6942 5749 6948 5783
rect 6982 5749 6988 5783
rect 6942 5711 6988 5749
rect 6942 5677 6948 5711
rect 6982 5677 6988 5711
rect 6942 5639 6988 5677
rect 6942 5605 6948 5639
rect 6982 5605 6988 5639
rect 6942 5590 6988 5605
rect 7038 6575 7084 6590
rect 7038 6541 7044 6575
rect 7078 6541 7084 6575
rect 7038 6503 7084 6541
rect 7038 6469 7044 6503
rect 7078 6469 7084 6503
rect 7038 6431 7084 6469
rect 7038 6397 7044 6431
rect 7078 6397 7084 6431
rect 7038 6359 7084 6397
rect 7038 6325 7044 6359
rect 7078 6325 7084 6359
rect 7038 6287 7084 6325
rect 7038 6253 7044 6287
rect 7078 6253 7084 6287
rect 7038 6215 7084 6253
rect 7038 6181 7044 6215
rect 7078 6181 7084 6215
rect 7038 6143 7084 6181
rect 7038 6109 7044 6143
rect 7078 6109 7084 6143
rect 7038 6071 7084 6109
rect 7038 6037 7044 6071
rect 7078 6037 7084 6071
rect 7038 5999 7084 6037
rect 7038 5965 7044 5999
rect 7078 5965 7084 5999
rect 7038 5927 7084 5965
rect 7038 5893 7044 5927
rect 7078 5893 7084 5927
rect 7038 5855 7084 5893
rect 7038 5821 7044 5855
rect 7078 5821 7084 5855
rect 7038 5783 7084 5821
rect 7038 5749 7044 5783
rect 7078 5749 7084 5783
rect 7038 5711 7084 5749
rect 7038 5677 7044 5711
rect 7078 5677 7084 5711
rect 7038 5639 7084 5677
rect 7038 5605 7044 5639
rect 7078 5605 7084 5639
rect 7038 5590 7084 5605
rect 7134 6575 7180 6590
rect 7134 6541 7140 6575
rect 7174 6541 7180 6575
rect 7134 6503 7180 6541
rect 7134 6469 7140 6503
rect 7174 6469 7180 6503
rect 7134 6431 7180 6469
rect 7134 6397 7140 6431
rect 7174 6397 7180 6431
rect 7134 6359 7180 6397
rect 7134 6325 7140 6359
rect 7174 6325 7180 6359
rect 7134 6287 7180 6325
rect 7134 6253 7140 6287
rect 7174 6253 7180 6287
rect 7134 6215 7180 6253
rect 7134 6181 7140 6215
rect 7174 6181 7180 6215
rect 7134 6143 7180 6181
rect 7134 6109 7140 6143
rect 7174 6109 7180 6143
rect 7134 6071 7180 6109
rect 7134 6037 7140 6071
rect 7174 6037 7180 6071
rect 7134 5999 7180 6037
rect 7134 5965 7140 5999
rect 7174 5965 7180 5999
rect 7134 5927 7180 5965
rect 7134 5893 7140 5927
rect 7174 5893 7180 5927
rect 7134 5855 7180 5893
rect 7134 5821 7140 5855
rect 7174 5821 7180 5855
rect 7134 5783 7180 5821
rect 7134 5749 7140 5783
rect 7174 5749 7180 5783
rect 7134 5711 7180 5749
rect 7134 5677 7140 5711
rect 7174 5677 7180 5711
rect 7134 5639 7180 5677
rect 7134 5605 7140 5639
rect 7174 5605 7180 5639
rect 7134 5590 7180 5605
rect 7230 6575 7276 6590
rect 7230 6541 7236 6575
rect 7270 6541 7276 6575
rect 7230 6503 7276 6541
rect 7230 6469 7236 6503
rect 7270 6469 7276 6503
rect 7230 6431 7276 6469
rect 7230 6397 7236 6431
rect 7270 6397 7276 6431
rect 7230 6359 7276 6397
rect 7230 6325 7236 6359
rect 7270 6325 7276 6359
rect 7230 6287 7276 6325
rect 7230 6253 7236 6287
rect 7270 6253 7276 6287
rect 7230 6215 7276 6253
rect 7230 6181 7236 6215
rect 7270 6181 7276 6215
rect 7230 6143 7276 6181
rect 7230 6109 7236 6143
rect 7270 6109 7276 6143
rect 7230 6071 7276 6109
rect 7230 6037 7236 6071
rect 7270 6037 7276 6071
rect 7230 5999 7276 6037
rect 7230 5965 7236 5999
rect 7270 5965 7276 5999
rect 7230 5927 7276 5965
rect 7230 5893 7236 5927
rect 7270 5893 7276 5927
rect 7230 5855 7276 5893
rect 7230 5821 7236 5855
rect 7270 5821 7276 5855
rect 7230 5783 7276 5821
rect 7230 5749 7236 5783
rect 7270 5749 7276 5783
rect 7230 5711 7276 5749
rect 7230 5677 7236 5711
rect 7270 5677 7276 5711
rect 7230 5639 7276 5677
rect 7230 5605 7236 5639
rect 7270 5605 7276 5639
rect 7230 5590 7276 5605
rect 7326 6575 7372 6590
rect 7326 6541 7332 6575
rect 7366 6541 7372 6575
rect 7326 6503 7372 6541
rect 7326 6469 7332 6503
rect 7366 6469 7372 6503
rect 7326 6431 7372 6469
rect 7326 6397 7332 6431
rect 7366 6397 7372 6431
rect 7326 6359 7372 6397
rect 7326 6325 7332 6359
rect 7366 6325 7372 6359
rect 7326 6287 7372 6325
rect 7326 6253 7332 6287
rect 7366 6253 7372 6287
rect 7326 6215 7372 6253
rect 7326 6181 7332 6215
rect 7366 6181 7372 6215
rect 7326 6143 7372 6181
rect 7326 6109 7332 6143
rect 7366 6109 7372 6143
rect 7326 6071 7372 6109
rect 7326 6037 7332 6071
rect 7366 6037 7372 6071
rect 7326 5999 7372 6037
rect 7326 5965 7332 5999
rect 7366 5965 7372 5999
rect 7326 5927 7372 5965
rect 7326 5893 7332 5927
rect 7366 5893 7372 5927
rect 7326 5855 7372 5893
rect 7326 5821 7332 5855
rect 7366 5821 7372 5855
rect 7326 5783 7372 5821
rect 7326 5749 7332 5783
rect 7366 5749 7372 5783
rect 7326 5711 7372 5749
rect 7326 5677 7332 5711
rect 7366 5677 7372 5711
rect 7326 5639 7372 5677
rect 7326 5605 7332 5639
rect 7366 5605 7372 5639
rect 7326 5590 7372 5605
rect 7940 6571 7986 6586
rect 7940 6537 7946 6571
rect 7980 6537 7986 6571
rect 7940 6499 7986 6537
rect 7940 6465 7946 6499
rect 7980 6465 7986 6499
rect 7940 6427 7986 6465
rect 7940 6393 7946 6427
rect 7980 6393 7986 6427
rect 7940 6355 7986 6393
rect 7940 6321 7946 6355
rect 7980 6321 7986 6355
rect 7940 6283 7986 6321
rect 7940 6249 7946 6283
rect 7980 6249 7986 6283
rect 7940 6211 7986 6249
rect 7940 6177 7946 6211
rect 7980 6177 7986 6211
rect 7940 6139 7986 6177
rect 7940 6105 7946 6139
rect 7980 6105 7986 6139
rect 7940 6067 7986 6105
rect 7940 6033 7946 6067
rect 7980 6033 7986 6067
rect 7940 5995 7986 6033
rect 7940 5961 7946 5995
rect 7980 5961 7986 5995
rect 7940 5923 7986 5961
rect 7940 5889 7946 5923
rect 7980 5889 7986 5923
rect 7940 5851 7986 5889
rect 7940 5817 7946 5851
rect 7980 5817 7986 5851
rect 7940 5779 7986 5817
rect 7940 5745 7946 5779
rect 7980 5745 7986 5779
rect 7940 5707 7986 5745
rect 7940 5673 7946 5707
rect 7980 5673 7986 5707
rect 7940 5635 7986 5673
rect 7940 5601 7946 5635
rect 7980 5601 7986 5635
rect 7940 5586 7986 5601
rect 8036 6571 8082 6586
rect 8036 6537 8042 6571
rect 8076 6537 8082 6571
rect 8036 6499 8082 6537
rect 8036 6465 8042 6499
rect 8076 6465 8082 6499
rect 8036 6427 8082 6465
rect 8036 6393 8042 6427
rect 8076 6393 8082 6427
rect 8036 6355 8082 6393
rect 8036 6321 8042 6355
rect 8076 6321 8082 6355
rect 8036 6283 8082 6321
rect 8036 6249 8042 6283
rect 8076 6249 8082 6283
rect 8036 6211 8082 6249
rect 8036 6177 8042 6211
rect 8076 6177 8082 6211
rect 8036 6139 8082 6177
rect 8036 6105 8042 6139
rect 8076 6105 8082 6139
rect 8036 6067 8082 6105
rect 8036 6033 8042 6067
rect 8076 6033 8082 6067
rect 8036 5995 8082 6033
rect 8036 5961 8042 5995
rect 8076 5961 8082 5995
rect 8036 5923 8082 5961
rect 8036 5889 8042 5923
rect 8076 5889 8082 5923
rect 8036 5851 8082 5889
rect 8036 5817 8042 5851
rect 8076 5817 8082 5851
rect 8036 5779 8082 5817
rect 8036 5745 8042 5779
rect 8076 5745 8082 5779
rect 8036 5707 8082 5745
rect 8036 5673 8042 5707
rect 8076 5673 8082 5707
rect 8036 5635 8082 5673
rect 8036 5601 8042 5635
rect 8076 5601 8082 5635
rect 8036 5586 8082 5601
rect 8132 6571 8178 6586
rect 8132 6537 8138 6571
rect 8172 6537 8178 6571
rect 8132 6499 8178 6537
rect 8132 6465 8138 6499
rect 8172 6465 8178 6499
rect 8132 6427 8178 6465
rect 8132 6393 8138 6427
rect 8172 6393 8178 6427
rect 8132 6355 8178 6393
rect 8132 6321 8138 6355
rect 8172 6321 8178 6355
rect 8132 6283 8178 6321
rect 8132 6249 8138 6283
rect 8172 6249 8178 6283
rect 8132 6211 8178 6249
rect 8132 6177 8138 6211
rect 8172 6177 8178 6211
rect 8132 6139 8178 6177
rect 8132 6105 8138 6139
rect 8172 6105 8178 6139
rect 8132 6067 8178 6105
rect 8132 6033 8138 6067
rect 8172 6033 8178 6067
rect 8132 5995 8178 6033
rect 8132 5961 8138 5995
rect 8172 5961 8178 5995
rect 8132 5923 8178 5961
rect 8132 5889 8138 5923
rect 8172 5889 8178 5923
rect 8132 5851 8178 5889
rect 8132 5817 8138 5851
rect 8172 5817 8178 5851
rect 8132 5779 8178 5817
rect 8132 5745 8138 5779
rect 8172 5745 8178 5779
rect 8132 5707 8178 5745
rect 8132 5673 8138 5707
rect 8172 5673 8178 5707
rect 8132 5635 8178 5673
rect 8132 5601 8138 5635
rect 8172 5601 8178 5635
rect 8132 5586 8178 5601
rect 8228 6571 8274 6586
rect 8228 6537 8234 6571
rect 8268 6537 8274 6571
rect 8228 6499 8274 6537
rect 8228 6465 8234 6499
rect 8268 6465 8274 6499
rect 8228 6427 8274 6465
rect 8228 6393 8234 6427
rect 8268 6393 8274 6427
rect 8228 6355 8274 6393
rect 8228 6321 8234 6355
rect 8268 6321 8274 6355
rect 8228 6283 8274 6321
rect 8228 6249 8234 6283
rect 8268 6249 8274 6283
rect 8228 6211 8274 6249
rect 8228 6177 8234 6211
rect 8268 6177 8274 6211
rect 8228 6139 8274 6177
rect 8228 6105 8234 6139
rect 8268 6105 8274 6139
rect 8228 6067 8274 6105
rect 8228 6033 8234 6067
rect 8268 6033 8274 6067
rect 8228 5995 8274 6033
rect 8228 5961 8234 5995
rect 8268 5961 8274 5995
rect 8228 5923 8274 5961
rect 8228 5889 8234 5923
rect 8268 5889 8274 5923
rect 8228 5851 8274 5889
rect 8228 5817 8234 5851
rect 8268 5817 8274 5851
rect 8228 5779 8274 5817
rect 8228 5745 8234 5779
rect 8268 5745 8274 5779
rect 8228 5707 8274 5745
rect 8228 5673 8234 5707
rect 8268 5673 8274 5707
rect 8228 5635 8274 5673
rect 8228 5601 8234 5635
rect 8268 5601 8274 5635
rect 8228 5586 8274 5601
rect 8324 6571 8370 6586
rect 8324 6537 8330 6571
rect 8364 6537 8370 6571
rect 8324 6499 8370 6537
rect 8324 6465 8330 6499
rect 8364 6465 8370 6499
rect 8324 6427 8370 6465
rect 8324 6393 8330 6427
rect 8364 6393 8370 6427
rect 8324 6355 8370 6393
rect 8324 6321 8330 6355
rect 8364 6321 8370 6355
rect 8324 6283 8370 6321
rect 8324 6249 8330 6283
rect 8364 6249 8370 6283
rect 8324 6211 8370 6249
rect 8324 6177 8330 6211
rect 8364 6177 8370 6211
rect 8324 6139 8370 6177
rect 8324 6105 8330 6139
rect 8364 6105 8370 6139
rect 8324 6067 8370 6105
rect 8324 6033 8330 6067
rect 8364 6033 8370 6067
rect 8324 5995 8370 6033
rect 8324 5961 8330 5995
rect 8364 5961 8370 5995
rect 8324 5923 8370 5961
rect 8324 5889 8330 5923
rect 8364 5889 8370 5923
rect 8324 5851 8370 5889
rect 8324 5817 8330 5851
rect 8364 5817 8370 5851
rect 8324 5779 8370 5817
rect 8324 5745 8330 5779
rect 8364 5745 8370 5779
rect 8324 5707 8370 5745
rect 8324 5673 8330 5707
rect 8364 5673 8370 5707
rect 8324 5635 8370 5673
rect 8324 5601 8330 5635
rect 8364 5601 8370 5635
rect 8324 5586 8370 5601
rect 8420 6571 8466 6586
rect 8420 6537 8426 6571
rect 8460 6537 8466 6571
rect 8420 6499 8466 6537
rect 8420 6465 8426 6499
rect 8460 6465 8466 6499
rect 8420 6427 8466 6465
rect 8420 6393 8426 6427
rect 8460 6393 8466 6427
rect 8420 6355 8466 6393
rect 8420 6321 8426 6355
rect 8460 6321 8466 6355
rect 8420 6283 8466 6321
rect 8420 6249 8426 6283
rect 8460 6249 8466 6283
rect 8420 6211 8466 6249
rect 8420 6177 8426 6211
rect 8460 6177 8466 6211
rect 8420 6139 8466 6177
rect 8420 6105 8426 6139
rect 8460 6105 8466 6139
rect 8420 6067 8466 6105
rect 8420 6033 8426 6067
rect 8460 6033 8466 6067
rect 8420 5995 8466 6033
rect 8420 5961 8426 5995
rect 8460 5961 8466 5995
rect 8420 5923 8466 5961
rect 8420 5889 8426 5923
rect 8460 5889 8466 5923
rect 8420 5851 8466 5889
rect 8420 5817 8426 5851
rect 8460 5817 8466 5851
rect 8420 5779 8466 5817
rect 8420 5745 8426 5779
rect 8460 5745 8466 5779
rect 8420 5707 8466 5745
rect 8420 5673 8426 5707
rect 8460 5673 8466 5707
rect 8420 5635 8466 5673
rect 8420 5601 8426 5635
rect 8460 5601 8466 5635
rect 8420 5586 8466 5601
rect 8516 6571 8562 6586
rect 8516 6537 8522 6571
rect 8556 6537 8562 6571
rect 8516 6499 8562 6537
rect 8516 6465 8522 6499
rect 8556 6465 8562 6499
rect 8516 6427 8562 6465
rect 8516 6393 8522 6427
rect 8556 6393 8562 6427
rect 8516 6355 8562 6393
rect 8516 6321 8522 6355
rect 8556 6321 8562 6355
rect 8516 6283 8562 6321
rect 8516 6249 8522 6283
rect 8556 6249 8562 6283
rect 8516 6211 8562 6249
rect 8516 6177 8522 6211
rect 8556 6177 8562 6211
rect 8516 6139 8562 6177
rect 8516 6105 8522 6139
rect 8556 6105 8562 6139
rect 8516 6067 8562 6105
rect 8516 6033 8522 6067
rect 8556 6033 8562 6067
rect 8516 5995 8562 6033
rect 8516 5961 8522 5995
rect 8556 5961 8562 5995
rect 8516 5923 8562 5961
rect 8516 5889 8522 5923
rect 8556 5889 8562 5923
rect 8516 5851 8562 5889
rect 8516 5817 8522 5851
rect 8556 5817 8562 5851
rect 8516 5779 8562 5817
rect 8516 5745 8522 5779
rect 8556 5745 8562 5779
rect 8516 5707 8562 5745
rect 8516 5673 8522 5707
rect 8556 5673 8562 5707
rect 8516 5635 8562 5673
rect 8516 5601 8522 5635
rect 8556 5601 8562 5635
rect 8516 5586 8562 5601
rect 8612 6571 8658 6586
rect 8612 6537 8618 6571
rect 8652 6537 8658 6571
rect 8612 6499 8658 6537
rect 8612 6465 8618 6499
rect 8652 6465 8658 6499
rect 8612 6427 8658 6465
rect 8612 6393 8618 6427
rect 8652 6393 8658 6427
rect 8612 6355 8658 6393
rect 8612 6321 8618 6355
rect 8652 6321 8658 6355
rect 8612 6283 8658 6321
rect 8612 6249 8618 6283
rect 8652 6249 8658 6283
rect 8612 6211 8658 6249
rect 8612 6177 8618 6211
rect 8652 6177 8658 6211
rect 8612 6139 8658 6177
rect 8612 6105 8618 6139
rect 8652 6105 8658 6139
rect 8612 6067 8658 6105
rect 8612 6033 8618 6067
rect 8652 6033 8658 6067
rect 8612 5995 8658 6033
rect 8612 5961 8618 5995
rect 8652 5961 8658 5995
rect 8612 5923 8658 5961
rect 8612 5889 8618 5923
rect 8652 5889 8658 5923
rect 8612 5851 8658 5889
rect 8612 5817 8618 5851
rect 8652 5817 8658 5851
rect 8612 5779 8658 5817
rect 8612 5745 8618 5779
rect 8652 5745 8658 5779
rect 8612 5707 8658 5745
rect 8612 5673 8618 5707
rect 8652 5673 8658 5707
rect 8612 5635 8658 5673
rect 8612 5601 8618 5635
rect 8652 5601 8658 5635
rect 8612 5586 8658 5601
rect 8708 6571 8754 6586
rect 8708 6537 8714 6571
rect 8748 6537 8754 6571
rect 8708 6499 8754 6537
rect 8708 6465 8714 6499
rect 8748 6465 8754 6499
rect 8708 6427 8754 6465
rect 8708 6393 8714 6427
rect 8748 6393 8754 6427
rect 8708 6355 8754 6393
rect 8708 6321 8714 6355
rect 8748 6321 8754 6355
rect 8708 6283 8754 6321
rect 8708 6249 8714 6283
rect 8748 6249 8754 6283
rect 8708 6211 8754 6249
rect 8708 6177 8714 6211
rect 8748 6177 8754 6211
rect 8708 6139 8754 6177
rect 8708 6105 8714 6139
rect 8748 6105 8754 6139
rect 8708 6067 8754 6105
rect 8708 6033 8714 6067
rect 8748 6033 8754 6067
rect 8708 5995 8754 6033
rect 8708 5961 8714 5995
rect 8748 5961 8754 5995
rect 8708 5923 8754 5961
rect 8708 5889 8714 5923
rect 8748 5889 8754 5923
rect 8708 5851 8754 5889
rect 8708 5817 8714 5851
rect 8748 5817 8754 5851
rect 8708 5779 8754 5817
rect 8708 5745 8714 5779
rect 8748 5745 8754 5779
rect 8708 5707 8754 5745
rect 8708 5673 8714 5707
rect 8748 5673 8754 5707
rect 8708 5635 8754 5673
rect 8708 5601 8714 5635
rect 8748 5601 8754 5635
rect 8708 5586 8754 5601
rect 9262 6573 9308 6588
rect 9262 6539 9268 6573
rect 9302 6539 9308 6573
rect 9262 6501 9308 6539
rect 9262 6467 9268 6501
rect 9302 6467 9308 6501
rect 9262 6429 9308 6467
rect 9262 6395 9268 6429
rect 9302 6395 9308 6429
rect 9262 6357 9308 6395
rect 9262 6323 9268 6357
rect 9302 6323 9308 6357
rect 9262 6285 9308 6323
rect 9262 6251 9268 6285
rect 9302 6251 9308 6285
rect 9262 6213 9308 6251
rect 9262 6179 9268 6213
rect 9302 6179 9308 6213
rect 9262 6141 9308 6179
rect 9262 6107 9268 6141
rect 9302 6107 9308 6141
rect 9262 6069 9308 6107
rect 9262 6035 9268 6069
rect 9302 6035 9308 6069
rect 9262 5997 9308 6035
rect 9262 5963 9268 5997
rect 9302 5963 9308 5997
rect 9262 5925 9308 5963
rect 9262 5891 9268 5925
rect 9302 5891 9308 5925
rect 9262 5853 9308 5891
rect 9262 5819 9268 5853
rect 9302 5819 9308 5853
rect 9262 5781 9308 5819
rect 9262 5747 9268 5781
rect 9302 5747 9308 5781
rect 9262 5709 9308 5747
rect 9262 5675 9268 5709
rect 9302 5675 9308 5709
rect 9262 5637 9308 5675
rect 9262 5603 9268 5637
rect 9302 5603 9308 5637
rect 9262 5588 9308 5603
rect 9358 6573 9404 6588
rect 9358 6539 9364 6573
rect 9398 6539 9404 6573
rect 9358 6501 9404 6539
rect 9358 6467 9364 6501
rect 9398 6467 9404 6501
rect 9358 6429 9404 6467
rect 9358 6395 9364 6429
rect 9398 6395 9404 6429
rect 9358 6357 9404 6395
rect 9358 6323 9364 6357
rect 9398 6323 9404 6357
rect 9358 6285 9404 6323
rect 9358 6251 9364 6285
rect 9398 6251 9404 6285
rect 9358 6213 9404 6251
rect 9358 6179 9364 6213
rect 9398 6179 9404 6213
rect 9358 6141 9404 6179
rect 9358 6107 9364 6141
rect 9398 6107 9404 6141
rect 9358 6069 9404 6107
rect 9358 6035 9364 6069
rect 9398 6035 9404 6069
rect 9358 5997 9404 6035
rect 9358 5963 9364 5997
rect 9398 5963 9404 5997
rect 9358 5925 9404 5963
rect 9358 5891 9364 5925
rect 9398 5891 9404 5925
rect 9358 5853 9404 5891
rect 9358 5819 9364 5853
rect 9398 5819 9404 5853
rect 9358 5781 9404 5819
rect 9358 5747 9364 5781
rect 9398 5747 9404 5781
rect 9358 5709 9404 5747
rect 9358 5675 9364 5709
rect 9398 5675 9404 5709
rect 9358 5637 9404 5675
rect 9358 5603 9364 5637
rect 9398 5603 9404 5637
rect 9358 5588 9404 5603
rect 9454 6573 9500 6588
rect 9454 6539 9460 6573
rect 9494 6539 9500 6573
rect 9454 6501 9500 6539
rect 9454 6467 9460 6501
rect 9494 6467 9500 6501
rect 9454 6429 9500 6467
rect 9454 6395 9460 6429
rect 9494 6395 9500 6429
rect 9454 6357 9500 6395
rect 9454 6323 9460 6357
rect 9494 6323 9500 6357
rect 9454 6285 9500 6323
rect 9454 6251 9460 6285
rect 9494 6251 9500 6285
rect 9454 6213 9500 6251
rect 9454 6179 9460 6213
rect 9494 6179 9500 6213
rect 9454 6141 9500 6179
rect 9454 6107 9460 6141
rect 9494 6107 9500 6141
rect 9454 6069 9500 6107
rect 9454 6035 9460 6069
rect 9494 6035 9500 6069
rect 9454 5997 9500 6035
rect 9454 5963 9460 5997
rect 9494 5963 9500 5997
rect 9454 5925 9500 5963
rect 9454 5891 9460 5925
rect 9494 5891 9500 5925
rect 9454 5853 9500 5891
rect 9454 5819 9460 5853
rect 9494 5819 9500 5853
rect 9454 5781 9500 5819
rect 9454 5747 9460 5781
rect 9494 5747 9500 5781
rect 9454 5709 9500 5747
rect 9454 5675 9460 5709
rect 9494 5675 9500 5709
rect 9454 5637 9500 5675
rect 9454 5603 9460 5637
rect 9494 5603 9500 5637
rect 9454 5588 9500 5603
rect 9550 6573 9596 6588
rect 9550 6539 9556 6573
rect 9590 6539 9596 6573
rect 9550 6501 9596 6539
rect 9550 6467 9556 6501
rect 9590 6467 9596 6501
rect 9550 6429 9596 6467
rect 9550 6395 9556 6429
rect 9590 6395 9596 6429
rect 9550 6357 9596 6395
rect 9550 6323 9556 6357
rect 9590 6323 9596 6357
rect 9550 6285 9596 6323
rect 9550 6251 9556 6285
rect 9590 6251 9596 6285
rect 9550 6213 9596 6251
rect 9550 6179 9556 6213
rect 9590 6179 9596 6213
rect 9550 6141 9596 6179
rect 9550 6107 9556 6141
rect 9590 6107 9596 6141
rect 9550 6069 9596 6107
rect 9550 6035 9556 6069
rect 9590 6035 9596 6069
rect 9550 5997 9596 6035
rect 9550 5963 9556 5997
rect 9590 5963 9596 5997
rect 9550 5925 9596 5963
rect 9550 5891 9556 5925
rect 9590 5891 9596 5925
rect 9550 5853 9596 5891
rect 9550 5819 9556 5853
rect 9590 5819 9596 5853
rect 9550 5781 9596 5819
rect 9550 5747 9556 5781
rect 9590 5747 9596 5781
rect 9550 5709 9596 5747
rect 9550 5675 9556 5709
rect 9590 5675 9596 5709
rect 9550 5637 9596 5675
rect 9550 5603 9556 5637
rect 9590 5603 9596 5637
rect 9550 5588 9596 5603
rect 9646 6573 9692 6588
rect 9646 6539 9652 6573
rect 9686 6539 9692 6573
rect 9646 6501 9692 6539
rect 9646 6467 9652 6501
rect 9686 6467 9692 6501
rect 9646 6429 9692 6467
rect 9646 6395 9652 6429
rect 9686 6395 9692 6429
rect 9646 6357 9692 6395
rect 9646 6323 9652 6357
rect 9686 6323 9692 6357
rect 9646 6285 9692 6323
rect 9646 6251 9652 6285
rect 9686 6251 9692 6285
rect 9646 6213 9692 6251
rect 9646 6179 9652 6213
rect 9686 6179 9692 6213
rect 9646 6141 9692 6179
rect 9646 6107 9652 6141
rect 9686 6107 9692 6141
rect 9646 6069 9692 6107
rect 9646 6035 9652 6069
rect 9686 6035 9692 6069
rect 9646 5997 9692 6035
rect 9646 5963 9652 5997
rect 9686 5963 9692 5997
rect 9646 5925 9692 5963
rect 9646 5891 9652 5925
rect 9686 5891 9692 5925
rect 9646 5853 9692 5891
rect 9646 5819 9652 5853
rect 9686 5819 9692 5853
rect 9646 5781 9692 5819
rect 9646 5747 9652 5781
rect 9686 5747 9692 5781
rect 9646 5709 9692 5747
rect 9646 5675 9652 5709
rect 9686 5675 9692 5709
rect 9646 5637 9692 5675
rect 9646 5603 9652 5637
rect 9686 5603 9692 5637
rect 9646 5588 9692 5603
rect 9742 6573 9788 6588
rect 9742 6539 9748 6573
rect 9782 6539 9788 6573
rect 9742 6501 9788 6539
rect 9742 6467 9748 6501
rect 9782 6467 9788 6501
rect 9742 6429 9788 6467
rect 9742 6395 9748 6429
rect 9782 6395 9788 6429
rect 9742 6357 9788 6395
rect 9742 6323 9748 6357
rect 9782 6323 9788 6357
rect 9742 6285 9788 6323
rect 9742 6251 9748 6285
rect 9782 6251 9788 6285
rect 9742 6213 9788 6251
rect 9742 6179 9748 6213
rect 9782 6179 9788 6213
rect 9742 6141 9788 6179
rect 9742 6107 9748 6141
rect 9782 6107 9788 6141
rect 9742 6069 9788 6107
rect 9742 6035 9748 6069
rect 9782 6035 9788 6069
rect 9742 5997 9788 6035
rect 9742 5963 9748 5997
rect 9782 5963 9788 5997
rect 9742 5925 9788 5963
rect 9742 5891 9748 5925
rect 9782 5891 9788 5925
rect 9742 5853 9788 5891
rect 9742 5819 9748 5853
rect 9782 5819 9788 5853
rect 9742 5781 9788 5819
rect 9742 5747 9748 5781
rect 9782 5747 9788 5781
rect 9742 5709 9788 5747
rect 9742 5675 9748 5709
rect 9782 5675 9788 5709
rect 9742 5637 9788 5675
rect 9742 5603 9748 5637
rect 9782 5603 9788 5637
rect 9742 5588 9788 5603
rect 9838 6573 9884 6588
rect 9838 6539 9844 6573
rect 9878 6539 9884 6573
rect 9838 6501 9884 6539
rect 9838 6467 9844 6501
rect 9878 6467 9884 6501
rect 9838 6429 9884 6467
rect 9838 6395 9844 6429
rect 9878 6395 9884 6429
rect 9838 6357 9884 6395
rect 9838 6323 9844 6357
rect 9878 6323 9884 6357
rect 9838 6285 9884 6323
rect 9838 6251 9844 6285
rect 9878 6251 9884 6285
rect 9838 6213 9884 6251
rect 9838 6179 9844 6213
rect 9878 6179 9884 6213
rect 9838 6141 9884 6179
rect 9838 6107 9844 6141
rect 9878 6107 9884 6141
rect 9838 6069 9884 6107
rect 9838 6035 9844 6069
rect 9878 6035 9884 6069
rect 9838 5997 9884 6035
rect 9838 5963 9844 5997
rect 9878 5963 9884 5997
rect 9838 5925 9884 5963
rect 9838 5891 9844 5925
rect 9878 5891 9884 5925
rect 9838 5853 9884 5891
rect 9838 5819 9844 5853
rect 9878 5819 9884 5853
rect 9838 5781 9884 5819
rect 9838 5747 9844 5781
rect 9878 5747 9884 5781
rect 9838 5709 9884 5747
rect 9838 5675 9844 5709
rect 9878 5675 9884 5709
rect 9838 5637 9884 5675
rect 9838 5603 9844 5637
rect 9878 5603 9884 5637
rect 9838 5588 9884 5603
rect 9934 6573 9980 6588
rect 9934 6539 9940 6573
rect 9974 6539 9980 6573
rect 9934 6501 9980 6539
rect 9934 6467 9940 6501
rect 9974 6467 9980 6501
rect 9934 6429 9980 6467
rect 9934 6395 9940 6429
rect 9974 6395 9980 6429
rect 9934 6357 9980 6395
rect 9934 6323 9940 6357
rect 9974 6323 9980 6357
rect 9934 6285 9980 6323
rect 9934 6251 9940 6285
rect 9974 6251 9980 6285
rect 9934 6213 9980 6251
rect 9934 6179 9940 6213
rect 9974 6179 9980 6213
rect 9934 6141 9980 6179
rect 9934 6107 9940 6141
rect 9974 6107 9980 6141
rect 9934 6069 9980 6107
rect 9934 6035 9940 6069
rect 9974 6035 9980 6069
rect 9934 5997 9980 6035
rect 9934 5963 9940 5997
rect 9974 5963 9980 5997
rect 9934 5925 9980 5963
rect 9934 5891 9940 5925
rect 9974 5891 9980 5925
rect 9934 5853 9980 5891
rect 9934 5819 9940 5853
rect 9974 5819 9980 5853
rect 9934 5781 9980 5819
rect 9934 5747 9940 5781
rect 9974 5747 9980 5781
rect 9934 5709 9980 5747
rect 9934 5675 9940 5709
rect 9974 5675 9980 5709
rect 9934 5637 9980 5675
rect 9934 5603 9940 5637
rect 9974 5603 9980 5637
rect 9934 5588 9980 5603
rect 10030 6573 10076 6588
rect 10030 6539 10036 6573
rect 10070 6539 10076 6573
rect 10030 6501 10076 6539
rect 10030 6467 10036 6501
rect 10070 6467 10076 6501
rect 10030 6429 10076 6467
rect 10030 6395 10036 6429
rect 10070 6395 10076 6429
rect 10030 6357 10076 6395
rect 10030 6323 10036 6357
rect 10070 6323 10076 6357
rect 10030 6285 10076 6323
rect 10030 6251 10036 6285
rect 10070 6251 10076 6285
rect 10030 6213 10076 6251
rect 10030 6179 10036 6213
rect 10070 6179 10076 6213
rect 10030 6141 10076 6179
rect 10030 6107 10036 6141
rect 10070 6107 10076 6141
rect 10030 6069 10076 6107
rect 10030 6035 10036 6069
rect 10070 6035 10076 6069
rect 10030 5997 10076 6035
rect 10030 5963 10036 5997
rect 10070 5963 10076 5997
rect 10030 5925 10076 5963
rect 10030 5891 10036 5925
rect 10070 5891 10076 5925
rect 10030 5853 10076 5891
rect 10030 5819 10036 5853
rect 10070 5819 10076 5853
rect 10030 5781 10076 5819
rect 10030 5747 10036 5781
rect 10070 5747 10076 5781
rect 10030 5709 10076 5747
rect 10030 5675 10036 5709
rect 10070 5675 10076 5709
rect 10030 5637 10076 5675
rect 10030 5603 10036 5637
rect 10070 5603 10076 5637
rect 10030 5588 10076 5603
rect 10126 6573 10172 6588
rect 10126 6539 10132 6573
rect 10166 6539 10172 6573
rect 10126 6501 10172 6539
rect 10126 6467 10132 6501
rect 10166 6467 10172 6501
rect 10126 6429 10172 6467
rect 10126 6395 10132 6429
rect 10166 6395 10172 6429
rect 10126 6357 10172 6395
rect 10126 6323 10132 6357
rect 10166 6323 10172 6357
rect 10126 6285 10172 6323
rect 10126 6251 10132 6285
rect 10166 6251 10172 6285
rect 10126 6213 10172 6251
rect 10126 6179 10132 6213
rect 10166 6179 10172 6213
rect 10126 6141 10172 6179
rect 10126 6107 10132 6141
rect 10166 6107 10172 6141
rect 10126 6069 10172 6107
rect 10126 6035 10132 6069
rect 10166 6035 10172 6069
rect 10126 5997 10172 6035
rect 10126 5963 10132 5997
rect 10166 5963 10172 5997
rect 10126 5925 10172 5963
rect 10126 5891 10132 5925
rect 10166 5891 10172 5925
rect 10126 5853 10172 5891
rect 10126 5819 10132 5853
rect 10166 5819 10172 5853
rect 10126 5781 10172 5819
rect 10126 5747 10132 5781
rect 10166 5747 10172 5781
rect 10126 5709 10172 5747
rect 10126 5675 10132 5709
rect 10166 5675 10172 5709
rect 10126 5637 10172 5675
rect 10126 5603 10132 5637
rect 10166 5603 10172 5637
rect 10126 5588 10172 5603
rect 10222 6573 10268 6588
rect 10222 6539 10228 6573
rect 10262 6539 10268 6573
rect 10222 6501 10268 6539
rect 10222 6467 10228 6501
rect 10262 6467 10268 6501
rect 10222 6429 10268 6467
rect 10222 6395 10228 6429
rect 10262 6395 10268 6429
rect 10222 6357 10268 6395
rect 10222 6323 10228 6357
rect 10262 6323 10268 6357
rect 10222 6285 10268 6323
rect 10222 6251 10228 6285
rect 10262 6251 10268 6285
rect 10222 6213 10268 6251
rect 10222 6179 10228 6213
rect 10262 6179 10268 6213
rect 10222 6141 10268 6179
rect 10222 6107 10228 6141
rect 10262 6107 10268 6141
rect 10222 6069 10268 6107
rect 10222 6035 10228 6069
rect 10262 6035 10268 6069
rect 10222 5997 10268 6035
rect 10222 5963 10228 5997
rect 10262 5963 10268 5997
rect 10222 5925 10268 5963
rect 10222 5891 10228 5925
rect 10262 5891 10268 5925
rect 10222 5853 10268 5891
rect 10222 5819 10228 5853
rect 10262 5819 10268 5853
rect 10222 5781 10268 5819
rect 10222 5747 10228 5781
rect 10262 5747 10268 5781
rect 10222 5709 10268 5747
rect 10222 5675 10228 5709
rect 10262 5675 10268 5709
rect 10222 5637 10268 5675
rect 10222 5603 10228 5637
rect 10262 5603 10268 5637
rect 10222 5588 10268 5603
rect 10318 6573 10364 6588
rect 10318 6539 10324 6573
rect 10358 6539 10364 6573
rect 10318 6501 10364 6539
rect 10318 6467 10324 6501
rect 10358 6467 10364 6501
rect 10318 6429 10364 6467
rect 10318 6395 10324 6429
rect 10358 6395 10364 6429
rect 10318 6357 10364 6395
rect 10318 6323 10324 6357
rect 10358 6323 10364 6357
rect 10318 6285 10364 6323
rect 10318 6251 10324 6285
rect 10358 6251 10364 6285
rect 10318 6213 10364 6251
rect 10318 6179 10324 6213
rect 10358 6179 10364 6213
rect 10318 6141 10364 6179
rect 10318 6107 10324 6141
rect 10358 6107 10364 6141
rect 10318 6069 10364 6107
rect 10318 6035 10324 6069
rect 10358 6035 10364 6069
rect 10318 5997 10364 6035
rect 10318 5963 10324 5997
rect 10358 5963 10364 5997
rect 10318 5925 10364 5963
rect 10318 5891 10324 5925
rect 10358 5891 10364 5925
rect 10318 5853 10364 5891
rect 10318 5819 10324 5853
rect 10358 5819 10364 5853
rect 10318 5781 10364 5819
rect 10318 5747 10324 5781
rect 10358 5747 10364 5781
rect 10318 5709 10364 5747
rect 10318 5675 10324 5709
rect 10358 5675 10364 5709
rect 10318 5637 10364 5675
rect 10318 5603 10324 5637
rect 10358 5603 10364 5637
rect 10318 5588 10364 5603
rect 10414 6573 10460 6588
rect 10414 6539 10420 6573
rect 10454 6539 10460 6573
rect 10414 6501 10460 6539
rect 10414 6467 10420 6501
rect 10454 6467 10460 6501
rect 10414 6429 10460 6467
rect 10414 6395 10420 6429
rect 10454 6395 10460 6429
rect 10414 6357 10460 6395
rect 10414 6323 10420 6357
rect 10454 6323 10460 6357
rect 10414 6285 10460 6323
rect 10414 6251 10420 6285
rect 10454 6251 10460 6285
rect 10414 6213 10460 6251
rect 10414 6179 10420 6213
rect 10454 6179 10460 6213
rect 10414 6141 10460 6179
rect 10414 6107 10420 6141
rect 10454 6107 10460 6141
rect 10414 6069 10460 6107
rect 10414 6035 10420 6069
rect 10454 6035 10460 6069
rect 10414 5997 10460 6035
rect 10414 5963 10420 5997
rect 10454 5963 10460 5997
rect 10414 5925 10460 5963
rect 10414 5891 10420 5925
rect 10454 5891 10460 5925
rect 10414 5853 10460 5891
rect 10414 5819 10420 5853
rect 10454 5819 10460 5853
rect 10414 5781 10460 5819
rect 10414 5747 10420 5781
rect 10454 5747 10460 5781
rect 10414 5709 10460 5747
rect 10414 5675 10420 5709
rect 10454 5675 10460 5709
rect 10414 5637 10460 5675
rect 10414 5603 10420 5637
rect 10454 5603 10460 5637
rect 10414 5588 10460 5603
rect 11028 6569 11074 6584
rect 11028 6535 11034 6569
rect 11068 6535 11074 6569
rect 11028 6497 11074 6535
rect 11028 6463 11034 6497
rect 11068 6463 11074 6497
rect 11028 6425 11074 6463
rect 11028 6391 11034 6425
rect 11068 6391 11074 6425
rect 11028 6353 11074 6391
rect 11028 6319 11034 6353
rect 11068 6319 11074 6353
rect 11028 6281 11074 6319
rect 11028 6247 11034 6281
rect 11068 6247 11074 6281
rect 11028 6209 11074 6247
rect 11028 6175 11034 6209
rect 11068 6175 11074 6209
rect 11028 6137 11074 6175
rect 11028 6103 11034 6137
rect 11068 6103 11074 6137
rect 11028 6065 11074 6103
rect 11028 6031 11034 6065
rect 11068 6031 11074 6065
rect 11028 5993 11074 6031
rect 11028 5959 11034 5993
rect 11068 5959 11074 5993
rect 11028 5921 11074 5959
rect 11028 5887 11034 5921
rect 11068 5887 11074 5921
rect 11028 5849 11074 5887
rect 11028 5815 11034 5849
rect 11068 5815 11074 5849
rect 11028 5777 11074 5815
rect 11028 5743 11034 5777
rect 11068 5743 11074 5777
rect 11028 5705 11074 5743
rect 11028 5671 11034 5705
rect 11068 5671 11074 5705
rect 11028 5633 11074 5671
rect 11028 5599 11034 5633
rect 11068 5599 11074 5633
rect 11028 5584 11074 5599
rect 11124 6569 11170 6584
rect 11124 6535 11130 6569
rect 11164 6535 11170 6569
rect 11124 6497 11170 6535
rect 11124 6463 11130 6497
rect 11164 6463 11170 6497
rect 11124 6425 11170 6463
rect 11124 6391 11130 6425
rect 11164 6391 11170 6425
rect 11124 6353 11170 6391
rect 11124 6319 11130 6353
rect 11164 6319 11170 6353
rect 11124 6281 11170 6319
rect 11124 6247 11130 6281
rect 11164 6247 11170 6281
rect 11124 6209 11170 6247
rect 11124 6175 11130 6209
rect 11164 6175 11170 6209
rect 11124 6137 11170 6175
rect 11124 6103 11130 6137
rect 11164 6103 11170 6137
rect 11124 6065 11170 6103
rect 11124 6031 11130 6065
rect 11164 6031 11170 6065
rect 11124 5993 11170 6031
rect 11124 5959 11130 5993
rect 11164 5959 11170 5993
rect 11124 5921 11170 5959
rect 11124 5887 11130 5921
rect 11164 5887 11170 5921
rect 11124 5849 11170 5887
rect 11124 5815 11130 5849
rect 11164 5815 11170 5849
rect 11124 5777 11170 5815
rect 11124 5743 11130 5777
rect 11164 5743 11170 5777
rect 11124 5705 11170 5743
rect 11124 5671 11130 5705
rect 11164 5671 11170 5705
rect 11124 5633 11170 5671
rect 11124 5599 11130 5633
rect 11164 5599 11170 5633
rect 11124 5584 11170 5599
rect 11220 6569 11266 6584
rect 11220 6535 11226 6569
rect 11260 6535 11266 6569
rect 11220 6497 11266 6535
rect 11220 6463 11226 6497
rect 11260 6463 11266 6497
rect 11220 6425 11266 6463
rect 11220 6391 11226 6425
rect 11260 6391 11266 6425
rect 11220 6353 11266 6391
rect 11220 6319 11226 6353
rect 11260 6319 11266 6353
rect 11220 6281 11266 6319
rect 11220 6247 11226 6281
rect 11260 6247 11266 6281
rect 11220 6209 11266 6247
rect 11220 6175 11226 6209
rect 11260 6175 11266 6209
rect 11220 6137 11266 6175
rect 11220 6103 11226 6137
rect 11260 6103 11266 6137
rect 11220 6065 11266 6103
rect 11220 6031 11226 6065
rect 11260 6031 11266 6065
rect 11220 5993 11266 6031
rect 11220 5959 11226 5993
rect 11260 5959 11266 5993
rect 11220 5921 11266 5959
rect 11220 5887 11226 5921
rect 11260 5887 11266 5921
rect 11220 5849 11266 5887
rect 11220 5815 11226 5849
rect 11260 5815 11266 5849
rect 11220 5777 11266 5815
rect 11220 5743 11226 5777
rect 11260 5743 11266 5777
rect 11220 5705 11266 5743
rect 11220 5671 11226 5705
rect 11260 5671 11266 5705
rect 11220 5633 11266 5671
rect 11220 5599 11226 5633
rect 11260 5599 11266 5633
rect 11220 5584 11266 5599
rect 11316 6569 11362 6584
rect 11316 6535 11322 6569
rect 11356 6535 11362 6569
rect 11316 6497 11362 6535
rect 11316 6463 11322 6497
rect 11356 6463 11362 6497
rect 11316 6425 11362 6463
rect 11316 6391 11322 6425
rect 11356 6391 11362 6425
rect 11316 6353 11362 6391
rect 11316 6319 11322 6353
rect 11356 6319 11362 6353
rect 11316 6281 11362 6319
rect 11316 6247 11322 6281
rect 11356 6247 11362 6281
rect 11316 6209 11362 6247
rect 11316 6175 11322 6209
rect 11356 6175 11362 6209
rect 11316 6137 11362 6175
rect 11316 6103 11322 6137
rect 11356 6103 11362 6137
rect 11316 6065 11362 6103
rect 11316 6031 11322 6065
rect 11356 6031 11362 6065
rect 11316 5993 11362 6031
rect 11316 5959 11322 5993
rect 11356 5959 11362 5993
rect 11316 5921 11362 5959
rect 11316 5887 11322 5921
rect 11356 5887 11362 5921
rect 11316 5849 11362 5887
rect 11316 5815 11322 5849
rect 11356 5815 11362 5849
rect 11316 5777 11362 5815
rect 11316 5743 11322 5777
rect 11356 5743 11362 5777
rect 11316 5705 11362 5743
rect 11316 5671 11322 5705
rect 11356 5671 11362 5705
rect 11316 5633 11362 5671
rect 11316 5599 11322 5633
rect 11356 5599 11362 5633
rect 11316 5584 11362 5599
rect 11412 6569 11458 6584
rect 11412 6535 11418 6569
rect 11452 6535 11458 6569
rect 11412 6497 11458 6535
rect 11412 6463 11418 6497
rect 11452 6463 11458 6497
rect 11412 6425 11458 6463
rect 11412 6391 11418 6425
rect 11452 6391 11458 6425
rect 11412 6353 11458 6391
rect 11412 6319 11418 6353
rect 11452 6319 11458 6353
rect 11412 6281 11458 6319
rect 11412 6247 11418 6281
rect 11452 6247 11458 6281
rect 11412 6209 11458 6247
rect 11412 6175 11418 6209
rect 11452 6175 11458 6209
rect 11412 6137 11458 6175
rect 11412 6103 11418 6137
rect 11452 6103 11458 6137
rect 11412 6065 11458 6103
rect 11412 6031 11418 6065
rect 11452 6031 11458 6065
rect 11412 5993 11458 6031
rect 11412 5959 11418 5993
rect 11452 5959 11458 5993
rect 11412 5921 11458 5959
rect 11412 5887 11418 5921
rect 11452 5887 11458 5921
rect 11412 5849 11458 5887
rect 11412 5815 11418 5849
rect 11452 5815 11458 5849
rect 11412 5777 11458 5815
rect 11412 5743 11418 5777
rect 11452 5743 11458 5777
rect 11412 5705 11458 5743
rect 11412 5671 11418 5705
rect 11452 5671 11458 5705
rect 11412 5633 11458 5671
rect 11412 5599 11418 5633
rect 11452 5599 11458 5633
rect 11412 5584 11458 5599
rect 11508 6569 11554 6584
rect 11508 6535 11514 6569
rect 11548 6535 11554 6569
rect 11508 6497 11554 6535
rect 11508 6463 11514 6497
rect 11548 6463 11554 6497
rect 11508 6425 11554 6463
rect 11508 6391 11514 6425
rect 11548 6391 11554 6425
rect 11508 6353 11554 6391
rect 11508 6319 11514 6353
rect 11548 6319 11554 6353
rect 11508 6281 11554 6319
rect 11508 6247 11514 6281
rect 11548 6247 11554 6281
rect 11508 6209 11554 6247
rect 11508 6175 11514 6209
rect 11548 6175 11554 6209
rect 11508 6137 11554 6175
rect 11508 6103 11514 6137
rect 11548 6103 11554 6137
rect 11508 6065 11554 6103
rect 11508 6031 11514 6065
rect 11548 6031 11554 6065
rect 11508 5993 11554 6031
rect 11508 5959 11514 5993
rect 11548 5959 11554 5993
rect 11508 5921 11554 5959
rect 11508 5887 11514 5921
rect 11548 5887 11554 5921
rect 11508 5849 11554 5887
rect 11508 5815 11514 5849
rect 11548 5815 11554 5849
rect 11508 5777 11554 5815
rect 11508 5743 11514 5777
rect 11548 5743 11554 5777
rect 11508 5705 11554 5743
rect 11508 5671 11514 5705
rect 11548 5671 11554 5705
rect 11508 5633 11554 5671
rect 11508 5599 11514 5633
rect 11548 5599 11554 5633
rect 11508 5584 11554 5599
rect 11604 6569 11650 6584
rect 11604 6535 11610 6569
rect 11644 6535 11650 6569
rect 11604 6497 11650 6535
rect 11604 6463 11610 6497
rect 11644 6463 11650 6497
rect 11604 6425 11650 6463
rect 11604 6391 11610 6425
rect 11644 6391 11650 6425
rect 11604 6353 11650 6391
rect 11604 6319 11610 6353
rect 11644 6319 11650 6353
rect 11604 6281 11650 6319
rect 11604 6247 11610 6281
rect 11644 6247 11650 6281
rect 11604 6209 11650 6247
rect 11604 6175 11610 6209
rect 11644 6175 11650 6209
rect 11604 6137 11650 6175
rect 11604 6103 11610 6137
rect 11644 6103 11650 6137
rect 11604 6065 11650 6103
rect 11604 6031 11610 6065
rect 11644 6031 11650 6065
rect 11604 5993 11650 6031
rect 11604 5959 11610 5993
rect 11644 5959 11650 5993
rect 11604 5921 11650 5959
rect 11604 5887 11610 5921
rect 11644 5887 11650 5921
rect 11604 5849 11650 5887
rect 11604 5815 11610 5849
rect 11644 5815 11650 5849
rect 11604 5777 11650 5815
rect 11604 5743 11610 5777
rect 11644 5743 11650 5777
rect 11604 5705 11650 5743
rect 11604 5671 11610 5705
rect 11644 5671 11650 5705
rect 11604 5633 11650 5671
rect 11604 5599 11610 5633
rect 11644 5599 11650 5633
rect 11604 5584 11650 5599
rect 11700 6569 11746 6584
rect 11700 6535 11706 6569
rect 11740 6535 11746 6569
rect 11700 6497 11746 6535
rect 11700 6463 11706 6497
rect 11740 6463 11746 6497
rect 11700 6425 11746 6463
rect 11700 6391 11706 6425
rect 11740 6391 11746 6425
rect 11700 6353 11746 6391
rect 11700 6319 11706 6353
rect 11740 6319 11746 6353
rect 11700 6281 11746 6319
rect 11700 6247 11706 6281
rect 11740 6247 11746 6281
rect 11700 6209 11746 6247
rect 11700 6175 11706 6209
rect 11740 6175 11746 6209
rect 11700 6137 11746 6175
rect 11700 6103 11706 6137
rect 11740 6103 11746 6137
rect 11700 6065 11746 6103
rect 11700 6031 11706 6065
rect 11740 6031 11746 6065
rect 11700 5993 11746 6031
rect 11700 5959 11706 5993
rect 11740 5959 11746 5993
rect 11700 5921 11746 5959
rect 11700 5887 11706 5921
rect 11740 5887 11746 5921
rect 11700 5849 11746 5887
rect 11700 5815 11706 5849
rect 11740 5815 11746 5849
rect 11700 5777 11746 5815
rect 11700 5743 11706 5777
rect 11740 5743 11746 5777
rect 11700 5705 11746 5743
rect 11700 5671 11706 5705
rect 11740 5671 11746 5705
rect 11700 5633 11746 5671
rect 11700 5599 11706 5633
rect 11740 5599 11746 5633
rect 11700 5584 11746 5599
rect 11796 6569 11842 6584
rect 11796 6535 11802 6569
rect 11836 6535 11842 6569
rect 11796 6497 11842 6535
rect 11796 6463 11802 6497
rect 11836 6463 11842 6497
rect 11796 6425 11842 6463
rect 11796 6391 11802 6425
rect 11836 6391 11842 6425
rect 11796 6353 11842 6391
rect 11796 6319 11802 6353
rect 11836 6319 11842 6353
rect 11796 6281 11842 6319
rect 11796 6247 11802 6281
rect 11836 6247 11842 6281
rect 11796 6209 11842 6247
rect 11796 6175 11802 6209
rect 11836 6175 11842 6209
rect 11796 6137 11842 6175
rect 11796 6103 11802 6137
rect 11836 6103 11842 6137
rect 11796 6065 11842 6103
rect 11796 6031 11802 6065
rect 11836 6031 11842 6065
rect 11796 5993 11842 6031
rect 11796 5959 11802 5993
rect 11836 5959 11842 5993
rect 11796 5921 11842 5959
rect 11796 5887 11802 5921
rect 11836 5887 11842 5921
rect 11796 5849 11842 5887
rect 11796 5815 11802 5849
rect 11836 5815 11842 5849
rect 11796 5777 11842 5815
rect 11796 5743 11802 5777
rect 11836 5743 11842 5777
rect 11796 5705 11842 5743
rect 11796 5671 11802 5705
rect 11836 5671 11842 5705
rect 11796 5633 11842 5671
rect 11796 5599 11802 5633
rect 11836 5599 11842 5633
rect 11796 5584 11842 5599
rect 12418 6547 12464 6562
rect 12418 6513 12424 6547
rect 12458 6513 12464 6547
rect 12418 6475 12464 6513
rect 12418 6441 12424 6475
rect 12458 6441 12464 6475
rect 12418 6403 12464 6441
rect 12418 6369 12424 6403
rect 12458 6369 12464 6403
rect 12418 6331 12464 6369
rect 12418 6297 12424 6331
rect 12458 6297 12464 6331
rect 12418 6259 12464 6297
rect 12418 6225 12424 6259
rect 12458 6225 12464 6259
rect 12418 6187 12464 6225
rect 12418 6153 12424 6187
rect 12458 6153 12464 6187
rect 12418 6115 12464 6153
rect 12418 6081 12424 6115
rect 12458 6081 12464 6115
rect 12418 6043 12464 6081
rect 12418 6009 12424 6043
rect 12458 6009 12464 6043
rect 12418 5971 12464 6009
rect 12418 5937 12424 5971
rect 12458 5937 12464 5971
rect 12418 5899 12464 5937
rect 12418 5865 12424 5899
rect 12458 5865 12464 5899
rect 12418 5827 12464 5865
rect 12418 5793 12424 5827
rect 12458 5793 12464 5827
rect 12418 5755 12464 5793
rect 12418 5721 12424 5755
rect 12458 5721 12464 5755
rect 12418 5683 12464 5721
rect 12418 5649 12424 5683
rect 12458 5649 12464 5683
rect 12418 5611 12464 5649
rect 12418 5577 12424 5611
rect 12458 5577 12464 5611
rect 12418 5562 12464 5577
rect 12514 6547 12560 6562
rect 12514 6513 12520 6547
rect 12554 6513 12560 6547
rect 12514 6475 12560 6513
rect 12514 6441 12520 6475
rect 12554 6441 12560 6475
rect 12514 6403 12560 6441
rect 12514 6369 12520 6403
rect 12554 6369 12560 6403
rect 12514 6331 12560 6369
rect 12514 6297 12520 6331
rect 12554 6297 12560 6331
rect 12514 6259 12560 6297
rect 12514 6225 12520 6259
rect 12554 6225 12560 6259
rect 12514 6187 12560 6225
rect 12514 6153 12520 6187
rect 12554 6153 12560 6187
rect 12514 6115 12560 6153
rect 12514 6081 12520 6115
rect 12554 6081 12560 6115
rect 12514 6043 12560 6081
rect 12514 6009 12520 6043
rect 12554 6009 12560 6043
rect 12514 5971 12560 6009
rect 12514 5937 12520 5971
rect 12554 5937 12560 5971
rect 12514 5899 12560 5937
rect 12514 5865 12520 5899
rect 12554 5865 12560 5899
rect 12514 5827 12560 5865
rect 12514 5793 12520 5827
rect 12554 5793 12560 5827
rect 12514 5755 12560 5793
rect 12514 5721 12520 5755
rect 12554 5721 12560 5755
rect 12514 5683 12560 5721
rect 12514 5649 12520 5683
rect 12554 5649 12560 5683
rect 12514 5611 12560 5649
rect 12514 5577 12520 5611
rect 12554 5577 12560 5611
rect 12514 5562 12560 5577
rect 12610 6547 12656 6562
rect 12610 6513 12616 6547
rect 12650 6513 12656 6547
rect 12610 6475 12656 6513
rect 12610 6441 12616 6475
rect 12650 6441 12656 6475
rect 12610 6403 12656 6441
rect 12610 6369 12616 6403
rect 12650 6369 12656 6403
rect 12610 6331 12656 6369
rect 12610 6297 12616 6331
rect 12650 6297 12656 6331
rect 12610 6259 12656 6297
rect 12610 6225 12616 6259
rect 12650 6225 12656 6259
rect 12610 6187 12656 6225
rect 12610 6153 12616 6187
rect 12650 6153 12656 6187
rect 12610 6115 12656 6153
rect 12610 6081 12616 6115
rect 12650 6081 12656 6115
rect 12610 6043 12656 6081
rect 12610 6009 12616 6043
rect 12650 6009 12656 6043
rect 12610 5971 12656 6009
rect 12610 5937 12616 5971
rect 12650 5937 12656 5971
rect 12610 5899 12656 5937
rect 12610 5865 12616 5899
rect 12650 5865 12656 5899
rect 12610 5827 12656 5865
rect 12610 5793 12616 5827
rect 12650 5793 12656 5827
rect 12610 5755 12656 5793
rect 12610 5721 12616 5755
rect 12650 5721 12656 5755
rect 12610 5683 12656 5721
rect 12610 5649 12616 5683
rect 12650 5649 12656 5683
rect 12610 5611 12656 5649
rect 12610 5577 12616 5611
rect 12650 5577 12656 5611
rect 12610 5562 12656 5577
rect 12706 6547 12752 6562
rect 12706 6513 12712 6547
rect 12746 6513 12752 6547
rect 12706 6475 12752 6513
rect 12706 6441 12712 6475
rect 12746 6441 12752 6475
rect 12706 6403 12752 6441
rect 12706 6369 12712 6403
rect 12746 6369 12752 6403
rect 12706 6331 12752 6369
rect 12706 6297 12712 6331
rect 12746 6297 12752 6331
rect 12706 6259 12752 6297
rect 12706 6225 12712 6259
rect 12746 6225 12752 6259
rect 12706 6187 12752 6225
rect 12706 6153 12712 6187
rect 12746 6153 12752 6187
rect 12706 6115 12752 6153
rect 12706 6081 12712 6115
rect 12746 6081 12752 6115
rect 12706 6043 12752 6081
rect 12706 6009 12712 6043
rect 12746 6009 12752 6043
rect 12706 5971 12752 6009
rect 12706 5937 12712 5971
rect 12746 5937 12752 5971
rect 12706 5899 12752 5937
rect 12706 5865 12712 5899
rect 12746 5865 12752 5899
rect 12706 5827 12752 5865
rect 12706 5793 12712 5827
rect 12746 5793 12752 5827
rect 12706 5755 12752 5793
rect 12706 5721 12712 5755
rect 12746 5721 12752 5755
rect 12706 5683 12752 5721
rect 12706 5649 12712 5683
rect 12746 5649 12752 5683
rect 12706 5611 12752 5649
rect 12706 5577 12712 5611
rect 12746 5577 12752 5611
rect 12706 5562 12752 5577
rect 12802 6547 12848 6562
rect 12802 6513 12808 6547
rect 12842 6513 12848 6547
rect 12802 6475 12848 6513
rect 12802 6441 12808 6475
rect 12842 6441 12848 6475
rect 12802 6403 12848 6441
rect 12802 6369 12808 6403
rect 12842 6369 12848 6403
rect 12802 6331 12848 6369
rect 12802 6297 12808 6331
rect 12842 6297 12848 6331
rect 12802 6259 12848 6297
rect 12802 6225 12808 6259
rect 12842 6225 12848 6259
rect 12802 6187 12848 6225
rect 12802 6153 12808 6187
rect 12842 6153 12848 6187
rect 12802 6115 12848 6153
rect 12802 6081 12808 6115
rect 12842 6081 12848 6115
rect 12802 6043 12848 6081
rect 12802 6009 12808 6043
rect 12842 6009 12848 6043
rect 12802 5971 12848 6009
rect 12802 5937 12808 5971
rect 12842 5937 12848 5971
rect 12802 5899 12848 5937
rect 12802 5865 12808 5899
rect 12842 5865 12848 5899
rect 12802 5827 12848 5865
rect 12802 5793 12808 5827
rect 12842 5793 12848 5827
rect 12802 5755 12848 5793
rect 12802 5721 12808 5755
rect 12842 5721 12848 5755
rect 12802 5683 12848 5721
rect 12802 5649 12808 5683
rect 12842 5649 12848 5683
rect 12802 5611 12848 5649
rect 12802 5577 12808 5611
rect 12842 5577 12848 5611
rect 12802 5562 12848 5577
rect 12898 6547 12944 6562
rect 12898 6513 12904 6547
rect 12938 6513 12944 6547
rect 12898 6475 12944 6513
rect 12898 6441 12904 6475
rect 12938 6441 12944 6475
rect 12898 6403 12944 6441
rect 12898 6369 12904 6403
rect 12938 6369 12944 6403
rect 12898 6331 12944 6369
rect 12898 6297 12904 6331
rect 12938 6297 12944 6331
rect 12898 6259 12944 6297
rect 12898 6225 12904 6259
rect 12938 6225 12944 6259
rect 12898 6187 12944 6225
rect 12898 6153 12904 6187
rect 12938 6153 12944 6187
rect 12898 6115 12944 6153
rect 12898 6081 12904 6115
rect 12938 6081 12944 6115
rect 12898 6043 12944 6081
rect 12898 6009 12904 6043
rect 12938 6009 12944 6043
rect 12898 5971 12944 6009
rect 12898 5937 12904 5971
rect 12938 5937 12944 5971
rect 12898 5899 12944 5937
rect 12898 5865 12904 5899
rect 12938 5865 12944 5899
rect 12898 5827 12944 5865
rect 12898 5793 12904 5827
rect 12938 5793 12944 5827
rect 12898 5755 12944 5793
rect 12898 5721 12904 5755
rect 12938 5721 12944 5755
rect 12898 5683 12944 5721
rect 12898 5649 12904 5683
rect 12938 5649 12944 5683
rect 12898 5611 12944 5649
rect 12898 5577 12904 5611
rect 12938 5577 12944 5611
rect 12898 5562 12944 5577
rect 12994 6547 13040 6562
rect 12994 6513 13000 6547
rect 13034 6513 13040 6547
rect 12994 6475 13040 6513
rect 12994 6441 13000 6475
rect 13034 6441 13040 6475
rect 12994 6403 13040 6441
rect 12994 6369 13000 6403
rect 13034 6369 13040 6403
rect 12994 6331 13040 6369
rect 12994 6297 13000 6331
rect 13034 6297 13040 6331
rect 12994 6259 13040 6297
rect 12994 6225 13000 6259
rect 13034 6225 13040 6259
rect 12994 6187 13040 6225
rect 12994 6153 13000 6187
rect 13034 6153 13040 6187
rect 12994 6115 13040 6153
rect 12994 6081 13000 6115
rect 13034 6081 13040 6115
rect 12994 6043 13040 6081
rect 12994 6009 13000 6043
rect 13034 6009 13040 6043
rect 12994 5971 13040 6009
rect 12994 5937 13000 5971
rect 13034 5937 13040 5971
rect 12994 5899 13040 5937
rect 12994 5865 13000 5899
rect 13034 5865 13040 5899
rect 12994 5827 13040 5865
rect 12994 5793 13000 5827
rect 13034 5793 13040 5827
rect 12994 5755 13040 5793
rect 12994 5721 13000 5755
rect 13034 5721 13040 5755
rect 12994 5683 13040 5721
rect 12994 5649 13000 5683
rect 13034 5649 13040 5683
rect 12994 5611 13040 5649
rect 12994 5577 13000 5611
rect 13034 5577 13040 5611
rect 12994 5562 13040 5577
rect 13090 6547 13136 6562
rect 13090 6513 13096 6547
rect 13130 6513 13136 6547
rect 13090 6475 13136 6513
rect 13090 6441 13096 6475
rect 13130 6441 13136 6475
rect 13090 6403 13136 6441
rect 13090 6369 13096 6403
rect 13130 6369 13136 6403
rect 13090 6331 13136 6369
rect 13090 6297 13096 6331
rect 13130 6297 13136 6331
rect 13090 6259 13136 6297
rect 13090 6225 13096 6259
rect 13130 6225 13136 6259
rect 13090 6187 13136 6225
rect 13090 6153 13096 6187
rect 13130 6153 13136 6187
rect 13090 6115 13136 6153
rect 13090 6081 13096 6115
rect 13130 6081 13136 6115
rect 13090 6043 13136 6081
rect 13090 6009 13096 6043
rect 13130 6009 13136 6043
rect 13090 5971 13136 6009
rect 13090 5937 13096 5971
rect 13130 5937 13136 5971
rect 13090 5899 13136 5937
rect 13090 5865 13096 5899
rect 13130 5865 13136 5899
rect 13090 5827 13136 5865
rect 13090 5793 13096 5827
rect 13130 5793 13136 5827
rect 13090 5755 13136 5793
rect 13090 5721 13096 5755
rect 13130 5721 13136 5755
rect 13090 5683 13136 5721
rect 13090 5649 13096 5683
rect 13130 5649 13136 5683
rect 13090 5611 13136 5649
rect 13090 5577 13096 5611
rect 13130 5577 13136 5611
rect 13090 5562 13136 5577
rect 13186 6547 13232 6562
rect 13186 6513 13192 6547
rect 13226 6513 13232 6547
rect 13186 6475 13232 6513
rect 13186 6441 13192 6475
rect 13226 6441 13232 6475
rect 13186 6403 13232 6441
rect 13186 6369 13192 6403
rect 13226 6369 13232 6403
rect 13186 6331 13232 6369
rect 13186 6297 13192 6331
rect 13226 6297 13232 6331
rect 13186 6259 13232 6297
rect 13186 6225 13192 6259
rect 13226 6225 13232 6259
rect 13186 6187 13232 6225
rect 13186 6153 13192 6187
rect 13226 6153 13232 6187
rect 13186 6115 13232 6153
rect 13186 6081 13192 6115
rect 13226 6081 13232 6115
rect 13186 6043 13232 6081
rect 13186 6009 13192 6043
rect 13226 6009 13232 6043
rect 13186 5971 13232 6009
rect 13186 5937 13192 5971
rect 13226 5937 13232 5971
rect 13186 5899 13232 5937
rect 13186 5865 13192 5899
rect 13226 5865 13232 5899
rect 13186 5827 13232 5865
rect 13186 5793 13192 5827
rect 13226 5793 13232 5827
rect 13186 5755 13232 5793
rect 13186 5721 13192 5755
rect 13226 5721 13232 5755
rect 13186 5683 13232 5721
rect 13186 5649 13192 5683
rect 13226 5649 13232 5683
rect 13186 5611 13232 5649
rect 13186 5577 13192 5611
rect 13226 5577 13232 5611
rect 13186 5562 13232 5577
rect 13282 6547 13328 6562
rect 13282 6513 13288 6547
rect 13322 6513 13328 6547
rect 13282 6475 13328 6513
rect 13282 6441 13288 6475
rect 13322 6441 13328 6475
rect 13282 6403 13328 6441
rect 13282 6369 13288 6403
rect 13322 6369 13328 6403
rect 13282 6331 13328 6369
rect 13282 6297 13288 6331
rect 13322 6297 13328 6331
rect 13282 6259 13328 6297
rect 13282 6225 13288 6259
rect 13322 6225 13328 6259
rect 13282 6187 13328 6225
rect 13282 6153 13288 6187
rect 13322 6153 13328 6187
rect 13282 6115 13328 6153
rect 13282 6081 13288 6115
rect 13322 6081 13328 6115
rect 13282 6043 13328 6081
rect 13282 6009 13288 6043
rect 13322 6009 13328 6043
rect 13282 5971 13328 6009
rect 13282 5937 13288 5971
rect 13322 5937 13328 5971
rect 13282 5899 13328 5937
rect 13282 5865 13288 5899
rect 13322 5865 13328 5899
rect 13282 5827 13328 5865
rect 13282 5793 13288 5827
rect 13322 5793 13328 5827
rect 13282 5755 13328 5793
rect 13282 5721 13288 5755
rect 13322 5721 13328 5755
rect 13282 5683 13328 5721
rect 13282 5649 13288 5683
rect 13322 5649 13328 5683
rect 13282 5611 13328 5649
rect 13282 5577 13288 5611
rect 13322 5577 13328 5611
rect 13282 5562 13328 5577
rect 13378 6547 13424 6562
rect 13378 6513 13384 6547
rect 13418 6513 13424 6547
rect 13378 6475 13424 6513
rect 13378 6441 13384 6475
rect 13418 6441 13424 6475
rect 13378 6403 13424 6441
rect 13378 6369 13384 6403
rect 13418 6369 13424 6403
rect 13378 6331 13424 6369
rect 13378 6297 13384 6331
rect 13418 6297 13424 6331
rect 13378 6259 13424 6297
rect 13378 6225 13384 6259
rect 13418 6225 13424 6259
rect 13378 6187 13424 6225
rect 13378 6153 13384 6187
rect 13418 6153 13424 6187
rect 13378 6115 13424 6153
rect 13378 6081 13384 6115
rect 13418 6081 13424 6115
rect 13378 6043 13424 6081
rect 13378 6009 13384 6043
rect 13418 6009 13424 6043
rect 13378 5971 13424 6009
rect 13378 5937 13384 5971
rect 13418 5937 13424 5971
rect 13378 5899 13424 5937
rect 13378 5865 13384 5899
rect 13418 5865 13424 5899
rect 13378 5827 13424 5865
rect 13378 5793 13384 5827
rect 13418 5793 13424 5827
rect 13378 5755 13424 5793
rect 13378 5721 13384 5755
rect 13418 5721 13424 5755
rect 13378 5683 13424 5721
rect 13378 5649 13384 5683
rect 13418 5649 13424 5683
rect 13378 5611 13424 5649
rect 13378 5577 13384 5611
rect 13418 5577 13424 5611
rect 13378 5562 13424 5577
rect 13474 6547 13520 6562
rect 13474 6513 13480 6547
rect 13514 6513 13520 6547
rect 13474 6475 13520 6513
rect 13474 6441 13480 6475
rect 13514 6441 13520 6475
rect 13474 6403 13520 6441
rect 13474 6369 13480 6403
rect 13514 6369 13520 6403
rect 13474 6331 13520 6369
rect 13474 6297 13480 6331
rect 13514 6297 13520 6331
rect 13474 6259 13520 6297
rect 13474 6225 13480 6259
rect 13514 6225 13520 6259
rect 13474 6187 13520 6225
rect 13474 6153 13480 6187
rect 13514 6153 13520 6187
rect 13474 6115 13520 6153
rect 13474 6081 13480 6115
rect 13514 6081 13520 6115
rect 13474 6043 13520 6081
rect 13474 6009 13480 6043
rect 13514 6009 13520 6043
rect 13474 5971 13520 6009
rect 13474 5937 13480 5971
rect 13514 5937 13520 5971
rect 13474 5899 13520 5937
rect 13474 5865 13480 5899
rect 13514 5865 13520 5899
rect 13474 5827 13520 5865
rect 13474 5793 13480 5827
rect 13514 5793 13520 5827
rect 13474 5755 13520 5793
rect 13474 5721 13480 5755
rect 13514 5721 13520 5755
rect 13474 5683 13520 5721
rect 13474 5649 13480 5683
rect 13514 5649 13520 5683
rect 13474 5611 13520 5649
rect 13474 5577 13480 5611
rect 13514 5577 13520 5611
rect 13474 5562 13520 5577
rect 13570 6547 13616 6562
rect 13570 6513 13576 6547
rect 13610 6513 13616 6547
rect 13570 6475 13616 6513
rect 13570 6441 13576 6475
rect 13610 6441 13616 6475
rect 13570 6403 13616 6441
rect 13570 6369 13576 6403
rect 13610 6369 13616 6403
rect 13570 6331 13616 6369
rect 13570 6297 13576 6331
rect 13610 6297 13616 6331
rect 13570 6259 13616 6297
rect 13570 6225 13576 6259
rect 13610 6225 13616 6259
rect 13570 6187 13616 6225
rect 13570 6153 13576 6187
rect 13610 6153 13616 6187
rect 13570 6115 13616 6153
rect 13570 6081 13576 6115
rect 13610 6081 13616 6115
rect 13570 6043 13616 6081
rect 13570 6009 13576 6043
rect 13610 6009 13616 6043
rect 13570 5971 13616 6009
rect 13570 5937 13576 5971
rect 13610 5937 13616 5971
rect 13570 5899 13616 5937
rect 13570 5865 13576 5899
rect 13610 5865 13616 5899
rect 13570 5827 13616 5865
rect 13570 5793 13576 5827
rect 13610 5793 13616 5827
rect 13570 5755 13616 5793
rect 13570 5721 13576 5755
rect 13610 5721 13616 5755
rect 13570 5683 13616 5721
rect 13570 5649 13576 5683
rect 13610 5649 13616 5683
rect 13570 5611 13616 5649
rect 13570 5577 13576 5611
rect 13610 5577 13616 5611
rect 13570 5562 13616 5577
rect 14184 6543 14230 6558
rect 14184 6509 14190 6543
rect 14224 6509 14230 6543
rect 14184 6471 14230 6509
rect 14184 6437 14190 6471
rect 14224 6437 14230 6471
rect 14184 6399 14230 6437
rect 14184 6365 14190 6399
rect 14224 6365 14230 6399
rect 14184 6327 14230 6365
rect 14184 6293 14190 6327
rect 14224 6293 14230 6327
rect 14184 6255 14230 6293
rect 14184 6221 14190 6255
rect 14224 6221 14230 6255
rect 14184 6183 14230 6221
rect 14184 6149 14190 6183
rect 14224 6149 14230 6183
rect 14184 6111 14230 6149
rect 14184 6077 14190 6111
rect 14224 6077 14230 6111
rect 14184 6039 14230 6077
rect 14184 6005 14190 6039
rect 14224 6005 14230 6039
rect 14184 5967 14230 6005
rect 14184 5933 14190 5967
rect 14224 5933 14230 5967
rect 14184 5895 14230 5933
rect 14184 5861 14190 5895
rect 14224 5861 14230 5895
rect 14184 5823 14230 5861
rect 14184 5789 14190 5823
rect 14224 5789 14230 5823
rect 14184 5751 14230 5789
rect 14184 5717 14190 5751
rect 14224 5717 14230 5751
rect 14184 5679 14230 5717
rect 14184 5645 14190 5679
rect 14224 5645 14230 5679
rect 14184 5607 14230 5645
rect 14184 5573 14190 5607
rect 14224 5573 14230 5607
rect 14184 5558 14230 5573
rect 14280 6543 14326 6558
rect 14280 6509 14286 6543
rect 14320 6509 14326 6543
rect 14280 6471 14326 6509
rect 14280 6437 14286 6471
rect 14320 6437 14326 6471
rect 14280 6399 14326 6437
rect 14280 6365 14286 6399
rect 14320 6365 14326 6399
rect 14280 6327 14326 6365
rect 14280 6293 14286 6327
rect 14320 6293 14326 6327
rect 14280 6255 14326 6293
rect 14280 6221 14286 6255
rect 14320 6221 14326 6255
rect 14280 6183 14326 6221
rect 14280 6149 14286 6183
rect 14320 6149 14326 6183
rect 14280 6111 14326 6149
rect 14280 6077 14286 6111
rect 14320 6077 14326 6111
rect 14280 6039 14326 6077
rect 14280 6005 14286 6039
rect 14320 6005 14326 6039
rect 14280 5967 14326 6005
rect 14280 5933 14286 5967
rect 14320 5933 14326 5967
rect 14280 5895 14326 5933
rect 14280 5861 14286 5895
rect 14320 5861 14326 5895
rect 14280 5823 14326 5861
rect 14280 5789 14286 5823
rect 14320 5789 14326 5823
rect 14280 5751 14326 5789
rect 14280 5717 14286 5751
rect 14320 5717 14326 5751
rect 14280 5679 14326 5717
rect 14280 5645 14286 5679
rect 14320 5645 14326 5679
rect 14280 5607 14326 5645
rect 14280 5573 14286 5607
rect 14320 5573 14326 5607
rect 14280 5558 14326 5573
rect 14376 6543 14422 6558
rect 14376 6509 14382 6543
rect 14416 6509 14422 6543
rect 14376 6471 14422 6509
rect 14376 6437 14382 6471
rect 14416 6437 14422 6471
rect 14376 6399 14422 6437
rect 14376 6365 14382 6399
rect 14416 6365 14422 6399
rect 14376 6327 14422 6365
rect 14376 6293 14382 6327
rect 14416 6293 14422 6327
rect 14376 6255 14422 6293
rect 14376 6221 14382 6255
rect 14416 6221 14422 6255
rect 14376 6183 14422 6221
rect 14376 6149 14382 6183
rect 14416 6149 14422 6183
rect 14376 6111 14422 6149
rect 14376 6077 14382 6111
rect 14416 6077 14422 6111
rect 14376 6039 14422 6077
rect 14376 6005 14382 6039
rect 14416 6005 14422 6039
rect 14376 5967 14422 6005
rect 14376 5933 14382 5967
rect 14416 5933 14422 5967
rect 14376 5895 14422 5933
rect 14376 5861 14382 5895
rect 14416 5861 14422 5895
rect 14376 5823 14422 5861
rect 14376 5789 14382 5823
rect 14416 5789 14422 5823
rect 14376 5751 14422 5789
rect 14376 5717 14382 5751
rect 14416 5717 14422 5751
rect 14376 5679 14422 5717
rect 14376 5645 14382 5679
rect 14416 5645 14422 5679
rect 14376 5607 14422 5645
rect 14376 5573 14382 5607
rect 14416 5573 14422 5607
rect 14376 5558 14422 5573
rect 14472 6543 14518 6558
rect 14472 6509 14478 6543
rect 14512 6509 14518 6543
rect 14472 6471 14518 6509
rect 14472 6437 14478 6471
rect 14512 6437 14518 6471
rect 14472 6399 14518 6437
rect 14472 6365 14478 6399
rect 14512 6365 14518 6399
rect 14472 6327 14518 6365
rect 14472 6293 14478 6327
rect 14512 6293 14518 6327
rect 14472 6255 14518 6293
rect 14472 6221 14478 6255
rect 14512 6221 14518 6255
rect 14472 6183 14518 6221
rect 14472 6149 14478 6183
rect 14512 6149 14518 6183
rect 14472 6111 14518 6149
rect 14472 6077 14478 6111
rect 14512 6077 14518 6111
rect 14472 6039 14518 6077
rect 14472 6005 14478 6039
rect 14512 6005 14518 6039
rect 14472 5967 14518 6005
rect 14472 5933 14478 5967
rect 14512 5933 14518 5967
rect 14472 5895 14518 5933
rect 14472 5861 14478 5895
rect 14512 5861 14518 5895
rect 14472 5823 14518 5861
rect 14472 5789 14478 5823
rect 14512 5789 14518 5823
rect 14472 5751 14518 5789
rect 14472 5717 14478 5751
rect 14512 5717 14518 5751
rect 14472 5679 14518 5717
rect 14472 5645 14478 5679
rect 14512 5645 14518 5679
rect 14472 5607 14518 5645
rect 14472 5573 14478 5607
rect 14512 5573 14518 5607
rect 14472 5558 14518 5573
rect 14568 6543 14614 6558
rect 14568 6509 14574 6543
rect 14608 6509 14614 6543
rect 14568 6471 14614 6509
rect 14568 6437 14574 6471
rect 14608 6437 14614 6471
rect 14568 6399 14614 6437
rect 14568 6365 14574 6399
rect 14608 6365 14614 6399
rect 14568 6327 14614 6365
rect 14568 6293 14574 6327
rect 14608 6293 14614 6327
rect 14568 6255 14614 6293
rect 14568 6221 14574 6255
rect 14608 6221 14614 6255
rect 14568 6183 14614 6221
rect 14568 6149 14574 6183
rect 14608 6149 14614 6183
rect 14568 6111 14614 6149
rect 14568 6077 14574 6111
rect 14608 6077 14614 6111
rect 14568 6039 14614 6077
rect 14568 6005 14574 6039
rect 14608 6005 14614 6039
rect 14568 5967 14614 6005
rect 14568 5933 14574 5967
rect 14608 5933 14614 5967
rect 14568 5895 14614 5933
rect 14568 5861 14574 5895
rect 14608 5861 14614 5895
rect 14568 5823 14614 5861
rect 14568 5789 14574 5823
rect 14608 5789 14614 5823
rect 14568 5751 14614 5789
rect 14568 5717 14574 5751
rect 14608 5717 14614 5751
rect 14568 5679 14614 5717
rect 14568 5645 14574 5679
rect 14608 5645 14614 5679
rect 14568 5607 14614 5645
rect 14568 5573 14574 5607
rect 14608 5573 14614 5607
rect 14568 5558 14614 5573
rect 14664 6543 14710 6558
rect 14664 6509 14670 6543
rect 14704 6509 14710 6543
rect 14664 6471 14710 6509
rect 14664 6437 14670 6471
rect 14704 6437 14710 6471
rect 14664 6399 14710 6437
rect 14664 6365 14670 6399
rect 14704 6365 14710 6399
rect 14664 6327 14710 6365
rect 14664 6293 14670 6327
rect 14704 6293 14710 6327
rect 14664 6255 14710 6293
rect 14664 6221 14670 6255
rect 14704 6221 14710 6255
rect 14664 6183 14710 6221
rect 14664 6149 14670 6183
rect 14704 6149 14710 6183
rect 14664 6111 14710 6149
rect 14664 6077 14670 6111
rect 14704 6077 14710 6111
rect 14664 6039 14710 6077
rect 14664 6005 14670 6039
rect 14704 6005 14710 6039
rect 14664 5967 14710 6005
rect 14664 5933 14670 5967
rect 14704 5933 14710 5967
rect 14664 5895 14710 5933
rect 14664 5861 14670 5895
rect 14704 5861 14710 5895
rect 14664 5823 14710 5861
rect 14664 5789 14670 5823
rect 14704 5789 14710 5823
rect 14664 5751 14710 5789
rect 14664 5717 14670 5751
rect 14704 5717 14710 5751
rect 14664 5679 14710 5717
rect 14664 5645 14670 5679
rect 14704 5645 14710 5679
rect 14664 5607 14710 5645
rect 14664 5573 14670 5607
rect 14704 5573 14710 5607
rect 14664 5558 14710 5573
rect 14760 6543 14806 6558
rect 14760 6509 14766 6543
rect 14800 6509 14806 6543
rect 14760 6471 14806 6509
rect 14760 6437 14766 6471
rect 14800 6437 14806 6471
rect 14760 6399 14806 6437
rect 14760 6365 14766 6399
rect 14800 6365 14806 6399
rect 14760 6327 14806 6365
rect 14760 6293 14766 6327
rect 14800 6293 14806 6327
rect 14760 6255 14806 6293
rect 14760 6221 14766 6255
rect 14800 6221 14806 6255
rect 14760 6183 14806 6221
rect 14760 6149 14766 6183
rect 14800 6149 14806 6183
rect 14760 6111 14806 6149
rect 14760 6077 14766 6111
rect 14800 6077 14806 6111
rect 14760 6039 14806 6077
rect 14760 6005 14766 6039
rect 14800 6005 14806 6039
rect 14760 5967 14806 6005
rect 14760 5933 14766 5967
rect 14800 5933 14806 5967
rect 14760 5895 14806 5933
rect 14760 5861 14766 5895
rect 14800 5861 14806 5895
rect 14760 5823 14806 5861
rect 14760 5789 14766 5823
rect 14800 5789 14806 5823
rect 14760 5751 14806 5789
rect 14760 5717 14766 5751
rect 14800 5717 14806 5751
rect 14760 5679 14806 5717
rect 14760 5645 14766 5679
rect 14800 5645 14806 5679
rect 14760 5607 14806 5645
rect 14760 5573 14766 5607
rect 14800 5573 14806 5607
rect 14760 5558 14806 5573
rect 14856 6543 14902 6558
rect 14856 6509 14862 6543
rect 14896 6509 14902 6543
rect 14856 6471 14902 6509
rect 14856 6437 14862 6471
rect 14896 6437 14902 6471
rect 14856 6399 14902 6437
rect 14856 6365 14862 6399
rect 14896 6365 14902 6399
rect 14856 6327 14902 6365
rect 14856 6293 14862 6327
rect 14896 6293 14902 6327
rect 14856 6255 14902 6293
rect 14856 6221 14862 6255
rect 14896 6221 14902 6255
rect 14856 6183 14902 6221
rect 14856 6149 14862 6183
rect 14896 6149 14902 6183
rect 14856 6111 14902 6149
rect 14856 6077 14862 6111
rect 14896 6077 14902 6111
rect 14856 6039 14902 6077
rect 14856 6005 14862 6039
rect 14896 6005 14902 6039
rect 14856 5967 14902 6005
rect 14856 5933 14862 5967
rect 14896 5933 14902 5967
rect 14856 5895 14902 5933
rect 14856 5861 14862 5895
rect 14896 5861 14902 5895
rect 14856 5823 14902 5861
rect 14856 5789 14862 5823
rect 14896 5789 14902 5823
rect 14856 5751 14902 5789
rect 14856 5717 14862 5751
rect 14896 5717 14902 5751
rect 14856 5679 14902 5717
rect 14856 5645 14862 5679
rect 14896 5645 14902 5679
rect 14856 5607 14902 5645
rect 14856 5573 14862 5607
rect 14896 5573 14902 5607
rect 14856 5558 14902 5573
rect 14952 6543 14998 6558
rect 14952 6509 14958 6543
rect 14992 6509 14998 6543
rect 14952 6471 14998 6509
rect 14952 6437 14958 6471
rect 14992 6437 14998 6471
rect 14952 6399 14998 6437
rect 14952 6365 14958 6399
rect 14992 6365 14998 6399
rect 14952 6327 14998 6365
rect 14952 6293 14958 6327
rect 14992 6293 14998 6327
rect 14952 6255 14998 6293
rect 14952 6221 14958 6255
rect 14992 6221 14998 6255
rect 14952 6183 14998 6221
rect 14952 6149 14958 6183
rect 14992 6149 14998 6183
rect 14952 6111 14998 6149
rect 15592 6182 15666 7832
rect 15592 6148 15614 6182
rect 15648 6148 15666 6182
rect 15592 6126 15666 6148
rect 14952 6077 14958 6111
rect 14992 6077 14998 6111
rect 14952 6039 14998 6077
rect 14952 6005 14958 6039
rect 14992 6005 14998 6039
rect 14952 5967 14998 6005
rect 14952 5933 14958 5967
rect 14992 5933 14998 5967
rect 14952 5895 14998 5933
rect 14952 5861 14958 5895
rect 14992 5861 14998 5895
rect 14952 5823 14998 5861
rect 14952 5789 14958 5823
rect 14992 5789 14998 5823
rect 14952 5751 14998 5789
rect 14952 5717 14958 5751
rect 14992 5717 14998 5751
rect 14952 5679 14998 5717
rect 14952 5645 14958 5679
rect 14992 5645 14998 5679
rect 14952 5607 14998 5645
rect 14952 5573 14958 5607
rect 14992 5573 14998 5607
rect 14952 5558 14998 5573
rect 15512 5879 15558 5926
rect 15512 5845 15518 5879
rect 15552 5845 15558 5879
rect 15512 5807 15558 5845
rect 15512 5773 15518 5807
rect 15552 5773 15558 5807
rect 15512 5735 15558 5773
rect 15512 5701 15518 5735
rect 15552 5701 15558 5735
rect 15512 5663 15558 5701
rect 15512 5629 15518 5663
rect 15552 5629 15558 5663
rect 15512 5591 15558 5629
rect 15512 5557 15518 5591
rect 15552 5557 15558 5591
rect 15512 5519 15558 5557
rect 15512 5485 15518 5519
rect 15552 5485 15558 5519
rect 15512 5447 15558 5485
rect 864 5420 2408 5430
rect 858 5418 2408 5420
rect 858 5372 880 5418
rect 982 5372 2278 5418
rect 2380 5372 2408 5418
rect 3806 5408 5364 5414
rect 858 5190 2408 5372
rect 3802 5400 5364 5408
rect 3802 5354 3824 5400
rect 3926 5398 5364 5400
rect 3926 5354 5234 5398
rect 3802 5352 5234 5354
rect 5336 5352 5364 5398
rect 3802 5248 5364 5352
rect 1570 5124 1624 5190
rect 3800 5164 5364 5248
rect 6828 5402 8396 5420
rect 6828 5398 8268 5402
rect 6828 5352 6854 5398
rect 6956 5356 8268 5398
rect 8370 5356 8396 5402
rect 6956 5352 8396 5356
rect 6828 5170 8396 5352
rect 9920 5398 11494 5414
rect 9920 5392 11354 5398
rect 9920 5346 9950 5392
rect 10052 5352 11354 5392
rect 11456 5352 11494 5398
rect 15512 5413 15518 5447
rect 15552 5413 15558 5447
rect 13096 5380 14650 5386
rect 10052 5346 11494 5352
rect 1570 5090 1580 5124
rect 1614 5090 1624 5124
rect 1570 5074 1624 5090
rect 4526 5108 4580 5164
rect 4526 5074 4536 5108
rect 4570 5074 4580 5108
rect 4526 5058 4580 5074
rect 7556 5108 7610 5170
rect 9920 5156 11494 5346
rect 13070 5372 14650 5380
rect 13070 5366 14510 5372
rect 13070 5320 13094 5366
rect 13196 5326 14510 5366
rect 14612 5326 14650 5372
rect 13196 5320 14650 5326
rect 7556 5074 7566 5108
rect 7600 5074 7610 5108
rect 7556 5058 7610 5074
rect 10644 5106 10698 5156
rect 13070 5122 14650 5320
rect 15512 5375 15558 5413
rect 15512 5341 15518 5375
rect 15552 5341 15558 5375
rect 15512 5303 15558 5341
rect 15512 5269 15518 5303
rect 15552 5269 15558 5303
rect 15512 5231 15558 5269
rect 15512 5197 15518 5231
rect 15552 5197 15558 5231
rect 15512 5159 15558 5197
rect 15512 5125 15518 5159
rect 15552 5125 15558 5159
rect 10644 5072 10654 5106
rect 10688 5072 10698 5106
rect 10644 5056 10698 5072
rect 13800 5080 13854 5122
rect 13800 5046 13810 5080
rect 13844 5046 13854 5080
rect 13800 5030 13854 5046
rect 15512 5087 15558 5125
rect 15512 5053 15518 5087
rect 15552 5053 15558 5087
rect 15512 5015 15558 5053
rect 15512 4981 15518 5015
rect 15552 4981 15558 5015
rect -1126 4769 -402 4792
rect -1126 4735 -1067 4769
rect -1033 4735 -402 4769
rect -1126 4630 -402 4735
rect 1478 4929 1524 4944
rect 1478 4895 1484 4929
rect 1518 4895 1524 4929
rect 1478 4857 1524 4895
rect 1478 4823 1484 4857
rect 1518 4823 1524 4857
rect 1478 4785 1524 4823
rect 1478 4751 1484 4785
rect 1518 4751 1524 4785
rect 1478 4713 1524 4751
rect 1478 4679 1484 4713
rect 1518 4679 1524 4713
rect 1478 4641 1524 4679
rect -23592 4427 -23546 4442
rect -23592 4393 -23586 4427
rect -23552 4393 -23546 4427
rect -23592 4355 -23546 4393
rect -23592 4321 -23586 4355
rect -23552 4321 -23546 4355
rect -23592 4283 -23546 4321
rect -23592 4249 -23586 4283
rect -23552 4249 -23546 4283
rect -23592 4211 -23546 4249
rect -23592 4177 -23586 4211
rect -23552 4177 -23546 4211
rect -23592 4139 -23546 4177
rect -23592 4105 -23586 4139
rect -23552 4105 -23546 4139
rect -23592 4067 -23546 4105
rect -23592 4033 -23586 4067
rect -23552 4033 -23546 4067
rect -23592 3995 -23546 4033
rect -23592 3961 -23586 3995
rect -23552 3961 -23546 3995
rect -23592 3923 -23546 3961
rect -23592 3889 -23586 3923
rect -23552 3889 -23546 3923
rect -23592 3851 -23546 3889
rect -23592 3817 -23586 3851
rect -23552 3817 -23546 3851
rect -23592 3779 -23546 3817
rect -23592 3745 -23586 3779
rect -23552 3745 -23546 3779
rect -23592 3707 -23546 3745
rect -23592 3673 -23586 3707
rect -23552 3673 -23546 3707
rect -23592 3635 -23546 3673
rect -23592 3601 -23586 3635
rect -23552 3601 -23546 3635
rect -23592 3563 -23546 3601
rect -23592 3529 -23586 3563
rect -23552 3529 -23546 3563
rect -23592 3491 -23546 3529
rect -23592 3457 -23586 3491
rect -23552 3457 -23546 3491
rect -23592 3442 -23546 3457
rect -23496 4427 -23450 4442
rect -23496 4393 -23490 4427
rect -23456 4393 -23450 4427
rect -23496 4355 -23450 4393
rect -23496 4321 -23490 4355
rect -23456 4321 -23450 4355
rect -23496 4283 -23450 4321
rect -23496 4249 -23490 4283
rect -23456 4249 -23450 4283
rect -23496 4211 -23450 4249
rect -23496 4177 -23490 4211
rect -23456 4177 -23450 4211
rect -23496 4139 -23450 4177
rect -23496 4105 -23490 4139
rect -23456 4105 -23450 4139
rect -23496 4067 -23450 4105
rect -23496 4033 -23490 4067
rect -23456 4033 -23450 4067
rect -23496 3995 -23450 4033
rect -23496 3961 -23490 3995
rect -23456 3961 -23450 3995
rect -23496 3923 -23450 3961
rect -23496 3889 -23490 3923
rect -23456 3889 -23450 3923
rect -23496 3851 -23450 3889
rect -23496 3817 -23490 3851
rect -23456 3817 -23450 3851
rect -23496 3779 -23450 3817
rect -23496 3745 -23490 3779
rect -23456 3745 -23450 3779
rect -23496 3707 -23450 3745
rect -23496 3673 -23490 3707
rect -23456 3673 -23450 3707
rect -23496 3635 -23450 3673
rect -23496 3601 -23490 3635
rect -23456 3601 -23450 3635
rect -23496 3563 -23450 3601
rect -23496 3529 -23490 3563
rect -23456 3529 -23450 3563
rect -23496 3491 -23450 3529
rect -23496 3457 -23490 3491
rect -23456 3457 -23450 3491
rect -23496 3442 -23450 3457
rect -23400 4427 -23354 4442
rect -23400 4393 -23394 4427
rect -23360 4393 -23354 4427
rect -23400 4355 -23354 4393
rect -23400 4321 -23394 4355
rect -23360 4321 -23354 4355
rect -23400 4283 -23354 4321
rect -23400 4249 -23394 4283
rect -23360 4249 -23354 4283
rect -23400 4211 -23354 4249
rect -23400 4177 -23394 4211
rect -23360 4177 -23354 4211
rect -23400 4139 -23354 4177
rect -23400 4105 -23394 4139
rect -23360 4105 -23354 4139
rect -23400 4067 -23354 4105
rect -23400 4033 -23394 4067
rect -23360 4033 -23354 4067
rect -23400 3995 -23354 4033
rect -23400 3961 -23394 3995
rect -23360 3961 -23354 3995
rect -23400 3923 -23354 3961
rect -23400 3889 -23394 3923
rect -23360 3889 -23354 3923
rect -23400 3851 -23354 3889
rect -23400 3817 -23394 3851
rect -23360 3817 -23354 3851
rect -23400 3779 -23354 3817
rect -23400 3745 -23394 3779
rect -23360 3745 -23354 3779
rect -23400 3707 -23354 3745
rect -23400 3673 -23394 3707
rect -23360 3673 -23354 3707
rect -23400 3635 -23354 3673
rect -23400 3601 -23394 3635
rect -23360 3601 -23354 3635
rect -23400 3563 -23354 3601
rect -23400 3529 -23394 3563
rect -23360 3529 -23354 3563
rect -23400 3491 -23354 3529
rect -23400 3457 -23394 3491
rect -23360 3457 -23354 3491
rect -23400 3442 -23354 3457
rect -23304 4427 -23258 4442
rect -23304 4393 -23298 4427
rect -23264 4393 -23258 4427
rect -23304 4355 -23258 4393
rect -23304 4321 -23298 4355
rect -23264 4321 -23258 4355
rect -23304 4283 -23258 4321
rect -23304 4249 -23298 4283
rect -23264 4249 -23258 4283
rect -23304 4211 -23258 4249
rect -23304 4177 -23298 4211
rect -23264 4177 -23258 4211
rect -23304 4139 -23258 4177
rect -23304 4105 -23298 4139
rect -23264 4105 -23258 4139
rect -23304 4067 -23258 4105
rect -23304 4033 -23298 4067
rect -23264 4033 -23258 4067
rect -23304 3995 -23258 4033
rect -23304 3961 -23298 3995
rect -23264 3961 -23258 3995
rect -23304 3923 -23258 3961
rect -23304 3889 -23298 3923
rect -23264 3889 -23258 3923
rect -23304 3851 -23258 3889
rect -23304 3817 -23298 3851
rect -23264 3817 -23258 3851
rect -23304 3779 -23258 3817
rect -23304 3745 -23298 3779
rect -23264 3745 -23258 3779
rect -23304 3707 -23258 3745
rect -23304 3673 -23298 3707
rect -23264 3673 -23258 3707
rect -23304 3635 -23258 3673
rect -23304 3601 -23298 3635
rect -23264 3601 -23258 3635
rect -23304 3563 -23258 3601
rect -23304 3529 -23298 3563
rect -23264 3529 -23258 3563
rect -23304 3491 -23258 3529
rect -23304 3457 -23298 3491
rect -23264 3457 -23258 3491
rect -23304 3442 -23258 3457
rect -23208 4427 -23162 4442
rect -23208 4393 -23202 4427
rect -23168 4393 -23162 4427
rect -23208 4355 -23162 4393
rect -23208 4321 -23202 4355
rect -23168 4321 -23162 4355
rect -23208 4283 -23162 4321
rect -23208 4249 -23202 4283
rect -23168 4249 -23162 4283
rect -23208 4211 -23162 4249
rect -23208 4177 -23202 4211
rect -23168 4177 -23162 4211
rect -23208 4139 -23162 4177
rect -23208 4105 -23202 4139
rect -23168 4105 -23162 4139
rect -23208 4067 -23162 4105
rect -23208 4033 -23202 4067
rect -23168 4033 -23162 4067
rect -23208 3995 -23162 4033
rect -23208 3961 -23202 3995
rect -23168 3961 -23162 3995
rect -23208 3923 -23162 3961
rect -23208 3889 -23202 3923
rect -23168 3889 -23162 3923
rect -23208 3851 -23162 3889
rect -23208 3817 -23202 3851
rect -23168 3817 -23162 3851
rect -23208 3779 -23162 3817
rect -23208 3745 -23202 3779
rect -23168 3745 -23162 3779
rect -23208 3707 -23162 3745
rect -23208 3673 -23202 3707
rect -23168 3673 -23162 3707
rect -23208 3635 -23162 3673
rect -23208 3601 -23202 3635
rect -23168 3601 -23162 3635
rect -23208 3563 -23162 3601
rect -23208 3529 -23202 3563
rect -23168 3529 -23162 3563
rect -23208 3491 -23162 3529
rect -23208 3457 -23202 3491
rect -23168 3457 -23162 3491
rect -23208 3442 -23162 3457
rect -23112 4427 -23066 4442
rect -23112 4393 -23106 4427
rect -23072 4393 -23066 4427
rect -23112 4355 -23066 4393
rect -23112 4321 -23106 4355
rect -23072 4321 -23066 4355
rect -23112 4283 -23066 4321
rect -23112 4249 -23106 4283
rect -23072 4249 -23066 4283
rect -23112 4211 -23066 4249
rect -23112 4177 -23106 4211
rect -23072 4177 -23066 4211
rect -23112 4139 -23066 4177
rect -23112 4105 -23106 4139
rect -23072 4105 -23066 4139
rect -23112 4067 -23066 4105
rect -23112 4033 -23106 4067
rect -23072 4033 -23066 4067
rect -23112 3995 -23066 4033
rect -23112 3961 -23106 3995
rect -23072 3961 -23066 3995
rect -23112 3923 -23066 3961
rect -23112 3889 -23106 3923
rect -23072 3889 -23066 3923
rect -23112 3851 -23066 3889
rect -23112 3817 -23106 3851
rect -23072 3817 -23066 3851
rect -23112 3779 -23066 3817
rect -23112 3745 -23106 3779
rect -23072 3745 -23066 3779
rect -23112 3707 -23066 3745
rect -23112 3673 -23106 3707
rect -23072 3673 -23066 3707
rect -23112 3635 -23066 3673
rect -23112 3601 -23106 3635
rect -23072 3601 -23066 3635
rect -23112 3563 -23066 3601
rect -23112 3529 -23106 3563
rect -23072 3529 -23066 3563
rect -23112 3491 -23066 3529
rect -23112 3457 -23106 3491
rect -23072 3457 -23066 3491
rect -23112 3442 -23066 3457
rect -23016 4427 -22970 4442
rect -23016 4393 -23010 4427
rect -22976 4393 -22970 4427
rect -23016 4355 -22970 4393
rect -23016 4321 -23010 4355
rect -22976 4321 -22970 4355
rect -23016 4283 -22970 4321
rect -23016 4249 -23010 4283
rect -22976 4249 -22970 4283
rect -23016 4211 -22970 4249
rect -23016 4177 -23010 4211
rect -22976 4177 -22970 4211
rect -23016 4139 -22970 4177
rect -23016 4105 -23010 4139
rect -22976 4105 -22970 4139
rect -23016 4067 -22970 4105
rect -23016 4033 -23010 4067
rect -22976 4033 -22970 4067
rect -23016 3995 -22970 4033
rect -23016 3961 -23010 3995
rect -22976 3961 -22970 3995
rect -23016 3923 -22970 3961
rect -23016 3889 -23010 3923
rect -22976 3889 -22970 3923
rect -23016 3851 -22970 3889
rect -23016 3817 -23010 3851
rect -22976 3817 -22970 3851
rect -23016 3779 -22970 3817
rect -23016 3745 -23010 3779
rect -22976 3745 -22970 3779
rect -23016 3707 -22970 3745
rect -23016 3673 -23010 3707
rect -22976 3673 -22970 3707
rect -23016 3635 -22970 3673
rect -23016 3601 -23010 3635
rect -22976 3601 -22970 3635
rect -23016 3563 -22970 3601
rect -23016 3529 -23010 3563
rect -22976 3529 -22970 3563
rect -23016 3491 -22970 3529
rect -23016 3457 -23010 3491
rect -22976 3457 -22970 3491
rect -23016 3442 -22970 3457
rect -22920 4427 -22874 4442
rect -22920 4393 -22914 4427
rect -22880 4393 -22874 4427
rect -22920 4355 -22874 4393
rect -22920 4321 -22914 4355
rect -22880 4321 -22874 4355
rect -22920 4283 -22874 4321
rect -22920 4249 -22914 4283
rect -22880 4249 -22874 4283
rect -22920 4211 -22874 4249
rect -22920 4177 -22914 4211
rect -22880 4177 -22874 4211
rect -22920 4139 -22874 4177
rect -22920 4105 -22914 4139
rect -22880 4105 -22874 4139
rect -22920 4067 -22874 4105
rect -22920 4033 -22914 4067
rect -22880 4033 -22874 4067
rect -22920 3995 -22874 4033
rect -22920 3961 -22914 3995
rect -22880 3961 -22874 3995
rect -22920 3923 -22874 3961
rect -22920 3889 -22914 3923
rect -22880 3889 -22874 3923
rect -22920 3851 -22874 3889
rect -22920 3817 -22914 3851
rect -22880 3817 -22874 3851
rect -22920 3779 -22874 3817
rect -22920 3745 -22914 3779
rect -22880 3745 -22874 3779
rect -22920 3707 -22874 3745
rect -22920 3673 -22914 3707
rect -22880 3673 -22874 3707
rect -22920 3635 -22874 3673
rect -22920 3601 -22914 3635
rect -22880 3601 -22874 3635
rect -22920 3563 -22874 3601
rect -22920 3529 -22914 3563
rect -22880 3529 -22874 3563
rect -22920 3491 -22874 3529
rect -22920 3457 -22914 3491
rect -22880 3457 -22874 3491
rect -22920 3442 -22874 3457
rect -22824 4427 -22778 4442
rect -22824 4393 -22818 4427
rect -22784 4393 -22778 4427
rect -22824 4355 -22778 4393
rect -22824 4321 -22818 4355
rect -22784 4321 -22778 4355
rect -22824 4283 -22778 4321
rect -22824 4249 -22818 4283
rect -22784 4249 -22778 4283
rect -22824 4211 -22778 4249
rect -22824 4177 -22818 4211
rect -22784 4177 -22778 4211
rect -22824 4139 -22778 4177
rect -22824 4105 -22818 4139
rect -22784 4105 -22778 4139
rect -22824 4067 -22778 4105
rect -22824 4033 -22818 4067
rect -22784 4033 -22778 4067
rect -22824 3995 -22778 4033
rect -22824 3961 -22818 3995
rect -22784 3961 -22778 3995
rect -22824 3923 -22778 3961
rect -22824 3889 -22818 3923
rect -22784 3889 -22778 3923
rect -22824 3851 -22778 3889
rect -22824 3817 -22818 3851
rect -22784 3817 -22778 3851
rect -22824 3779 -22778 3817
rect -22824 3745 -22818 3779
rect -22784 3745 -22778 3779
rect -22824 3707 -22778 3745
rect -22824 3673 -22818 3707
rect -22784 3673 -22778 3707
rect -22824 3635 -22778 3673
rect -22824 3601 -22818 3635
rect -22784 3601 -22778 3635
rect -22824 3563 -22778 3601
rect -22824 3529 -22818 3563
rect -22784 3529 -22778 3563
rect -22824 3491 -22778 3529
rect -22824 3457 -22818 3491
rect -22784 3457 -22778 3491
rect -22824 3442 -22778 3457
rect -22728 4427 -22682 4442
rect -22728 4393 -22722 4427
rect -22688 4393 -22682 4427
rect -22728 4355 -22682 4393
rect -22728 4321 -22722 4355
rect -22688 4321 -22682 4355
rect -22728 4283 -22682 4321
rect -22728 4249 -22722 4283
rect -22688 4249 -22682 4283
rect -22728 4211 -22682 4249
rect -22728 4177 -22722 4211
rect -22688 4177 -22682 4211
rect -22728 4139 -22682 4177
rect -22728 4105 -22722 4139
rect -22688 4105 -22682 4139
rect -22728 4067 -22682 4105
rect -22728 4033 -22722 4067
rect -22688 4033 -22682 4067
rect -22728 3995 -22682 4033
rect -22728 3961 -22722 3995
rect -22688 3961 -22682 3995
rect -22728 3923 -22682 3961
rect -22728 3889 -22722 3923
rect -22688 3889 -22682 3923
rect -22728 3851 -22682 3889
rect -22728 3817 -22722 3851
rect -22688 3817 -22682 3851
rect -22728 3779 -22682 3817
rect -22728 3745 -22722 3779
rect -22688 3745 -22682 3779
rect -22728 3707 -22682 3745
rect -22728 3673 -22722 3707
rect -22688 3673 -22682 3707
rect -22728 3635 -22682 3673
rect -22728 3601 -22722 3635
rect -22688 3601 -22682 3635
rect -22728 3563 -22682 3601
rect -22728 3529 -22722 3563
rect -22688 3529 -22682 3563
rect -22728 3491 -22682 3529
rect -22728 3457 -22722 3491
rect -22688 3457 -22682 3491
rect -22728 3442 -22682 3457
rect -22632 4427 -22586 4442
rect -22632 4393 -22626 4427
rect -22592 4393 -22586 4427
rect -22632 4355 -22586 4393
rect -22632 4321 -22626 4355
rect -22592 4321 -22586 4355
rect -22632 4283 -22586 4321
rect -22632 4249 -22626 4283
rect -22592 4249 -22586 4283
rect -22632 4211 -22586 4249
rect -22632 4177 -22626 4211
rect -22592 4177 -22586 4211
rect -22632 4139 -22586 4177
rect -22632 4105 -22626 4139
rect -22592 4105 -22586 4139
rect -22632 4067 -22586 4105
rect -22632 4033 -22626 4067
rect -22592 4033 -22586 4067
rect -22632 3995 -22586 4033
rect -22632 3961 -22626 3995
rect -22592 3961 -22586 3995
rect -22632 3923 -22586 3961
rect -22632 3889 -22626 3923
rect -22592 3889 -22586 3923
rect -22632 3851 -22586 3889
rect -22632 3817 -22626 3851
rect -22592 3817 -22586 3851
rect -22632 3779 -22586 3817
rect -22632 3745 -22626 3779
rect -22592 3745 -22586 3779
rect -22632 3707 -22586 3745
rect -22632 3673 -22626 3707
rect -22592 3673 -22586 3707
rect -22632 3635 -22586 3673
rect -22632 3601 -22626 3635
rect -22592 3601 -22586 3635
rect -22632 3563 -22586 3601
rect -22632 3529 -22626 3563
rect -22592 3529 -22586 3563
rect -22632 3491 -22586 3529
rect -22632 3457 -22626 3491
rect -22592 3457 -22586 3491
rect -22632 3442 -22586 3457
rect -22536 4427 -22490 4442
rect -22536 4393 -22530 4427
rect -22496 4393 -22490 4427
rect -22536 4355 -22490 4393
rect -22536 4321 -22530 4355
rect -22496 4321 -22490 4355
rect -22536 4283 -22490 4321
rect -22536 4249 -22530 4283
rect -22496 4249 -22490 4283
rect -22536 4211 -22490 4249
rect -22536 4177 -22530 4211
rect -22496 4177 -22490 4211
rect -22536 4139 -22490 4177
rect -22536 4105 -22530 4139
rect -22496 4105 -22490 4139
rect -22536 4067 -22490 4105
rect -22536 4033 -22530 4067
rect -22496 4033 -22490 4067
rect -22536 3995 -22490 4033
rect -22536 3961 -22530 3995
rect -22496 3961 -22490 3995
rect -22536 3923 -22490 3961
rect -22536 3889 -22530 3923
rect -22496 3889 -22490 3923
rect -22536 3851 -22490 3889
rect -22536 3817 -22530 3851
rect -22496 3817 -22490 3851
rect -22536 3779 -22490 3817
rect -22536 3745 -22530 3779
rect -22496 3745 -22490 3779
rect -22536 3707 -22490 3745
rect -22536 3673 -22530 3707
rect -22496 3673 -22490 3707
rect -22536 3635 -22490 3673
rect -22536 3601 -22530 3635
rect -22496 3601 -22490 3635
rect -22536 3563 -22490 3601
rect -22536 3529 -22530 3563
rect -22496 3529 -22490 3563
rect -22536 3491 -22490 3529
rect -22536 3457 -22530 3491
rect -22496 3457 -22490 3491
rect -22536 3442 -22490 3457
rect -22440 4427 -22394 4442
rect -22440 4393 -22434 4427
rect -22400 4393 -22394 4427
rect -22440 4355 -22394 4393
rect -22440 4321 -22434 4355
rect -22400 4321 -22394 4355
rect -22440 4283 -22394 4321
rect -22440 4249 -22434 4283
rect -22400 4249 -22394 4283
rect -22440 4211 -22394 4249
rect -22440 4177 -22434 4211
rect -22400 4177 -22394 4211
rect -22440 4139 -22394 4177
rect -22440 4105 -22434 4139
rect -22400 4105 -22394 4139
rect -22440 4067 -22394 4105
rect -22440 4033 -22434 4067
rect -22400 4033 -22394 4067
rect -22440 3995 -22394 4033
rect -22440 3961 -22434 3995
rect -22400 3961 -22394 3995
rect -22440 3923 -22394 3961
rect -22440 3889 -22434 3923
rect -22400 3889 -22394 3923
rect -22440 3851 -22394 3889
rect -22440 3817 -22434 3851
rect -22400 3817 -22394 3851
rect -22440 3779 -22394 3817
rect -22440 3745 -22434 3779
rect -22400 3745 -22394 3779
rect -22440 3707 -22394 3745
rect -22440 3673 -22434 3707
rect -22400 3673 -22394 3707
rect -22440 3635 -22394 3673
rect -22440 3601 -22434 3635
rect -22400 3601 -22394 3635
rect -22440 3563 -22394 3601
rect -22440 3529 -22434 3563
rect -22400 3529 -22394 3563
rect -22440 3491 -22394 3529
rect -22440 3457 -22434 3491
rect -22400 3457 -22394 3491
rect -22440 3442 -22394 3457
rect -22344 4427 -22298 4442
rect -22344 4393 -22338 4427
rect -22304 4393 -22298 4427
rect -22344 4355 -22298 4393
rect -22344 4321 -22338 4355
rect -22304 4321 -22298 4355
rect -22344 4283 -22298 4321
rect -22344 4249 -22338 4283
rect -22304 4249 -22298 4283
rect -22344 4211 -22298 4249
rect -22344 4177 -22338 4211
rect -22304 4177 -22298 4211
rect -22344 4139 -22298 4177
rect -22344 4105 -22338 4139
rect -22304 4105 -22298 4139
rect -22344 4067 -22298 4105
rect -22344 4033 -22338 4067
rect -22304 4033 -22298 4067
rect -22344 3995 -22298 4033
rect -22344 3961 -22338 3995
rect -22304 3961 -22298 3995
rect -22344 3923 -22298 3961
rect -22344 3889 -22338 3923
rect -22304 3889 -22298 3923
rect -22344 3851 -22298 3889
rect -22344 3817 -22338 3851
rect -22304 3817 -22298 3851
rect -22344 3779 -22298 3817
rect -22344 3745 -22338 3779
rect -22304 3745 -22298 3779
rect -22344 3707 -22298 3745
rect -22344 3673 -22338 3707
rect -22304 3673 -22298 3707
rect -22344 3635 -22298 3673
rect -22344 3601 -22338 3635
rect -22304 3601 -22298 3635
rect -22344 3563 -22298 3601
rect -22344 3529 -22338 3563
rect -22304 3529 -22298 3563
rect -22344 3491 -22298 3529
rect -22344 3457 -22338 3491
rect -22304 3457 -22298 3491
rect -22344 3442 -22298 3457
rect -22248 4427 -22202 4442
rect -22248 4393 -22242 4427
rect -22208 4393 -22202 4427
rect -22248 4355 -22202 4393
rect -22248 4321 -22242 4355
rect -22208 4321 -22202 4355
rect -22248 4283 -22202 4321
rect -22248 4249 -22242 4283
rect -22208 4249 -22202 4283
rect -22248 4211 -22202 4249
rect -22248 4177 -22242 4211
rect -22208 4177 -22202 4211
rect -22248 4139 -22202 4177
rect -22248 4105 -22242 4139
rect -22208 4105 -22202 4139
rect -22248 4067 -22202 4105
rect -22248 4033 -22242 4067
rect -22208 4033 -22202 4067
rect -22248 3995 -22202 4033
rect -22248 3961 -22242 3995
rect -22208 3961 -22202 3995
rect -22248 3923 -22202 3961
rect -22248 3889 -22242 3923
rect -22208 3889 -22202 3923
rect -22248 3851 -22202 3889
rect -22248 3817 -22242 3851
rect -22208 3817 -22202 3851
rect -22248 3779 -22202 3817
rect -22248 3745 -22242 3779
rect -22208 3745 -22202 3779
rect -22248 3707 -22202 3745
rect -22248 3673 -22242 3707
rect -22208 3673 -22202 3707
rect -22248 3635 -22202 3673
rect -22248 3601 -22242 3635
rect -22208 3601 -22202 3635
rect -22248 3563 -22202 3601
rect -22248 3529 -22242 3563
rect -22208 3529 -22202 3563
rect -22248 3491 -22202 3529
rect -22248 3457 -22242 3491
rect -22208 3457 -22202 3491
rect -22248 3442 -22202 3457
rect -22152 4427 -22106 4442
rect -22152 4393 -22146 4427
rect -22112 4393 -22106 4427
rect -22152 4355 -22106 4393
rect -22152 4321 -22146 4355
rect -22112 4321 -22106 4355
rect -22152 4283 -22106 4321
rect -22152 4249 -22146 4283
rect -22112 4249 -22106 4283
rect -22152 4211 -22106 4249
rect -22152 4177 -22146 4211
rect -22112 4177 -22106 4211
rect -22152 4139 -22106 4177
rect -22152 4105 -22146 4139
rect -22112 4105 -22106 4139
rect -22152 4067 -22106 4105
rect -22152 4033 -22146 4067
rect -22112 4033 -22106 4067
rect -22152 3995 -22106 4033
rect -22152 3961 -22146 3995
rect -22112 3961 -22106 3995
rect -22152 3923 -22106 3961
rect -22152 3889 -22146 3923
rect -22112 3889 -22106 3923
rect -22152 3851 -22106 3889
rect -22152 3817 -22146 3851
rect -22112 3817 -22106 3851
rect -22152 3779 -22106 3817
rect -22152 3745 -22146 3779
rect -22112 3745 -22106 3779
rect -22152 3707 -22106 3745
rect -22152 3673 -22146 3707
rect -22112 3673 -22106 3707
rect -22152 3635 -22106 3673
rect -22152 3601 -22146 3635
rect -22112 3601 -22106 3635
rect -22152 3563 -22106 3601
rect -22152 3529 -22146 3563
rect -22112 3529 -22106 3563
rect -22152 3491 -22106 3529
rect -22152 3457 -22146 3491
rect -22112 3457 -22106 3491
rect -22152 3442 -22106 3457
rect -22056 4427 -22010 4442
rect -22056 4393 -22050 4427
rect -22016 4393 -22010 4427
rect -22056 4355 -22010 4393
rect -22056 4321 -22050 4355
rect -22016 4321 -22010 4355
rect -22056 4283 -22010 4321
rect -22056 4249 -22050 4283
rect -22016 4249 -22010 4283
rect -22056 4211 -22010 4249
rect -22056 4177 -22050 4211
rect -22016 4177 -22010 4211
rect -22056 4139 -22010 4177
rect -22056 4105 -22050 4139
rect -22016 4105 -22010 4139
rect -22056 4067 -22010 4105
rect -22056 4033 -22050 4067
rect -22016 4033 -22010 4067
rect -22056 3995 -22010 4033
rect -22056 3961 -22050 3995
rect -22016 3961 -22010 3995
rect -22056 3923 -22010 3961
rect -22056 3889 -22050 3923
rect -22016 3889 -22010 3923
rect -22056 3851 -22010 3889
rect -22056 3817 -22050 3851
rect -22016 3817 -22010 3851
rect -22056 3779 -22010 3817
rect -22056 3745 -22050 3779
rect -22016 3745 -22010 3779
rect -22056 3707 -22010 3745
rect -22056 3673 -22050 3707
rect -22016 3673 -22010 3707
rect -22056 3635 -22010 3673
rect -22056 3601 -22050 3635
rect -22016 3601 -22010 3635
rect -22056 3563 -22010 3601
rect -22056 3529 -22050 3563
rect -22016 3529 -22010 3563
rect -22056 3491 -22010 3529
rect -22056 3457 -22050 3491
rect -22016 3457 -22010 3491
rect -22056 3442 -22010 3457
rect -21960 4427 -21914 4442
rect -21960 4393 -21954 4427
rect -21920 4393 -21914 4427
rect -21960 4355 -21914 4393
rect -21960 4321 -21954 4355
rect -21920 4321 -21914 4355
rect -21960 4283 -21914 4321
rect -21960 4249 -21954 4283
rect -21920 4249 -21914 4283
rect -21960 4211 -21914 4249
rect -21960 4177 -21954 4211
rect -21920 4177 -21914 4211
rect -21960 4139 -21914 4177
rect -21960 4105 -21954 4139
rect -21920 4105 -21914 4139
rect -21960 4067 -21914 4105
rect -21960 4033 -21954 4067
rect -21920 4033 -21914 4067
rect -21960 3995 -21914 4033
rect -21960 3961 -21954 3995
rect -21920 3961 -21914 3995
rect -21960 3923 -21914 3961
rect -21960 3889 -21954 3923
rect -21920 3889 -21914 3923
rect -21960 3851 -21914 3889
rect -21960 3817 -21954 3851
rect -21920 3817 -21914 3851
rect -21960 3779 -21914 3817
rect -21960 3745 -21954 3779
rect -21920 3745 -21914 3779
rect -21960 3707 -21914 3745
rect -21960 3673 -21954 3707
rect -21920 3673 -21914 3707
rect -21960 3635 -21914 3673
rect -21960 3601 -21954 3635
rect -21920 3601 -21914 3635
rect -21960 3563 -21914 3601
rect -21960 3529 -21954 3563
rect -21920 3529 -21914 3563
rect -21960 3491 -21914 3529
rect -21960 3457 -21954 3491
rect -21920 3457 -21914 3491
rect -21960 3442 -21914 3457
rect -21864 4427 -21818 4442
rect -21864 4393 -21858 4427
rect -21824 4393 -21818 4427
rect -21864 4355 -21818 4393
rect -21864 4321 -21858 4355
rect -21824 4321 -21818 4355
rect -21864 4283 -21818 4321
rect -21864 4249 -21858 4283
rect -21824 4249 -21818 4283
rect -21864 4211 -21818 4249
rect -21864 4177 -21858 4211
rect -21824 4177 -21818 4211
rect -21864 4139 -21818 4177
rect -21864 4105 -21858 4139
rect -21824 4105 -21818 4139
rect -21864 4067 -21818 4105
rect -21864 4033 -21858 4067
rect -21824 4033 -21818 4067
rect -21864 3995 -21818 4033
rect -21864 3961 -21858 3995
rect -21824 3961 -21818 3995
rect -21864 3923 -21818 3961
rect -21864 3889 -21858 3923
rect -21824 3889 -21818 3923
rect -21864 3851 -21818 3889
rect -21864 3817 -21858 3851
rect -21824 3817 -21818 3851
rect -21864 3779 -21818 3817
rect -21864 3745 -21858 3779
rect -21824 3745 -21818 3779
rect -21864 3707 -21818 3745
rect -21864 3673 -21858 3707
rect -21824 3673 -21818 3707
rect -21864 3635 -21818 3673
rect -21864 3601 -21858 3635
rect -21824 3601 -21818 3635
rect -21864 3563 -21818 3601
rect -21864 3529 -21858 3563
rect -21824 3529 -21818 3563
rect -21864 3491 -21818 3529
rect -21864 3457 -21858 3491
rect -21824 3457 -21818 3491
rect -21864 3442 -21818 3457
rect -21768 4427 -21722 4442
rect -21768 4393 -21762 4427
rect -21728 4393 -21722 4427
rect -21768 4355 -21722 4393
rect -21768 4321 -21762 4355
rect -21728 4321 -21722 4355
rect -21768 4283 -21722 4321
rect -21768 4249 -21762 4283
rect -21728 4249 -21722 4283
rect -21768 4211 -21722 4249
rect -21768 4177 -21762 4211
rect -21728 4177 -21722 4211
rect -21768 4139 -21722 4177
rect -21768 4105 -21762 4139
rect -21728 4105 -21722 4139
rect -21768 4067 -21722 4105
rect -21768 4033 -21762 4067
rect -21728 4033 -21722 4067
rect -21768 3995 -21722 4033
rect -21768 3961 -21762 3995
rect -21728 3961 -21722 3995
rect -21768 3923 -21722 3961
rect -21768 3889 -21762 3923
rect -21728 3889 -21722 3923
rect -21768 3851 -21722 3889
rect -21768 3817 -21762 3851
rect -21728 3817 -21722 3851
rect -21768 3779 -21722 3817
rect -21768 3745 -21762 3779
rect -21728 3745 -21722 3779
rect -21768 3707 -21722 3745
rect -21768 3673 -21762 3707
rect -21728 3673 -21722 3707
rect -21768 3635 -21722 3673
rect -21768 3601 -21762 3635
rect -21728 3601 -21722 3635
rect -21768 3563 -21722 3601
rect -21768 3529 -21762 3563
rect -21728 3529 -21722 3563
rect -21768 3491 -21722 3529
rect -21768 3457 -21762 3491
rect -21728 3457 -21722 3491
rect -21768 3442 -21722 3457
rect -21672 4427 -21626 4442
rect -21672 4393 -21666 4427
rect -21632 4393 -21626 4427
rect -21672 4355 -21626 4393
rect -21672 4321 -21666 4355
rect -21632 4321 -21626 4355
rect -21672 4283 -21626 4321
rect -21672 4249 -21666 4283
rect -21632 4249 -21626 4283
rect -21672 4211 -21626 4249
rect -21672 4177 -21666 4211
rect -21632 4177 -21626 4211
rect -21672 4139 -21626 4177
rect -21672 4105 -21666 4139
rect -21632 4105 -21626 4139
rect -21672 4067 -21626 4105
rect -21672 4033 -21666 4067
rect -21632 4033 -21626 4067
rect -21672 3995 -21626 4033
rect -21672 3961 -21666 3995
rect -21632 3961 -21626 3995
rect -21672 3923 -21626 3961
rect -21672 3889 -21666 3923
rect -21632 3889 -21626 3923
rect -21672 3851 -21626 3889
rect -21672 3817 -21666 3851
rect -21632 3817 -21626 3851
rect -21672 3779 -21626 3817
rect -21672 3745 -21666 3779
rect -21632 3745 -21626 3779
rect -21672 3707 -21626 3745
rect -21672 3673 -21666 3707
rect -21632 3673 -21626 3707
rect -21672 3635 -21626 3673
rect -21672 3601 -21666 3635
rect -21632 3601 -21626 3635
rect -21672 3563 -21626 3601
rect -21672 3529 -21666 3563
rect -21632 3529 -21626 3563
rect -21672 3491 -21626 3529
rect -21672 3457 -21666 3491
rect -21632 3457 -21626 3491
rect -21672 3442 -21626 3457
rect -21448 4433 -21402 4448
rect -21448 4399 -21442 4433
rect -21408 4399 -21402 4433
rect -21448 4361 -21402 4399
rect -21448 4327 -21442 4361
rect -21408 4327 -21402 4361
rect -21448 4289 -21402 4327
rect -21448 4255 -21442 4289
rect -21408 4255 -21402 4289
rect -21448 4217 -21402 4255
rect -21448 4183 -21442 4217
rect -21408 4183 -21402 4217
rect -21448 4145 -21402 4183
rect -21448 4111 -21442 4145
rect -21408 4111 -21402 4145
rect -21448 4073 -21402 4111
rect -21448 4039 -21442 4073
rect -21408 4039 -21402 4073
rect -21448 4001 -21402 4039
rect -21448 3967 -21442 4001
rect -21408 3967 -21402 4001
rect -21448 3929 -21402 3967
rect -21448 3895 -21442 3929
rect -21408 3895 -21402 3929
rect -21448 3857 -21402 3895
rect -21448 3823 -21442 3857
rect -21408 3823 -21402 3857
rect -21448 3785 -21402 3823
rect -21448 3751 -21442 3785
rect -21408 3751 -21402 3785
rect -21448 3713 -21402 3751
rect -21448 3679 -21442 3713
rect -21408 3679 -21402 3713
rect -21448 3641 -21402 3679
rect -21448 3607 -21442 3641
rect -21408 3607 -21402 3641
rect -21448 3569 -21402 3607
rect -21448 3535 -21442 3569
rect -21408 3535 -21402 3569
rect -21448 3497 -21402 3535
rect -21448 3463 -21442 3497
rect -21408 3463 -21402 3497
rect -21448 3448 -21402 3463
rect -21352 4433 -21306 4448
rect -21352 4399 -21346 4433
rect -21312 4399 -21306 4433
rect -21352 4361 -21306 4399
rect -21352 4327 -21346 4361
rect -21312 4327 -21306 4361
rect -21352 4289 -21306 4327
rect -21352 4255 -21346 4289
rect -21312 4255 -21306 4289
rect -21352 4217 -21306 4255
rect -21352 4183 -21346 4217
rect -21312 4183 -21306 4217
rect -21352 4145 -21306 4183
rect -21352 4111 -21346 4145
rect -21312 4111 -21306 4145
rect -21352 4073 -21306 4111
rect -21352 4039 -21346 4073
rect -21312 4039 -21306 4073
rect -21352 4001 -21306 4039
rect -21352 3967 -21346 4001
rect -21312 3967 -21306 4001
rect -21352 3929 -21306 3967
rect -21352 3895 -21346 3929
rect -21312 3895 -21306 3929
rect -21352 3857 -21306 3895
rect -21352 3823 -21346 3857
rect -21312 3823 -21306 3857
rect -21352 3785 -21306 3823
rect -21352 3751 -21346 3785
rect -21312 3751 -21306 3785
rect -21352 3713 -21306 3751
rect -21352 3679 -21346 3713
rect -21312 3679 -21306 3713
rect -21352 3641 -21306 3679
rect -21352 3607 -21346 3641
rect -21312 3607 -21306 3641
rect -21352 3569 -21306 3607
rect -21352 3535 -21346 3569
rect -21312 3535 -21306 3569
rect -21352 3497 -21306 3535
rect -21352 3463 -21346 3497
rect -21312 3463 -21306 3497
rect -21352 3448 -21306 3463
rect -21256 4433 -21210 4448
rect -21256 4399 -21250 4433
rect -21216 4399 -21210 4433
rect -21256 4361 -21210 4399
rect -21256 4327 -21250 4361
rect -21216 4327 -21210 4361
rect -21256 4289 -21210 4327
rect -21256 4255 -21250 4289
rect -21216 4255 -21210 4289
rect -21256 4217 -21210 4255
rect -21256 4183 -21250 4217
rect -21216 4183 -21210 4217
rect -21256 4145 -21210 4183
rect -21256 4111 -21250 4145
rect -21216 4111 -21210 4145
rect -21256 4073 -21210 4111
rect -21256 4039 -21250 4073
rect -21216 4039 -21210 4073
rect -21256 4001 -21210 4039
rect -21256 3967 -21250 4001
rect -21216 3967 -21210 4001
rect -21256 3929 -21210 3967
rect -21256 3895 -21250 3929
rect -21216 3895 -21210 3929
rect -21256 3857 -21210 3895
rect -21256 3823 -21250 3857
rect -21216 3823 -21210 3857
rect -21256 3785 -21210 3823
rect -21256 3751 -21250 3785
rect -21216 3751 -21210 3785
rect -21256 3713 -21210 3751
rect -21256 3679 -21250 3713
rect -21216 3679 -21210 3713
rect -21256 3641 -21210 3679
rect -21256 3607 -21250 3641
rect -21216 3607 -21210 3641
rect -21256 3569 -21210 3607
rect -21256 3535 -21250 3569
rect -21216 3535 -21210 3569
rect -21256 3497 -21210 3535
rect -21256 3463 -21250 3497
rect -21216 3463 -21210 3497
rect -21256 3448 -21210 3463
rect -21160 4433 -21114 4448
rect -21160 4399 -21154 4433
rect -21120 4399 -21114 4433
rect -21160 4361 -21114 4399
rect -21160 4327 -21154 4361
rect -21120 4327 -21114 4361
rect -21160 4289 -21114 4327
rect -21160 4255 -21154 4289
rect -21120 4255 -21114 4289
rect -21160 4217 -21114 4255
rect -21160 4183 -21154 4217
rect -21120 4183 -21114 4217
rect -21160 4145 -21114 4183
rect -21160 4111 -21154 4145
rect -21120 4111 -21114 4145
rect -21160 4073 -21114 4111
rect -21160 4039 -21154 4073
rect -21120 4039 -21114 4073
rect -21160 4001 -21114 4039
rect -21160 3967 -21154 4001
rect -21120 3967 -21114 4001
rect -21160 3929 -21114 3967
rect -21160 3895 -21154 3929
rect -21120 3895 -21114 3929
rect -21160 3857 -21114 3895
rect -21160 3823 -21154 3857
rect -21120 3823 -21114 3857
rect -21160 3785 -21114 3823
rect -21160 3751 -21154 3785
rect -21120 3751 -21114 3785
rect -21160 3713 -21114 3751
rect -21160 3679 -21154 3713
rect -21120 3679 -21114 3713
rect -21160 3641 -21114 3679
rect -21160 3607 -21154 3641
rect -21120 3607 -21114 3641
rect -21160 3569 -21114 3607
rect -21160 3535 -21154 3569
rect -21120 3535 -21114 3569
rect -21160 3497 -21114 3535
rect -21160 3463 -21154 3497
rect -21120 3463 -21114 3497
rect -21160 3448 -21114 3463
rect -21064 4433 -21018 4448
rect -21064 4399 -21058 4433
rect -21024 4399 -21018 4433
rect -21064 4361 -21018 4399
rect -21064 4327 -21058 4361
rect -21024 4327 -21018 4361
rect -21064 4289 -21018 4327
rect -21064 4255 -21058 4289
rect -21024 4255 -21018 4289
rect -21064 4217 -21018 4255
rect -21064 4183 -21058 4217
rect -21024 4183 -21018 4217
rect -21064 4145 -21018 4183
rect -21064 4111 -21058 4145
rect -21024 4111 -21018 4145
rect -21064 4073 -21018 4111
rect -21064 4039 -21058 4073
rect -21024 4039 -21018 4073
rect -21064 4001 -21018 4039
rect -21064 3967 -21058 4001
rect -21024 3967 -21018 4001
rect -21064 3929 -21018 3967
rect -21064 3895 -21058 3929
rect -21024 3895 -21018 3929
rect -21064 3857 -21018 3895
rect -21064 3823 -21058 3857
rect -21024 3823 -21018 3857
rect -21064 3785 -21018 3823
rect -21064 3751 -21058 3785
rect -21024 3751 -21018 3785
rect -21064 3713 -21018 3751
rect -21064 3679 -21058 3713
rect -21024 3679 -21018 3713
rect -21064 3641 -21018 3679
rect -21064 3607 -21058 3641
rect -21024 3607 -21018 3641
rect -21064 3569 -21018 3607
rect -21064 3535 -21058 3569
rect -21024 3535 -21018 3569
rect -21064 3497 -21018 3535
rect -21064 3463 -21058 3497
rect -21024 3463 -21018 3497
rect -21064 3448 -21018 3463
rect -20968 4433 -20922 4448
rect -20968 4399 -20962 4433
rect -20928 4399 -20922 4433
rect -20968 4361 -20922 4399
rect -20968 4327 -20962 4361
rect -20928 4327 -20922 4361
rect -20968 4289 -20922 4327
rect -20968 4255 -20962 4289
rect -20928 4255 -20922 4289
rect -20968 4217 -20922 4255
rect -20968 4183 -20962 4217
rect -20928 4183 -20922 4217
rect -20968 4145 -20922 4183
rect -20968 4111 -20962 4145
rect -20928 4111 -20922 4145
rect -20968 4073 -20922 4111
rect -20968 4039 -20962 4073
rect -20928 4039 -20922 4073
rect -20968 4001 -20922 4039
rect -20968 3967 -20962 4001
rect -20928 3967 -20922 4001
rect -20968 3929 -20922 3967
rect -20968 3895 -20962 3929
rect -20928 3895 -20922 3929
rect -20968 3857 -20922 3895
rect -20968 3823 -20962 3857
rect -20928 3823 -20922 3857
rect -20968 3785 -20922 3823
rect -20968 3751 -20962 3785
rect -20928 3751 -20922 3785
rect -20968 3713 -20922 3751
rect -20968 3679 -20962 3713
rect -20928 3679 -20922 3713
rect -20968 3641 -20922 3679
rect -20968 3607 -20962 3641
rect -20928 3607 -20922 3641
rect -20968 3569 -20922 3607
rect -20968 3535 -20962 3569
rect -20928 3535 -20922 3569
rect -20968 3497 -20922 3535
rect -20968 3463 -20962 3497
rect -20928 3463 -20922 3497
rect -20968 3448 -20922 3463
rect -20872 4433 -20826 4448
rect -20872 4399 -20866 4433
rect -20832 4399 -20826 4433
rect -20872 4361 -20826 4399
rect -20872 4327 -20866 4361
rect -20832 4327 -20826 4361
rect -20872 4289 -20826 4327
rect -20872 4255 -20866 4289
rect -20832 4255 -20826 4289
rect -20872 4217 -20826 4255
rect -20872 4183 -20866 4217
rect -20832 4183 -20826 4217
rect -20872 4145 -20826 4183
rect -20872 4111 -20866 4145
rect -20832 4111 -20826 4145
rect -20872 4073 -20826 4111
rect -20872 4039 -20866 4073
rect -20832 4039 -20826 4073
rect -20872 4001 -20826 4039
rect -20872 3967 -20866 4001
rect -20832 3967 -20826 4001
rect -20872 3929 -20826 3967
rect -20872 3895 -20866 3929
rect -20832 3895 -20826 3929
rect -20872 3857 -20826 3895
rect -20872 3823 -20866 3857
rect -20832 3823 -20826 3857
rect -20872 3785 -20826 3823
rect -20872 3751 -20866 3785
rect -20832 3751 -20826 3785
rect -20872 3713 -20826 3751
rect -20872 3679 -20866 3713
rect -20832 3679 -20826 3713
rect -20872 3641 -20826 3679
rect -20872 3607 -20866 3641
rect -20832 3607 -20826 3641
rect -20872 3569 -20826 3607
rect -20872 3535 -20866 3569
rect -20832 3535 -20826 3569
rect -20872 3497 -20826 3535
rect -20872 3463 -20866 3497
rect -20832 3463 -20826 3497
rect -20872 3448 -20826 3463
rect -20776 4433 -20730 4448
rect -20776 4399 -20770 4433
rect -20736 4399 -20730 4433
rect -20776 4361 -20730 4399
rect -20776 4327 -20770 4361
rect -20736 4327 -20730 4361
rect -20776 4289 -20730 4327
rect -20776 4255 -20770 4289
rect -20736 4255 -20730 4289
rect -20776 4217 -20730 4255
rect -20776 4183 -20770 4217
rect -20736 4183 -20730 4217
rect -20776 4145 -20730 4183
rect -20776 4111 -20770 4145
rect -20736 4111 -20730 4145
rect -20776 4073 -20730 4111
rect -20776 4039 -20770 4073
rect -20736 4039 -20730 4073
rect -20776 4001 -20730 4039
rect -20776 3967 -20770 4001
rect -20736 3967 -20730 4001
rect -20776 3929 -20730 3967
rect -20776 3895 -20770 3929
rect -20736 3895 -20730 3929
rect -20776 3857 -20730 3895
rect -20776 3823 -20770 3857
rect -20736 3823 -20730 3857
rect -20776 3785 -20730 3823
rect -20776 3751 -20770 3785
rect -20736 3751 -20730 3785
rect -20776 3713 -20730 3751
rect -20776 3679 -20770 3713
rect -20736 3679 -20730 3713
rect -20776 3641 -20730 3679
rect -20776 3607 -20770 3641
rect -20736 3607 -20730 3641
rect -20776 3569 -20730 3607
rect -20776 3535 -20770 3569
rect -20736 3535 -20730 3569
rect -20776 3497 -20730 3535
rect -20776 3463 -20770 3497
rect -20736 3463 -20730 3497
rect -20776 3448 -20730 3463
rect -20680 4433 -20634 4448
rect -20680 4399 -20674 4433
rect -20640 4399 -20634 4433
rect -20680 4361 -20634 4399
rect -20680 4327 -20674 4361
rect -20640 4327 -20634 4361
rect -20680 4289 -20634 4327
rect -20680 4255 -20674 4289
rect -20640 4255 -20634 4289
rect -20680 4217 -20634 4255
rect -20680 4183 -20674 4217
rect -20640 4183 -20634 4217
rect -20680 4145 -20634 4183
rect -20680 4111 -20674 4145
rect -20640 4111 -20634 4145
rect -20680 4073 -20634 4111
rect -20680 4039 -20674 4073
rect -20640 4039 -20634 4073
rect -20680 4001 -20634 4039
rect -20680 3967 -20674 4001
rect -20640 3967 -20634 4001
rect -20680 3929 -20634 3967
rect -20680 3895 -20674 3929
rect -20640 3895 -20634 3929
rect -20680 3857 -20634 3895
rect -20680 3823 -20674 3857
rect -20640 3823 -20634 3857
rect -20680 3785 -20634 3823
rect -20680 3751 -20674 3785
rect -20640 3751 -20634 3785
rect -20680 3713 -20634 3751
rect -20680 3679 -20674 3713
rect -20640 3679 -20634 3713
rect -20680 3641 -20634 3679
rect -20680 3607 -20674 3641
rect -20640 3607 -20634 3641
rect -20680 3569 -20634 3607
rect -20680 3535 -20674 3569
rect -20640 3535 -20634 3569
rect -20680 3497 -20634 3535
rect -20680 3463 -20674 3497
rect -20640 3463 -20634 3497
rect -20680 3448 -20634 3463
rect -20584 4433 -20538 4448
rect -20584 4399 -20578 4433
rect -20544 4399 -20538 4433
rect -20584 4361 -20538 4399
rect -20584 4327 -20578 4361
rect -20544 4327 -20538 4361
rect -20584 4289 -20538 4327
rect -20584 4255 -20578 4289
rect -20544 4255 -20538 4289
rect -20584 4217 -20538 4255
rect -20584 4183 -20578 4217
rect -20544 4183 -20538 4217
rect -20584 4145 -20538 4183
rect -20584 4111 -20578 4145
rect -20544 4111 -20538 4145
rect -20584 4073 -20538 4111
rect -20584 4039 -20578 4073
rect -20544 4039 -20538 4073
rect -20584 4001 -20538 4039
rect -20584 3967 -20578 4001
rect -20544 3967 -20538 4001
rect -20584 3929 -20538 3967
rect -20584 3895 -20578 3929
rect -20544 3895 -20538 3929
rect -20584 3857 -20538 3895
rect -20584 3823 -20578 3857
rect -20544 3823 -20538 3857
rect -20584 3785 -20538 3823
rect -20584 3751 -20578 3785
rect -20544 3751 -20538 3785
rect -20584 3713 -20538 3751
rect -20584 3679 -20578 3713
rect -20544 3679 -20538 3713
rect -20584 3641 -20538 3679
rect -20584 3607 -20578 3641
rect -20544 3607 -20538 3641
rect -20584 3569 -20538 3607
rect -20584 3535 -20578 3569
rect -20544 3535 -20538 3569
rect -20584 3497 -20538 3535
rect -20584 3463 -20578 3497
rect -20544 3463 -20538 3497
rect -20584 3448 -20538 3463
rect -20488 4433 -20442 4448
rect -20488 4399 -20482 4433
rect -20448 4399 -20442 4433
rect -20488 4361 -20442 4399
rect -20488 4327 -20482 4361
rect -20448 4327 -20442 4361
rect -20488 4289 -20442 4327
rect -20488 4255 -20482 4289
rect -20448 4255 -20442 4289
rect -20488 4217 -20442 4255
rect -20488 4183 -20482 4217
rect -20448 4183 -20442 4217
rect -20488 4145 -20442 4183
rect -20488 4111 -20482 4145
rect -20448 4111 -20442 4145
rect -20488 4073 -20442 4111
rect -20488 4039 -20482 4073
rect -20448 4039 -20442 4073
rect -20488 4001 -20442 4039
rect -20488 3967 -20482 4001
rect -20448 3967 -20442 4001
rect -20488 3929 -20442 3967
rect -20488 3895 -20482 3929
rect -20448 3895 -20442 3929
rect -20488 3857 -20442 3895
rect -20488 3823 -20482 3857
rect -20448 3823 -20442 3857
rect -20488 3785 -20442 3823
rect -20488 3751 -20482 3785
rect -20448 3751 -20442 3785
rect -20488 3713 -20442 3751
rect -20488 3679 -20482 3713
rect -20448 3679 -20442 3713
rect -20488 3641 -20442 3679
rect -20488 3607 -20482 3641
rect -20448 3607 -20442 3641
rect -20488 3569 -20442 3607
rect -20488 3535 -20482 3569
rect -20448 3535 -20442 3569
rect -20488 3497 -20442 3535
rect -20488 3463 -20482 3497
rect -20448 3463 -20442 3497
rect -20488 3448 -20442 3463
rect -20392 4433 -20346 4448
rect -20392 4399 -20386 4433
rect -20352 4399 -20346 4433
rect -20392 4361 -20346 4399
rect -20392 4327 -20386 4361
rect -20352 4327 -20346 4361
rect -20392 4289 -20346 4327
rect -20392 4255 -20386 4289
rect -20352 4255 -20346 4289
rect -20392 4217 -20346 4255
rect -20392 4183 -20386 4217
rect -20352 4183 -20346 4217
rect -20392 4145 -20346 4183
rect -20392 4111 -20386 4145
rect -20352 4111 -20346 4145
rect -20392 4073 -20346 4111
rect -20392 4039 -20386 4073
rect -20352 4039 -20346 4073
rect -20392 4001 -20346 4039
rect -20392 3967 -20386 4001
rect -20352 3967 -20346 4001
rect -20392 3929 -20346 3967
rect -20392 3895 -20386 3929
rect -20352 3895 -20346 3929
rect -20392 3857 -20346 3895
rect -20392 3823 -20386 3857
rect -20352 3823 -20346 3857
rect -20392 3785 -20346 3823
rect -20392 3751 -20386 3785
rect -20352 3751 -20346 3785
rect -20392 3713 -20346 3751
rect -20392 3679 -20386 3713
rect -20352 3679 -20346 3713
rect -20392 3641 -20346 3679
rect -20392 3607 -20386 3641
rect -20352 3607 -20346 3641
rect -20392 3569 -20346 3607
rect -20392 3535 -20386 3569
rect -20352 3535 -20346 3569
rect -20392 3497 -20346 3535
rect -20392 3463 -20386 3497
rect -20352 3463 -20346 3497
rect -20392 3448 -20346 3463
rect -20296 4433 -20250 4448
rect -20296 4399 -20290 4433
rect -20256 4399 -20250 4433
rect -20296 4361 -20250 4399
rect -20296 4327 -20290 4361
rect -20256 4327 -20250 4361
rect -20296 4289 -20250 4327
rect -20296 4255 -20290 4289
rect -20256 4255 -20250 4289
rect -20296 4217 -20250 4255
rect -20296 4183 -20290 4217
rect -20256 4183 -20250 4217
rect -20296 4145 -20250 4183
rect -20296 4111 -20290 4145
rect -20256 4111 -20250 4145
rect -20296 4073 -20250 4111
rect -20296 4039 -20290 4073
rect -20256 4039 -20250 4073
rect -20296 4001 -20250 4039
rect -20296 3967 -20290 4001
rect -20256 3967 -20250 4001
rect -20296 3929 -20250 3967
rect -20296 3895 -20290 3929
rect -20256 3895 -20250 3929
rect -20296 3857 -20250 3895
rect -20296 3823 -20290 3857
rect -20256 3823 -20250 3857
rect -20296 3785 -20250 3823
rect -20296 3751 -20290 3785
rect -20256 3751 -20250 3785
rect -20296 3713 -20250 3751
rect -20296 3679 -20290 3713
rect -20256 3679 -20250 3713
rect -20296 3641 -20250 3679
rect -20296 3607 -20290 3641
rect -20256 3607 -20250 3641
rect -20296 3569 -20250 3607
rect -20296 3535 -20290 3569
rect -20256 3535 -20250 3569
rect -20296 3497 -20250 3535
rect -20296 3463 -20290 3497
rect -20256 3463 -20250 3497
rect -20296 3448 -20250 3463
rect -20200 4433 -20154 4448
rect -20200 4399 -20194 4433
rect -20160 4399 -20154 4433
rect -20200 4361 -20154 4399
rect -20200 4327 -20194 4361
rect -20160 4327 -20154 4361
rect -20200 4289 -20154 4327
rect -20200 4255 -20194 4289
rect -20160 4255 -20154 4289
rect -20200 4217 -20154 4255
rect -20200 4183 -20194 4217
rect -20160 4183 -20154 4217
rect -20200 4145 -20154 4183
rect -20200 4111 -20194 4145
rect -20160 4111 -20154 4145
rect -20200 4073 -20154 4111
rect -20200 4039 -20194 4073
rect -20160 4039 -20154 4073
rect -20200 4001 -20154 4039
rect -20200 3967 -20194 4001
rect -20160 3967 -20154 4001
rect -20200 3929 -20154 3967
rect -20200 3895 -20194 3929
rect -20160 3895 -20154 3929
rect -20200 3857 -20154 3895
rect -20200 3823 -20194 3857
rect -20160 3823 -20154 3857
rect -20200 3785 -20154 3823
rect -20200 3751 -20194 3785
rect -20160 3751 -20154 3785
rect -20200 3713 -20154 3751
rect -20200 3679 -20194 3713
rect -20160 3679 -20154 3713
rect -20200 3641 -20154 3679
rect -20200 3607 -20194 3641
rect -20160 3607 -20154 3641
rect -20200 3569 -20154 3607
rect -20200 3535 -20194 3569
rect -20160 3535 -20154 3569
rect -20200 3497 -20154 3535
rect -20200 3463 -20194 3497
rect -20160 3463 -20154 3497
rect -20200 3448 -20154 3463
rect -20104 4433 -20058 4448
rect -20104 4399 -20098 4433
rect -20064 4399 -20058 4433
rect -20104 4361 -20058 4399
rect -20104 4327 -20098 4361
rect -20064 4327 -20058 4361
rect -20104 4289 -20058 4327
rect -20104 4255 -20098 4289
rect -20064 4255 -20058 4289
rect -20104 4217 -20058 4255
rect -20104 4183 -20098 4217
rect -20064 4183 -20058 4217
rect -20104 4145 -20058 4183
rect -20104 4111 -20098 4145
rect -20064 4111 -20058 4145
rect -20104 4073 -20058 4111
rect -20104 4039 -20098 4073
rect -20064 4039 -20058 4073
rect -20104 4001 -20058 4039
rect -20104 3967 -20098 4001
rect -20064 3967 -20058 4001
rect -20104 3929 -20058 3967
rect -20104 3895 -20098 3929
rect -20064 3895 -20058 3929
rect -20104 3857 -20058 3895
rect -20104 3823 -20098 3857
rect -20064 3823 -20058 3857
rect -20104 3785 -20058 3823
rect -20104 3751 -20098 3785
rect -20064 3751 -20058 3785
rect -20104 3713 -20058 3751
rect -20104 3679 -20098 3713
rect -20064 3679 -20058 3713
rect -20104 3641 -20058 3679
rect -20104 3607 -20098 3641
rect -20064 3607 -20058 3641
rect -20104 3569 -20058 3607
rect -20104 3535 -20098 3569
rect -20064 3535 -20058 3569
rect -20104 3497 -20058 3535
rect -20104 3463 -20098 3497
rect -20064 3463 -20058 3497
rect -20104 3448 -20058 3463
rect -20008 4433 -19962 4448
rect -20008 4399 -20002 4433
rect -19968 4399 -19962 4433
rect -20008 4361 -19962 4399
rect -20008 4327 -20002 4361
rect -19968 4327 -19962 4361
rect -20008 4289 -19962 4327
rect -20008 4255 -20002 4289
rect -19968 4255 -19962 4289
rect -20008 4217 -19962 4255
rect -20008 4183 -20002 4217
rect -19968 4183 -19962 4217
rect -20008 4145 -19962 4183
rect -20008 4111 -20002 4145
rect -19968 4111 -19962 4145
rect -20008 4073 -19962 4111
rect -20008 4039 -20002 4073
rect -19968 4039 -19962 4073
rect -20008 4001 -19962 4039
rect -20008 3967 -20002 4001
rect -19968 3967 -19962 4001
rect -20008 3929 -19962 3967
rect -20008 3895 -20002 3929
rect -19968 3895 -19962 3929
rect -20008 3857 -19962 3895
rect -20008 3823 -20002 3857
rect -19968 3823 -19962 3857
rect -20008 3785 -19962 3823
rect -20008 3751 -20002 3785
rect -19968 3751 -19962 3785
rect -20008 3713 -19962 3751
rect -20008 3679 -20002 3713
rect -19968 3679 -19962 3713
rect -20008 3641 -19962 3679
rect -20008 3607 -20002 3641
rect -19968 3607 -19962 3641
rect -20008 3569 -19962 3607
rect -20008 3535 -20002 3569
rect -19968 3535 -19962 3569
rect -20008 3497 -19962 3535
rect -20008 3463 -20002 3497
rect -19968 3463 -19962 3497
rect -20008 3448 -19962 3463
rect -19764 4439 -19718 4454
rect -19764 4405 -19758 4439
rect -19724 4405 -19718 4439
rect -19764 4367 -19718 4405
rect -19764 4333 -19758 4367
rect -19724 4333 -19718 4367
rect -19764 4295 -19718 4333
rect -19764 4261 -19758 4295
rect -19724 4261 -19718 4295
rect -19764 4223 -19718 4261
rect -19764 4189 -19758 4223
rect -19724 4189 -19718 4223
rect -19764 4151 -19718 4189
rect -19764 4117 -19758 4151
rect -19724 4117 -19718 4151
rect -19764 4079 -19718 4117
rect -19764 4045 -19758 4079
rect -19724 4045 -19718 4079
rect -19764 4007 -19718 4045
rect -19764 3973 -19758 4007
rect -19724 3973 -19718 4007
rect -19764 3935 -19718 3973
rect -19764 3901 -19758 3935
rect -19724 3901 -19718 3935
rect -19764 3863 -19718 3901
rect -19764 3829 -19758 3863
rect -19724 3829 -19718 3863
rect -19764 3791 -19718 3829
rect -19764 3757 -19758 3791
rect -19724 3757 -19718 3791
rect -19764 3719 -19718 3757
rect -19764 3685 -19758 3719
rect -19724 3685 -19718 3719
rect -19764 3647 -19718 3685
rect -19764 3613 -19758 3647
rect -19724 3613 -19718 3647
rect -19764 3575 -19718 3613
rect -19764 3541 -19758 3575
rect -19724 3541 -19718 3575
rect -19764 3503 -19718 3541
rect -19764 3469 -19758 3503
rect -19724 3469 -19718 3503
rect -19764 3454 -19718 3469
rect -19668 4439 -19622 4454
rect -19668 4405 -19662 4439
rect -19628 4405 -19622 4439
rect -19668 4367 -19622 4405
rect -19668 4333 -19662 4367
rect -19628 4333 -19622 4367
rect -19668 4295 -19622 4333
rect -19668 4261 -19662 4295
rect -19628 4261 -19622 4295
rect -19668 4223 -19622 4261
rect -19668 4189 -19662 4223
rect -19628 4189 -19622 4223
rect -19668 4151 -19622 4189
rect -19668 4117 -19662 4151
rect -19628 4117 -19622 4151
rect -19668 4079 -19622 4117
rect -19668 4045 -19662 4079
rect -19628 4045 -19622 4079
rect -19668 4007 -19622 4045
rect -19668 3973 -19662 4007
rect -19628 3973 -19622 4007
rect -19668 3935 -19622 3973
rect -19668 3901 -19662 3935
rect -19628 3901 -19622 3935
rect -19668 3863 -19622 3901
rect -19668 3829 -19662 3863
rect -19628 3829 -19622 3863
rect -19668 3791 -19622 3829
rect -19668 3757 -19662 3791
rect -19628 3757 -19622 3791
rect -19668 3719 -19622 3757
rect -19668 3685 -19662 3719
rect -19628 3685 -19622 3719
rect -19668 3647 -19622 3685
rect -19668 3613 -19662 3647
rect -19628 3613 -19622 3647
rect -19668 3575 -19622 3613
rect -19668 3541 -19662 3575
rect -19628 3541 -19622 3575
rect -19668 3503 -19622 3541
rect -19668 3469 -19662 3503
rect -19628 3469 -19622 3503
rect -19668 3454 -19622 3469
rect -19572 4439 -19526 4454
rect -19572 4405 -19566 4439
rect -19532 4405 -19526 4439
rect -19572 4367 -19526 4405
rect -19572 4333 -19566 4367
rect -19532 4333 -19526 4367
rect -19572 4295 -19526 4333
rect -19572 4261 -19566 4295
rect -19532 4261 -19526 4295
rect -19572 4223 -19526 4261
rect -19572 4189 -19566 4223
rect -19532 4189 -19526 4223
rect -19572 4151 -19526 4189
rect -19572 4117 -19566 4151
rect -19532 4117 -19526 4151
rect -19572 4079 -19526 4117
rect -19572 4045 -19566 4079
rect -19532 4045 -19526 4079
rect -19572 4007 -19526 4045
rect -19572 3973 -19566 4007
rect -19532 3973 -19526 4007
rect -19572 3935 -19526 3973
rect -19572 3901 -19566 3935
rect -19532 3901 -19526 3935
rect -19572 3863 -19526 3901
rect -19572 3829 -19566 3863
rect -19532 3829 -19526 3863
rect -19572 3791 -19526 3829
rect -19572 3757 -19566 3791
rect -19532 3757 -19526 3791
rect -19572 3719 -19526 3757
rect -19572 3685 -19566 3719
rect -19532 3685 -19526 3719
rect -19572 3647 -19526 3685
rect -19572 3613 -19566 3647
rect -19532 3613 -19526 3647
rect -19572 3575 -19526 3613
rect -19572 3541 -19566 3575
rect -19532 3541 -19526 3575
rect -19572 3503 -19526 3541
rect -19572 3469 -19566 3503
rect -19532 3469 -19526 3503
rect -19572 3454 -19526 3469
rect -19476 4439 -19430 4454
rect -19476 4405 -19470 4439
rect -19436 4405 -19430 4439
rect -19476 4367 -19430 4405
rect -19476 4333 -19470 4367
rect -19436 4333 -19430 4367
rect -19476 4295 -19430 4333
rect -19476 4261 -19470 4295
rect -19436 4261 -19430 4295
rect -19476 4223 -19430 4261
rect -19476 4189 -19470 4223
rect -19436 4189 -19430 4223
rect -19476 4151 -19430 4189
rect -19476 4117 -19470 4151
rect -19436 4117 -19430 4151
rect -19476 4079 -19430 4117
rect -19476 4045 -19470 4079
rect -19436 4045 -19430 4079
rect -19476 4007 -19430 4045
rect -19476 3973 -19470 4007
rect -19436 3973 -19430 4007
rect -19476 3935 -19430 3973
rect -19476 3901 -19470 3935
rect -19436 3901 -19430 3935
rect -19476 3863 -19430 3901
rect -19476 3829 -19470 3863
rect -19436 3829 -19430 3863
rect -19476 3791 -19430 3829
rect -19476 3757 -19470 3791
rect -19436 3757 -19430 3791
rect -19476 3719 -19430 3757
rect -19476 3685 -19470 3719
rect -19436 3685 -19430 3719
rect -19476 3647 -19430 3685
rect -19476 3613 -19470 3647
rect -19436 3613 -19430 3647
rect -19476 3575 -19430 3613
rect -19476 3541 -19470 3575
rect -19436 3541 -19430 3575
rect -19476 3503 -19430 3541
rect -19476 3469 -19470 3503
rect -19436 3469 -19430 3503
rect -19476 3454 -19430 3469
rect -19380 4439 -19334 4454
rect -19380 4405 -19374 4439
rect -19340 4405 -19334 4439
rect -19380 4367 -19334 4405
rect -19380 4333 -19374 4367
rect -19340 4333 -19334 4367
rect -19380 4295 -19334 4333
rect -19380 4261 -19374 4295
rect -19340 4261 -19334 4295
rect -19380 4223 -19334 4261
rect -19380 4189 -19374 4223
rect -19340 4189 -19334 4223
rect -19380 4151 -19334 4189
rect -19380 4117 -19374 4151
rect -19340 4117 -19334 4151
rect -19380 4079 -19334 4117
rect -19380 4045 -19374 4079
rect -19340 4045 -19334 4079
rect -19380 4007 -19334 4045
rect -19380 3973 -19374 4007
rect -19340 3973 -19334 4007
rect -19380 3935 -19334 3973
rect -19380 3901 -19374 3935
rect -19340 3901 -19334 3935
rect -19380 3863 -19334 3901
rect -19380 3829 -19374 3863
rect -19340 3829 -19334 3863
rect -19380 3791 -19334 3829
rect -19380 3757 -19374 3791
rect -19340 3757 -19334 3791
rect -19380 3719 -19334 3757
rect -19380 3685 -19374 3719
rect -19340 3685 -19334 3719
rect -19380 3647 -19334 3685
rect -19380 3613 -19374 3647
rect -19340 3613 -19334 3647
rect -19380 3575 -19334 3613
rect -19380 3541 -19374 3575
rect -19340 3541 -19334 3575
rect -19380 3503 -19334 3541
rect -19380 3469 -19374 3503
rect -19340 3469 -19334 3503
rect -19380 3454 -19334 3469
rect -19284 4439 -19238 4454
rect -19284 4405 -19278 4439
rect -19244 4405 -19238 4439
rect -19284 4367 -19238 4405
rect -19284 4333 -19278 4367
rect -19244 4333 -19238 4367
rect -19284 4295 -19238 4333
rect -19284 4261 -19278 4295
rect -19244 4261 -19238 4295
rect -19284 4223 -19238 4261
rect -19284 4189 -19278 4223
rect -19244 4189 -19238 4223
rect -19284 4151 -19238 4189
rect -19284 4117 -19278 4151
rect -19244 4117 -19238 4151
rect -19284 4079 -19238 4117
rect -19284 4045 -19278 4079
rect -19244 4045 -19238 4079
rect -19284 4007 -19238 4045
rect -19284 3973 -19278 4007
rect -19244 3973 -19238 4007
rect -19284 3935 -19238 3973
rect -19284 3901 -19278 3935
rect -19244 3901 -19238 3935
rect -19284 3863 -19238 3901
rect -19284 3829 -19278 3863
rect -19244 3829 -19238 3863
rect -19284 3791 -19238 3829
rect -19284 3757 -19278 3791
rect -19244 3757 -19238 3791
rect -19284 3719 -19238 3757
rect -19284 3685 -19278 3719
rect -19244 3685 -19238 3719
rect -19284 3647 -19238 3685
rect -19284 3613 -19278 3647
rect -19244 3613 -19238 3647
rect -19284 3575 -19238 3613
rect -19284 3541 -19278 3575
rect -19244 3541 -19238 3575
rect -19284 3503 -19238 3541
rect -19284 3469 -19278 3503
rect -19244 3469 -19238 3503
rect -19284 3454 -19238 3469
rect -19188 4439 -19142 4454
rect -19188 4405 -19182 4439
rect -19148 4405 -19142 4439
rect -19188 4367 -19142 4405
rect -19188 4333 -19182 4367
rect -19148 4333 -19142 4367
rect -19188 4295 -19142 4333
rect -19188 4261 -19182 4295
rect -19148 4261 -19142 4295
rect -19188 4223 -19142 4261
rect -19188 4189 -19182 4223
rect -19148 4189 -19142 4223
rect -19188 4151 -19142 4189
rect -19188 4117 -19182 4151
rect -19148 4117 -19142 4151
rect -19188 4079 -19142 4117
rect -19188 4045 -19182 4079
rect -19148 4045 -19142 4079
rect -19188 4007 -19142 4045
rect -19188 3973 -19182 4007
rect -19148 3973 -19142 4007
rect -19188 3935 -19142 3973
rect -19188 3901 -19182 3935
rect -19148 3901 -19142 3935
rect -19188 3863 -19142 3901
rect -19188 3829 -19182 3863
rect -19148 3829 -19142 3863
rect -19188 3791 -19142 3829
rect -19188 3757 -19182 3791
rect -19148 3757 -19142 3791
rect -19188 3719 -19142 3757
rect -19188 3685 -19182 3719
rect -19148 3685 -19142 3719
rect -19188 3647 -19142 3685
rect -19188 3613 -19182 3647
rect -19148 3613 -19142 3647
rect -19188 3575 -19142 3613
rect -19188 3541 -19182 3575
rect -19148 3541 -19142 3575
rect -19188 3503 -19142 3541
rect -19188 3469 -19182 3503
rect -19148 3469 -19142 3503
rect -19188 3454 -19142 3469
rect -19092 4439 -19046 4454
rect -19092 4405 -19086 4439
rect -19052 4405 -19046 4439
rect -19092 4367 -19046 4405
rect -19092 4333 -19086 4367
rect -19052 4333 -19046 4367
rect -19092 4295 -19046 4333
rect -19092 4261 -19086 4295
rect -19052 4261 -19046 4295
rect -19092 4223 -19046 4261
rect -19092 4189 -19086 4223
rect -19052 4189 -19046 4223
rect -19092 4151 -19046 4189
rect -19092 4117 -19086 4151
rect -19052 4117 -19046 4151
rect -19092 4079 -19046 4117
rect -19092 4045 -19086 4079
rect -19052 4045 -19046 4079
rect -19092 4007 -19046 4045
rect -19092 3973 -19086 4007
rect -19052 3973 -19046 4007
rect -19092 3935 -19046 3973
rect -19092 3901 -19086 3935
rect -19052 3901 -19046 3935
rect -19092 3863 -19046 3901
rect -19092 3829 -19086 3863
rect -19052 3829 -19046 3863
rect -19092 3791 -19046 3829
rect -19092 3757 -19086 3791
rect -19052 3757 -19046 3791
rect -19092 3719 -19046 3757
rect -19092 3685 -19086 3719
rect -19052 3685 -19046 3719
rect -19092 3647 -19046 3685
rect -19092 3613 -19086 3647
rect -19052 3613 -19046 3647
rect -19092 3575 -19046 3613
rect -19092 3541 -19086 3575
rect -19052 3541 -19046 3575
rect -19092 3503 -19046 3541
rect -19092 3469 -19086 3503
rect -19052 3469 -19046 3503
rect -19092 3454 -19046 3469
rect -18996 4439 -18950 4454
rect -18996 4405 -18990 4439
rect -18956 4405 -18950 4439
rect -18996 4367 -18950 4405
rect -18996 4333 -18990 4367
rect -18956 4333 -18950 4367
rect -18996 4295 -18950 4333
rect -18996 4261 -18990 4295
rect -18956 4261 -18950 4295
rect -18996 4223 -18950 4261
rect -18996 4189 -18990 4223
rect -18956 4189 -18950 4223
rect -18996 4151 -18950 4189
rect -18996 4117 -18990 4151
rect -18956 4117 -18950 4151
rect -18996 4079 -18950 4117
rect -18996 4045 -18990 4079
rect -18956 4045 -18950 4079
rect -18996 4007 -18950 4045
rect -18996 3973 -18990 4007
rect -18956 3973 -18950 4007
rect -18996 3935 -18950 3973
rect -18996 3901 -18990 3935
rect -18956 3901 -18950 3935
rect -18996 3863 -18950 3901
rect -18996 3829 -18990 3863
rect -18956 3829 -18950 3863
rect -18996 3791 -18950 3829
rect -18996 3757 -18990 3791
rect -18956 3757 -18950 3791
rect -18996 3719 -18950 3757
rect -18996 3685 -18990 3719
rect -18956 3685 -18950 3719
rect -18996 3647 -18950 3685
rect -18996 3613 -18990 3647
rect -18956 3613 -18950 3647
rect -18996 3575 -18950 3613
rect -18996 3541 -18990 3575
rect -18956 3541 -18950 3575
rect -18996 3503 -18950 3541
rect -18996 3469 -18990 3503
rect -18956 3469 -18950 3503
rect -18996 3454 -18950 3469
rect -18900 4439 -18854 4454
rect -18900 4405 -18894 4439
rect -18860 4405 -18854 4439
rect -18900 4367 -18854 4405
rect -18900 4333 -18894 4367
rect -18860 4333 -18854 4367
rect -18900 4295 -18854 4333
rect -18900 4261 -18894 4295
rect -18860 4261 -18854 4295
rect -18900 4223 -18854 4261
rect -18900 4189 -18894 4223
rect -18860 4189 -18854 4223
rect -18900 4151 -18854 4189
rect -18900 4117 -18894 4151
rect -18860 4117 -18854 4151
rect -18900 4079 -18854 4117
rect -18900 4045 -18894 4079
rect -18860 4045 -18854 4079
rect -18900 4007 -18854 4045
rect -18900 3973 -18894 4007
rect -18860 3973 -18854 4007
rect -18900 3935 -18854 3973
rect -18900 3901 -18894 3935
rect -18860 3901 -18854 3935
rect -18900 3863 -18854 3901
rect -18900 3829 -18894 3863
rect -18860 3829 -18854 3863
rect -18900 3791 -18854 3829
rect -18900 3757 -18894 3791
rect -18860 3757 -18854 3791
rect -18900 3719 -18854 3757
rect -18900 3685 -18894 3719
rect -18860 3685 -18854 3719
rect -18900 3647 -18854 3685
rect -18900 3613 -18894 3647
rect -18860 3613 -18854 3647
rect -18900 3575 -18854 3613
rect -18900 3541 -18894 3575
rect -18860 3541 -18854 3575
rect -18900 3503 -18854 3541
rect -18900 3469 -18894 3503
rect -18860 3469 -18854 3503
rect -18900 3454 -18854 3469
rect -18804 4439 -18758 4454
rect -18804 4405 -18798 4439
rect -18764 4405 -18758 4439
rect -18804 4367 -18758 4405
rect -18804 4333 -18798 4367
rect -18764 4333 -18758 4367
rect -18804 4295 -18758 4333
rect -18804 4261 -18798 4295
rect -18764 4261 -18758 4295
rect -18804 4223 -18758 4261
rect -18804 4189 -18798 4223
rect -18764 4189 -18758 4223
rect -18804 4151 -18758 4189
rect -18804 4117 -18798 4151
rect -18764 4117 -18758 4151
rect -18804 4079 -18758 4117
rect -18804 4045 -18798 4079
rect -18764 4045 -18758 4079
rect -18804 4007 -18758 4045
rect -18804 3973 -18798 4007
rect -18764 3973 -18758 4007
rect -18804 3935 -18758 3973
rect -18804 3901 -18798 3935
rect -18764 3901 -18758 3935
rect -18804 3863 -18758 3901
rect -18804 3829 -18798 3863
rect -18764 3829 -18758 3863
rect -18804 3791 -18758 3829
rect -18804 3757 -18798 3791
rect -18764 3757 -18758 3791
rect -18804 3719 -18758 3757
rect -18804 3685 -18798 3719
rect -18764 3685 -18758 3719
rect -18804 3647 -18758 3685
rect -18804 3613 -18798 3647
rect -18764 3613 -18758 3647
rect -18804 3575 -18758 3613
rect -18804 3541 -18798 3575
rect -18764 3541 -18758 3575
rect -18804 3503 -18758 3541
rect -18804 3469 -18798 3503
rect -18764 3469 -18758 3503
rect -18804 3454 -18758 3469
rect -18596 4441 -18550 4456
rect -18596 4407 -18590 4441
rect -18556 4407 -18550 4441
rect -18596 4369 -18550 4407
rect -18596 4335 -18590 4369
rect -18556 4335 -18550 4369
rect -18596 4297 -18550 4335
rect -18596 4263 -18590 4297
rect -18556 4263 -18550 4297
rect -18596 4225 -18550 4263
rect -18596 4191 -18590 4225
rect -18556 4191 -18550 4225
rect -18596 4153 -18550 4191
rect -18596 4119 -18590 4153
rect -18556 4119 -18550 4153
rect -18596 4081 -18550 4119
rect -18596 4047 -18590 4081
rect -18556 4047 -18550 4081
rect -18596 4009 -18550 4047
rect -18596 3975 -18590 4009
rect -18556 3975 -18550 4009
rect -18596 3937 -18550 3975
rect -18596 3903 -18590 3937
rect -18556 3903 -18550 3937
rect -18596 3865 -18550 3903
rect -18596 3831 -18590 3865
rect -18556 3831 -18550 3865
rect -18596 3793 -18550 3831
rect -18596 3759 -18590 3793
rect -18556 3759 -18550 3793
rect -18596 3721 -18550 3759
rect -18596 3687 -18590 3721
rect -18556 3687 -18550 3721
rect -18596 3649 -18550 3687
rect -18596 3615 -18590 3649
rect -18556 3615 -18550 3649
rect -18596 3577 -18550 3615
rect -18596 3543 -18590 3577
rect -18556 3543 -18550 3577
rect -18596 3505 -18550 3543
rect -18596 3471 -18590 3505
rect -18556 3471 -18550 3505
rect -18596 3456 -18550 3471
rect -18500 4441 -18454 4456
rect -18500 4407 -18494 4441
rect -18460 4407 -18454 4441
rect -18500 4369 -18454 4407
rect -18500 4335 -18494 4369
rect -18460 4335 -18454 4369
rect -18500 4297 -18454 4335
rect -18500 4263 -18494 4297
rect -18460 4263 -18454 4297
rect -18500 4225 -18454 4263
rect -18500 4191 -18494 4225
rect -18460 4191 -18454 4225
rect -18500 4153 -18454 4191
rect -18500 4119 -18494 4153
rect -18460 4119 -18454 4153
rect -18500 4081 -18454 4119
rect -18500 4047 -18494 4081
rect -18460 4047 -18454 4081
rect -18500 4009 -18454 4047
rect -18500 3975 -18494 4009
rect -18460 3975 -18454 4009
rect -18500 3937 -18454 3975
rect -18500 3903 -18494 3937
rect -18460 3903 -18454 3937
rect -18500 3865 -18454 3903
rect -18500 3831 -18494 3865
rect -18460 3831 -18454 3865
rect -18500 3793 -18454 3831
rect -18500 3759 -18494 3793
rect -18460 3759 -18454 3793
rect -18500 3721 -18454 3759
rect -18500 3687 -18494 3721
rect -18460 3687 -18454 3721
rect -18500 3649 -18454 3687
rect -18500 3615 -18494 3649
rect -18460 3615 -18454 3649
rect -18500 3577 -18454 3615
rect -18500 3543 -18494 3577
rect -18460 3543 -18454 3577
rect -18500 3505 -18454 3543
rect -18500 3471 -18494 3505
rect -18460 3471 -18454 3505
rect -18500 3456 -18454 3471
rect -18404 4441 -18358 4456
rect -18404 4407 -18398 4441
rect -18364 4407 -18358 4441
rect -18404 4369 -18358 4407
rect -18404 4335 -18398 4369
rect -18364 4335 -18358 4369
rect -18404 4297 -18358 4335
rect -18404 4263 -18398 4297
rect -18364 4263 -18358 4297
rect -18404 4225 -18358 4263
rect -18404 4191 -18398 4225
rect -18364 4191 -18358 4225
rect -18404 4153 -18358 4191
rect -18404 4119 -18398 4153
rect -18364 4119 -18358 4153
rect -18404 4081 -18358 4119
rect -18404 4047 -18398 4081
rect -18364 4047 -18358 4081
rect -18404 4009 -18358 4047
rect -18404 3975 -18398 4009
rect -18364 3975 -18358 4009
rect -18404 3937 -18358 3975
rect -18404 3903 -18398 3937
rect -18364 3903 -18358 3937
rect -18404 3865 -18358 3903
rect -18404 3831 -18398 3865
rect -18364 3831 -18358 3865
rect -18404 3793 -18358 3831
rect -18404 3759 -18398 3793
rect -18364 3759 -18358 3793
rect -18404 3721 -18358 3759
rect -18404 3687 -18398 3721
rect -18364 3687 -18358 3721
rect -18404 3649 -18358 3687
rect -18404 3615 -18398 3649
rect -18364 3615 -18358 3649
rect -18404 3577 -18358 3615
rect -18404 3543 -18398 3577
rect -18364 3543 -18358 3577
rect -18404 3505 -18358 3543
rect -18404 3471 -18398 3505
rect -18364 3471 -18358 3505
rect -18404 3456 -18358 3471
rect -18308 4441 -18262 4456
rect -18308 4407 -18302 4441
rect -18268 4407 -18262 4441
rect -18308 4369 -18262 4407
rect -18308 4335 -18302 4369
rect -18268 4335 -18262 4369
rect -18308 4297 -18262 4335
rect -18308 4263 -18302 4297
rect -18268 4263 -18262 4297
rect -18308 4225 -18262 4263
rect -18308 4191 -18302 4225
rect -18268 4191 -18262 4225
rect -18308 4153 -18262 4191
rect -18308 4119 -18302 4153
rect -18268 4119 -18262 4153
rect -18308 4081 -18262 4119
rect -18308 4047 -18302 4081
rect -18268 4047 -18262 4081
rect -18308 4009 -18262 4047
rect -18308 3975 -18302 4009
rect -18268 3975 -18262 4009
rect -18308 3937 -18262 3975
rect -18308 3903 -18302 3937
rect -18268 3903 -18262 3937
rect -18308 3865 -18262 3903
rect -18308 3831 -18302 3865
rect -18268 3831 -18262 3865
rect -18308 3793 -18262 3831
rect -18308 3759 -18302 3793
rect -18268 3759 -18262 3793
rect -18308 3721 -18262 3759
rect -18308 3687 -18302 3721
rect -18268 3687 -18262 3721
rect -18308 3649 -18262 3687
rect -18308 3615 -18302 3649
rect -18268 3615 -18262 3649
rect -18308 3577 -18262 3615
rect -18308 3543 -18302 3577
rect -18268 3543 -18262 3577
rect -18308 3505 -18262 3543
rect -18308 3471 -18302 3505
rect -18268 3471 -18262 3505
rect -18308 3456 -18262 3471
rect -18212 4441 -18166 4456
rect -18212 4407 -18206 4441
rect -18172 4407 -18166 4441
rect -18212 4369 -18166 4407
rect -18212 4335 -18206 4369
rect -18172 4335 -18166 4369
rect -18212 4297 -18166 4335
rect -18212 4263 -18206 4297
rect -18172 4263 -18166 4297
rect -18212 4225 -18166 4263
rect -18212 4191 -18206 4225
rect -18172 4191 -18166 4225
rect -18212 4153 -18166 4191
rect -18212 4119 -18206 4153
rect -18172 4119 -18166 4153
rect -18212 4081 -18166 4119
rect -18212 4047 -18206 4081
rect -18172 4047 -18166 4081
rect -18212 4009 -18166 4047
rect -18212 3975 -18206 4009
rect -18172 3975 -18166 4009
rect -18212 3937 -18166 3975
rect -18212 3903 -18206 3937
rect -18172 3903 -18166 3937
rect -18212 3865 -18166 3903
rect -18212 3831 -18206 3865
rect -18172 3831 -18166 3865
rect -18212 3793 -18166 3831
rect -18212 3759 -18206 3793
rect -18172 3759 -18166 3793
rect -18212 3721 -18166 3759
rect -18212 3687 -18206 3721
rect -18172 3687 -18166 3721
rect -18212 3649 -18166 3687
rect -18212 3615 -18206 3649
rect -18172 3615 -18166 3649
rect -18212 3577 -18166 3615
rect -18212 3543 -18206 3577
rect -18172 3543 -18166 3577
rect -18212 3505 -18166 3543
rect -18212 3471 -18206 3505
rect -18172 3471 -18166 3505
rect -18212 3456 -18166 3471
rect -18116 4441 -18070 4456
rect -18116 4407 -18110 4441
rect -18076 4407 -18070 4441
rect -18116 4369 -18070 4407
rect -18116 4335 -18110 4369
rect -18076 4335 -18070 4369
rect -18116 4297 -18070 4335
rect -18116 4263 -18110 4297
rect -18076 4263 -18070 4297
rect -18116 4225 -18070 4263
rect -18116 4191 -18110 4225
rect -18076 4191 -18070 4225
rect -18116 4153 -18070 4191
rect -18116 4119 -18110 4153
rect -18076 4119 -18070 4153
rect -18116 4081 -18070 4119
rect -18116 4047 -18110 4081
rect -18076 4047 -18070 4081
rect -18116 4009 -18070 4047
rect -18116 3975 -18110 4009
rect -18076 3975 -18070 4009
rect -18116 3937 -18070 3975
rect -18116 3903 -18110 3937
rect -18076 3903 -18070 3937
rect -18116 3865 -18070 3903
rect -18116 3831 -18110 3865
rect -18076 3831 -18070 3865
rect -18116 3793 -18070 3831
rect -18116 3759 -18110 3793
rect -18076 3759 -18070 3793
rect -18116 3721 -18070 3759
rect -18116 3687 -18110 3721
rect -18076 3687 -18070 3721
rect -18116 3649 -18070 3687
rect -18116 3615 -18110 3649
rect -18076 3615 -18070 3649
rect -18116 3577 -18070 3615
rect -18116 3543 -18110 3577
rect -18076 3543 -18070 3577
rect -18116 3505 -18070 3543
rect -18116 3471 -18110 3505
rect -18076 3471 -18070 3505
rect -18116 3456 -18070 3471
rect -16762 4439 -16716 4454
rect -16762 4405 -16756 4439
rect -16722 4405 -16716 4439
rect -16762 4367 -16716 4405
rect -16762 4333 -16756 4367
rect -16722 4333 -16716 4367
rect -16762 4295 -16716 4333
rect -16762 4261 -16756 4295
rect -16722 4261 -16716 4295
rect -16762 4223 -16716 4261
rect -16762 4189 -16756 4223
rect -16722 4189 -16716 4223
rect -16762 4151 -16716 4189
rect -16762 4117 -16756 4151
rect -16722 4117 -16716 4151
rect -16762 4079 -16716 4117
rect -16762 4045 -16756 4079
rect -16722 4045 -16716 4079
rect -16762 4007 -16716 4045
rect -16762 3973 -16756 4007
rect -16722 3973 -16716 4007
rect -16762 3935 -16716 3973
rect -16762 3901 -16756 3935
rect -16722 3901 -16716 3935
rect -16762 3863 -16716 3901
rect -16762 3829 -16756 3863
rect -16722 3829 -16716 3863
rect -16762 3791 -16716 3829
rect -16762 3757 -16756 3791
rect -16722 3757 -16716 3791
rect -16762 3719 -16716 3757
rect -16762 3685 -16756 3719
rect -16722 3685 -16716 3719
rect -16762 3647 -16716 3685
rect -16762 3613 -16756 3647
rect -16722 3613 -16716 3647
rect -16762 3575 -16716 3613
rect -16762 3541 -16756 3575
rect -16722 3541 -16716 3575
rect -16762 3503 -16716 3541
rect -16762 3469 -16756 3503
rect -16722 3469 -16716 3503
rect -16762 3454 -16716 3469
rect -16666 4439 -16620 4454
rect -16666 4405 -16660 4439
rect -16626 4405 -16620 4439
rect -16666 4367 -16620 4405
rect -16666 4333 -16660 4367
rect -16626 4333 -16620 4367
rect -16666 4295 -16620 4333
rect -16666 4261 -16660 4295
rect -16626 4261 -16620 4295
rect -16666 4223 -16620 4261
rect -16666 4189 -16660 4223
rect -16626 4189 -16620 4223
rect -16666 4151 -16620 4189
rect -16666 4117 -16660 4151
rect -16626 4117 -16620 4151
rect -16666 4079 -16620 4117
rect -16666 4045 -16660 4079
rect -16626 4045 -16620 4079
rect -16666 4007 -16620 4045
rect -16666 3973 -16660 4007
rect -16626 3973 -16620 4007
rect -16666 3935 -16620 3973
rect -16666 3901 -16660 3935
rect -16626 3901 -16620 3935
rect -16666 3863 -16620 3901
rect -16666 3829 -16660 3863
rect -16626 3829 -16620 3863
rect -16666 3791 -16620 3829
rect -16666 3757 -16660 3791
rect -16626 3757 -16620 3791
rect -16666 3719 -16620 3757
rect -16666 3685 -16660 3719
rect -16626 3685 -16620 3719
rect -16666 3647 -16620 3685
rect -16666 3613 -16660 3647
rect -16626 3613 -16620 3647
rect -16666 3575 -16620 3613
rect -16666 3541 -16660 3575
rect -16626 3541 -16620 3575
rect -16666 3503 -16620 3541
rect -16666 3469 -16660 3503
rect -16626 3469 -16620 3503
rect -16666 3454 -16620 3469
rect -16570 4439 -16524 4454
rect -16570 4405 -16564 4439
rect -16530 4405 -16524 4439
rect -16570 4367 -16524 4405
rect -16570 4333 -16564 4367
rect -16530 4333 -16524 4367
rect -16570 4295 -16524 4333
rect -16570 4261 -16564 4295
rect -16530 4261 -16524 4295
rect -16570 4223 -16524 4261
rect -16570 4189 -16564 4223
rect -16530 4189 -16524 4223
rect -16570 4151 -16524 4189
rect -16570 4117 -16564 4151
rect -16530 4117 -16524 4151
rect -16570 4079 -16524 4117
rect -16570 4045 -16564 4079
rect -16530 4045 -16524 4079
rect -16570 4007 -16524 4045
rect -16570 3973 -16564 4007
rect -16530 3973 -16524 4007
rect -16570 3935 -16524 3973
rect -16570 3901 -16564 3935
rect -16530 3901 -16524 3935
rect -16570 3863 -16524 3901
rect -16570 3829 -16564 3863
rect -16530 3829 -16524 3863
rect -16570 3791 -16524 3829
rect -16570 3757 -16564 3791
rect -16530 3757 -16524 3791
rect -16570 3719 -16524 3757
rect -16570 3685 -16564 3719
rect -16530 3685 -16524 3719
rect -16570 3647 -16524 3685
rect -16570 3613 -16564 3647
rect -16530 3613 -16524 3647
rect -16570 3575 -16524 3613
rect -16570 3541 -16564 3575
rect -16530 3541 -16524 3575
rect -16570 3503 -16524 3541
rect -16570 3469 -16564 3503
rect -16530 3469 -16524 3503
rect -16570 3454 -16524 3469
rect -16474 4439 -16428 4454
rect -16474 4405 -16468 4439
rect -16434 4405 -16428 4439
rect -16474 4367 -16428 4405
rect -16474 4333 -16468 4367
rect -16434 4333 -16428 4367
rect -16474 4295 -16428 4333
rect -16474 4261 -16468 4295
rect -16434 4261 -16428 4295
rect -16474 4223 -16428 4261
rect -16474 4189 -16468 4223
rect -16434 4189 -16428 4223
rect -16474 4151 -16428 4189
rect -16474 4117 -16468 4151
rect -16434 4117 -16428 4151
rect -16474 4079 -16428 4117
rect -16474 4045 -16468 4079
rect -16434 4045 -16428 4079
rect -16474 4007 -16428 4045
rect -16474 3973 -16468 4007
rect -16434 3973 -16428 4007
rect -16474 3935 -16428 3973
rect -16474 3901 -16468 3935
rect -16434 3901 -16428 3935
rect -16474 3863 -16428 3901
rect -16474 3829 -16468 3863
rect -16434 3829 -16428 3863
rect -16474 3791 -16428 3829
rect -16474 3757 -16468 3791
rect -16434 3757 -16428 3791
rect -16474 3719 -16428 3757
rect -16474 3685 -16468 3719
rect -16434 3685 -16428 3719
rect -16474 3647 -16428 3685
rect -16474 3613 -16468 3647
rect -16434 3613 -16428 3647
rect -16474 3575 -16428 3613
rect -16474 3541 -16468 3575
rect -16434 3541 -16428 3575
rect -16474 3503 -16428 3541
rect -16474 3469 -16468 3503
rect -16434 3469 -16428 3503
rect -16474 3454 -16428 3469
rect -16378 4439 -16332 4454
rect -16378 4405 -16372 4439
rect -16338 4405 -16332 4439
rect -16378 4367 -16332 4405
rect -16378 4333 -16372 4367
rect -16338 4333 -16332 4367
rect -16378 4295 -16332 4333
rect -16378 4261 -16372 4295
rect -16338 4261 -16332 4295
rect -16378 4223 -16332 4261
rect -16378 4189 -16372 4223
rect -16338 4189 -16332 4223
rect -16378 4151 -16332 4189
rect -16378 4117 -16372 4151
rect -16338 4117 -16332 4151
rect -16378 4079 -16332 4117
rect -16378 4045 -16372 4079
rect -16338 4045 -16332 4079
rect -16378 4007 -16332 4045
rect -16378 3973 -16372 4007
rect -16338 3973 -16332 4007
rect -16378 3935 -16332 3973
rect -16378 3901 -16372 3935
rect -16338 3901 -16332 3935
rect -16378 3863 -16332 3901
rect -16378 3829 -16372 3863
rect -16338 3829 -16332 3863
rect -16378 3791 -16332 3829
rect -16378 3757 -16372 3791
rect -16338 3757 -16332 3791
rect -16378 3719 -16332 3757
rect -16378 3685 -16372 3719
rect -16338 3685 -16332 3719
rect -16378 3647 -16332 3685
rect -16378 3613 -16372 3647
rect -16338 3613 -16332 3647
rect -16378 3575 -16332 3613
rect -16378 3541 -16372 3575
rect -16338 3541 -16332 3575
rect -16378 3503 -16332 3541
rect -16378 3469 -16372 3503
rect -16338 3469 -16332 3503
rect -16378 3454 -16332 3469
rect -16282 4439 -16236 4454
rect -16282 4405 -16276 4439
rect -16242 4405 -16236 4439
rect -16282 4367 -16236 4405
rect -16282 4333 -16276 4367
rect -16242 4333 -16236 4367
rect -16282 4295 -16236 4333
rect -16282 4261 -16276 4295
rect -16242 4261 -16236 4295
rect -16282 4223 -16236 4261
rect -16282 4189 -16276 4223
rect -16242 4189 -16236 4223
rect -16282 4151 -16236 4189
rect -16282 4117 -16276 4151
rect -16242 4117 -16236 4151
rect -16282 4079 -16236 4117
rect -16282 4045 -16276 4079
rect -16242 4045 -16236 4079
rect -16282 4007 -16236 4045
rect -16282 3973 -16276 4007
rect -16242 3973 -16236 4007
rect -16282 3935 -16236 3973
rect -16282 3901 -16276 3935
rect -16242 3901 -16236 3935
rect -16282 3863 -16236 3901
rect -16282 3829 -16276 3863
rect -16242 3829 -16236 3863
rect -16282 3791 -16236 3829
rect -16282 3757 -16276 3791
rect -16242 3757 -16236 3791
rect -16282 3719 -16236 3757
rect -16282 3685 -16276 3719
rect -16242 3685 -16236 3719
rect -16282 3647 -16236 3685
rect -16282 3613 -16276 3647
rect -16242 3613 -16236 3647
rect -16282 3575 -16236 3613
rect -16282 3541 -16276 3575
rect -16242 3541 -16236 3575
rect -16282 3503 -16236 3541
rect -16282 3469 -16276 3503
rect -16242 3469 -16236 3503
rect -16282 3454 -16236 3469
rect -16186 4439 -16140 4454
rect -16186 4405 -16180 4439
rect -16146 4405 -16140 4439
rect -16186 4367 -16140 4405
rect -16186 4333 -16180 4367
rect -16146 4333 -16140 4367
rect -16186 4295 -16140 4333
rect -16186 4261 -16180 4295
rect -16146 4261 -16140 4295
rect -16186 4223 -16140 4261
rect -16186 4189 -16180 4223
rect -16146 4189 -16140 4223
rect -16186 4151 -16140 4189
rect -16186 4117 -16180 4151
rect -16146 4117 -16140 4151
rect -16186 4079 -16140 4117
rect -16186 4045 -16180 4079
rect -16146 4045 -16140 4079
rect -16186 4007 -16140 4045
rect -16186 3973 -16180 4007
rect -16146 3973 -16140 4007
rect -16186 3935 -16140 3973
rect -16186 3901 -16180 3935
rect -16146 3901 -16140 3935
rect -16186 3863 -16140 3901
rect -16186 3829 -16180 3863
rect -16146 3829 -16140 3863
rect -16186 3791 -16140 3829
rect -16186 3757 -16180 3791
rect -16146 3757 -16140 3791
rect -16186 3719 -16140 3757
rect -16186 3685 -16180 3719
rect -16146 3685 -16140 3719
rect -16186 3647 -16140 3685
rect -16186 3613 -16180 3647
rect -16146 3613 -16140 3647
rect -16186 3575 -16140 3613
rect -16186 3541 -16180 3575
rect -16146 3541 -16140 3575
rect -16186 3503 -16140 3541
rect -16186 3469 -16180 3503
rect -16146 3469 -16140 3503
rect -16186 3454 -16140 3469
rect -16090 4439 -16044 4454
rect -16090 4405 -16084 4439
rect -16050 4405 -16044 4439
rect -16090 4367 -16044 4405
rect -16090 4333 -16084 4367
rect -16050 4333 -16044 4367
rect -16090 4295 -16044 4333
rect -16090 4261 -16084 4295
rect -16050 4261 -16044 4295
rect -16090 4223 -16044 4261
rect -16090 4189 -16084 4223
rect -16050 4189 -16044 4223
rect -16090 4151 -16044 4189
rect -16090 4117 -16084 4151
rect -16050 4117 -16044 4151
rect -16090 4079 -16044 4117
rect -16090 4045 -16084 4079
rect -16050 4045 -16044 4079
rect -16090 4007 -16044 4045
rect -16090 3973 -16084 4007
rect -16050 3973 -16044 4007
rect -16090 3935 -16044 3973
rect -16090 3901 -16084 3935
rect -16050 3901 -16044 3935
rect -16090 3863 -16044 3901
rect -16090 3829 -16084 3863
rect -16050 3829 -16044 3863
rect -16090 3791 -16044 3829
rect -16090 3757 -16084 3791
rect -16050 3757 -16044 3791
rect -16090 3719 -16044 3757
rect -16090 3685 -16084 3719
rect -16050 3685 -16044 3719
rect -16090 3647 -16044 3685
rect -16090 3613 -16084 3647
rect -16050 3613 -16044 3647
rect -16090 3575 -16044 3613
rect -16090 3541 -16084 3575
rect -16050 3541 -16044 3575
rect -16090 3503 -16044 3541
rect -16090 3469 -16084 3503
rect -16050 3469 -16044 3503
rect -16090 3454 -16044 3469
rect -15994 4439 -15948 4454
rect -15994 4405 -15988 4439
rect -15954 4405 -15948 4439
rect -15994 4367 -15948 4405
rect -15994 4333 -15988 4367
rect -15954 4333 -15948 4367
rect -15994 4295 -15948 4333
rect -15994 4261 -15988 4295
rect -15954 4261 -15948 4295
rect -15994 4223 -15948 4261
rect -15994 4189 -15988 4223
rect -15954 4189 -15948 4223
rect -15994 4151 -15948 4189
rect -15994 4117 -15988 4151
rect -15954 4117 -15948 4151
rect -15994 4079 -15948 4117
rect -15994 4045 -15988 4079
rect -15954 4045 -15948 4079
rect -15994 4007 -15948 4045
rect -15994 3973 -15988 4007
rect -15954 3973 -15948 4007
rect -15994 3935 -15948 3973
rect -15994 3901 -15988 3935
rect -15954 3901 -15948 3935
rect -15994 3863 -15948 3901
rect -15994 3829 -15988 3863
rect -15954 3829 -15948 3863
rect -15994 3791 -15948 3829
rect -15994 3757 -15988 3791
rect -15954 3757 -15948 3791
rect -15994 3719 -15948 3757
rect -15994 3685 -15988 3719
rect -15954 3685 -15948 3719
rect -15994 3647 -15948 3685
rect -15994 3613 -15988 3647
rect -15954 3613 -15948 3647
rect -15994 3575 -15948 3613
rect -15994 3541 -15988 3575
rect -15954 3541 -15948 3575
rect -15994 3503 -15948 3541
rect -15994 3469 -15988 3503
rect -15954 3469 -15948 3503
rect -15994 3454 -15948 3469
rect -15898 4439 -15852 4454
rect -15898 4405 -15892 4439
rect -15858 4405 -15852 4439
rect -15898 4367 -15852 4405
rect -15898 4333 -15892 4367
rect -15858 4333 -15852 4367
rect -15898 4295 -15852 4333
rect -15898 4261 -15892 4295
rect -15858 4261 -15852 4295
rect -15898 4223 -15852 4261
rect -15898 4189 -15892 4223
rect -15858 4189 -15852 4223
rect -15898 4151 -15852 4189
rect -15898 4117 -15892 4151
rect -15858 4117 -15852 4151
rect -15898 4079 -15852 4117
rect -15898 4045 -15892 4079
rect -15858 4045 -15852 4079
rect -15898 4007 -15852 4045
rect -15898 3973 -15892 4007
rect -15858 3973 -15852 4007
rect -15898 3935 -15852 3973
rect -15898 3901 -15892 3935
rect -15858 3901 -15852 3935
rect -15898 3863 -15852 3901
rect -15898 3829 -15892 3863
rect -15858 3829 -15852 3863
rect -15898 3791 -15852 3829
rect -15898 3757 -15892 3791
rect -15858 3757 -15852 3791
rect -15898 3719 -15852 3757
rect -15898 3685 -15892 3719
rect -15858 3685 -15852 3719
rect -15898 3647 -15852 3685
rect -15898 3613 -15892 3647
rect -15858 3613 -15852 3647
rect -15898 3575 -15852 3613
rect -15898 3541 -15892 3575
rect -15858 3541 -15852 3575
rect -15898 3503 -15852 3541
rect -15898 3469 -15892 3503
rect -15858 3469 -15852 3503
rect -15898 3454 -15852 3469
rect -15802 4439 -15756 4454
rect -15802 4405 -15796 4439
rect -15762 4405 -15756 4439
rect -15802 4367 -15756 4405
rect -15802 4333 -15796 4367
rect -15762 4333 -15756 4367
rect -15802 4295 -15756 4333
rect -15802 4261 -15796 4295
rect -15762 4261 -15756 4295
rect -15802 4223 -15756 4261
rect -15802 4189 -15796 4223
rect -15762 4189 -15756 4223
rect -15802 4151 -15756 4189
rect -15802 4117 -15796 4151
rect -15762 4117 -15756 4151
rect -15802 4079 -15756 4117
rect -15802 4045 -15796 4079
rect -15762 4045 -15756 4079
rect -15802 4007 -15756 4045
rect -15802 3973 -15796 4007
rect -15762 3973 -15756 4007
rect -15802 3935 -15756 3973
rect -15802 3901 -15796 3935
rect -15762 3901 -15756 3935
rect -15802 3863 -15756 3901
rect -15802 3829 -15796 3863
rect -15762 3829 -15756 3863
rect -15802 3791 -15756 3829
rect -15802 3757 -15796 3791
rect -15762 3757 -15756 3791
rect -15802 3719 -15756 3757
rect -15802 3685 -15796 3719
rect -15762 3685 -15756 3719
rect -15802 3647 -15756 3685
rect -15802 3613 -15796 3647
rect -15762 3613 -15756 3647
rect -15802 3575 -15756 3613
rect -15802 3541 -15796 3575
rect -15762 3541 -15756 3575
rect -15802 3503 -15756 3541
rect -15802 3469 -15796 3503
rect -15762 3469 -15756 3503
rect -15802 3454 -15756 3469
rect -15706 4439 -15660 4454
rect -15706 4405 -15700 4439
rect -15666 4405 -15660 4439
rect -15706 4367 -15660 4405
rect -15706 4333 -15700 4367
rect -15666 4333 -15660 4367
rect -15706 4295 -15660 4333
rect -15706 4261 -15700 4295
rect -15666 4261 -15660 4295
rect -15706 4223 -15660 4261
rect -15706 4189 -15700 4223
rect -15666 4189 -15660 4223
rect -15706 4151 -15660 4189
rect -15706 4117 -15700 4151
rect -15666 4117 -15660 4151
rect -15706 4079 -15660 4117
rect -15706 4045 -15700 4079
rect -15666 4045 -15660 4079
rect -15706 4007 -15660 4045
rect -15706 3973 -15700 4007
rect -15666 3973 -15660 4007
rect -15706 3935 -15660 3973
rect -15706 3901 -15700 3935
rect -15666 3901 -15660 3935
rect -15706 3863 -15660 3901
rect -15706 3829 -15700 3863
rect -15666 3829 -15660 3863
rect -15706 3791 -15660 3829
rect -15706 3757 -15700 3791
rect -15666 3757 -15660 3791
rect -15706 3719 -15660 3757
rect -15706 3685 -15700 3719
rect -15666 3685 -15660 3719
rect -15706 3647 -15660 3685
rect -15706 3613 -15700 3647
rect -15666 3613 -15660 3647
rect -15706 3575 -15660 3613
rect -15706 3541 -15700 3575
rect -15666 3541 -15660 3575
rect -15706 3503 -15660 3541
rect -15706 3469 -15700 3503
rect -15666 3469 -15660 3503
rect -15706 3454 -15660 3469
rect -15610 4439 -15564 4454
rect -15610 4405 -15604 4439
rect -15570 4405 -15564 4439
rect -15610 4367 -15564 4405
rect -15610 4333 -15604 4367
rect -15570 4333 -15564 4367
rect -15610 4295 -15564 4333
rect -15610 4261 -15604 4295
rect -15570 4261 -15564 4295
rect -15610 4223 -15564 4261
rect -15610 4189 -15604 4223
rect -15570 4189 -15564 4223
rect -15610 4151 -15564 4189
rect -15610 4117 -15604 4151
rect -15570 4117 -15564 4151
rect -15610 4079 -15564 4117
rect -15610 4045 -15604 4079
rect -15570 4045 -15564 4079
rect -15610 4007 -15564 4045
rect -15610 3973 -15604 4007
rect -15570 3973 -15564 4007
rect -15610 3935 -15564 3973
rect -15610 3901 -15604 3935
rect -15570 3901 -15564 3935
rect -15610 3863 -15564 3901
rect -15610 3829 -15604 3863
rect -15570 3829 -15564 3863
rect -15610 3791 -15564 3829
rect -15610 3757 -15604 3791
rect -15570 3757 -15564 3791
rect -15610 3719 -15564 3757
rect -15610 3685 -15604 3719
rect -15570 3685 -15564 3719
rect -15610 3647 -15564 3685
rect -15610 3613 -15604 3647
rect -15570 3613 -15564 3647
rect -15610 3575 -15564 3613
rect -15610 3541 -15604 3575
rect -15570 3541 -15564 3575
rect -15610 3503 -15564 3541
rect -15610 3469 -15604 3503
rect -15570 3469 -15564 3503
rect -15610 3454 -15564 3469
rect -15514 4439 -15468 4454
rect -15514 4405 -15508 4439
rect -15474 4405 -15468 4439
rect -15514 4367 -15468 4405
rect -15514 4333 -15508 4367
rect -15474 4333 -15468 4367
rect -15514 4295 -15468 4333
rect -15514 4261 -15508 4295
rect -15474 4261 -15468 4295
rect -15514 4223 -15468 4261
rect -15514 4189 -15508 4223
rect -15474 4189 -15468 4223
rect -15514 4151 -15468 4189
rect -15514 4117 -15508 4151
rect -15474 4117 -15468 4151
rect -15514 4079 -15468 4117
rect -15514 4045 -15508 4079
rect -15474 4045 -15468 4079
rect -15514 4007 -15468 4045
rect -15514 3973 -15508 4007
rect -15474 3973 -15468 4007
rect -15514 3935 -15468 3973
rect -15514 3901 -15508 3935
rect -15474 3901 -15468 3935
rect -15514 3863 -15468 3901
rect -15514 3829 -15508 3863
rect -15474 3829 -15468 3863
rect -15514 3791 -15468 3829
rect -15514 3757 -15508 3791
rect -15474 3757 -15468 3791
rect -15514 3719 -15468 3757
rect -15514 3685 -15508 3719
rect -15474 3685 -15468 3719
rect -15514 3647 -15468 3685
rect -15514 3613 -15508 3647
rect -15474 3613 -15468 3647
rect -15514 3575 -15468 3613
rect -15514 3541 -15508 3575
rect -15474 3541 -15468 3575
rect -15514 3503 -15468 3541
rect -15514 3469 -15508 3503
rect -15474 3469 -15468 3503
rect -15514 3454 -15468 3469
rect -15418 4439 -15372 4454
rect -15418 4405 -15412 4439
rect -15378 4405 -15372 4439
rect -15418 4367 -15372 4405
rect -15418 4333 -15412 4367
rect -15378 4333 -15372 4367
rect -15418 4295 -15372 4333
rect -15418 4261 -15412 4295
rect -15378 4261 -15372 4295
rect -15418 4223 -15372 4261
rect -15418 4189 -15412 4223
rect -15378 4189 -15372 4223
rect -15418 4151 -15372 4189
rect -15418 4117 -15412 4151
rect -15378 4117 -15372 4151
rect -15418 4079 -15372 4117
rect -15418 4045 -15412 4079
rect -15378 4045 -15372 4079
rect -15418 4007 -15372 4045
rect -15418 3973 -15412 4007
rect -15378 3973 -15372 4007
rect -15418 3935 -15372 3973
rect -15418 3901 -15412 3935
rect -15378 3901 -15372 3935
rect -15418 3863 -15372 3901
rect -15418 3829 -15412 3863
rect -15378 3829 -15372 3863
rect -15418 3791 -15372 3829
rect -15418 3757 -15412 3791
rect -15378 3757 -15372 3791
rect -15418 3719 -15372 3757
rect -15418 3685 -15412 3719
rect -15378 3685 -15372 3719
rect -15418 3647 -15372 3685
rect -15418 3613 -15412 3647
rect -15378 3613 -15372 3647
rect -15418 3575 -15372 3613
rect -15418 3541 -15412 3575
rect -15378 3541 -15372 3575
rect -15418 3503 -15372 3541
rect -15418 3469 -15412 3503
rect -15378 3469 -15372 3503
rect -15418 3454 -15372 3469
rect -15322 4439 -15276 4454
rect -15322 4405 -15316 4439
rect -15282 4405 -15276 4439
rect -15322 4367 -15276 4405
rect -15322 4333 -15316 4367
rect -15282 4333 -15276 4367
rect -15322 4295 -15276 4333
rect -15322 4261 -15316 4295
rect -15282 4261 -15276 4295
rect -15322 4223 -15276 4261
rect -15322 4189 -15316 4223
rect -15282 4189 -15276 4223
rect -15322 4151 -15276 4189
rect -15322 4117 -15316 4151
rect -15282 4117 -15276 4151
rect -15322 4079 -15276 4117
rect -15322 4045 -15316 4079
rect -15282 4045 -15276 4079
rect -15322 4007 -15276 4045
rect -15322 3973 -15316 4007
rect -15282 3973 -15276 4007
rect -15322 3935 -15276 3973
rect -15322 3901 -15316 3935
rect -15282 3901 -15276 3935
rect -15322 3863 -15276 3901
rect -15322 3829 -15316 3863
rect -15282 3829 -15276 3863
rect -15322 3791 -15276 3829
rect -15322 3757 -15316 3791
rect -15282 3757 -15276 3791
rect -15322 3719 -15276 3757
rect -15322 3685 -15316 3719
rect -15282 3685 -15276 3719
rect -15322 3647 -15276 3685
rect -15322 3613 -15316 3647
rect -15282 3613 -15276 3647
rect -15322 3575 -15276 3613
rect -15322 3541 -15316 3575
rect -15282 3541 -15276 3575
rect -15322 3503 -15276 3541
rect -15322 3469 -15316 3503
rect -15282 3469 -15276 3503
rect -15322 3454 -15276 3469
rect -15226 4439 -15180 4454
rect -15226 4405 -15220 4439
rect -15186 4405 -15180 4439
rect -15226 4367 -15180 4405
rect -15226 4333 -15220 4367
rect -15186 4333 -15180 4367
rect -15226 4295 -15180 4333
rect -15226 4261 -15220 4295
rect -15186 4261 -15180 4295
rect -15226 4223 -15180 4261
rect -15226 4189 -15220 4223
rect -15186 4189 -15180 4223
rect -15226 4151 -15180 4189
rect -15226 4117 -15220 4151
rect -15186 4117 -15180 4151
rect -15226 4079 -15180 4117
rect -15226 4045 -15220 4079
rect -15186 4045 -15180 4079
rect -15226 4007 -15180 4045
rect -15226 3973 -15220 4007
rect -15186 3973 -15180 4007
rect -15226 3935 -15180 3973
rect -15226 3901 -15220 3935
rect -15186 3901 -15180 3935
rect -15226 3863 -15180 3901
rect -15226 3829 -15220 3863
rect -15186 3829 -15180 3863
rect -15226 3791 -15180 3829
rect -15226 3757 -15220 3791
rect -15186 3757 -15180 3791
rect -15226 3719 -15180 3757
rect -15226 3685 -15220 3719
rect -15186 3685 -15180 3719
rect -15226 3647 -15180 3685
rect -15226 3613 -15220 3647
rect -15186 3613 -15180 3647
rect -15226 3575 -15180 3613
rect -15226 3541 -15220 3575
rect -15186 3541 -15180 3575
rect -15226 3503 -15180 3541
rect -15226 3469 -15220 3503
rect -15186 3469 -15180 3503
rect -15226 3454 -15180 3469
rect -15130 4439 -15084 4454
rect -15130 4405 -15124 4439
rect -15090 4405 -15084 4439
rect -15130 4367 -15084 4405
rect -15130 4333 -15124 4367
rect -15090 4333 -15084 4367
rect -15130 4295 -15084 4333
rect -15130 4261 -15124 4295
rect -15090 4261 -15084 4295
rect -15130 4223 -15084 4261
rect -15130 4189 -15124 4223
rect -15090 4189 -15084 4223
rect -15130 4151 -15084 4189
rect -15130 4117 -15124 4151
rect -15090 4117 -15084 4151
rect -15130 4079 -15084 4117
rect -15130 4045 -15124 4079
rect -15090 4045 -15084 4079
rect -15130 4007 -15084 4045
rect -15130 3973 -15124 4007
rect -15090 3973 -15084 4007
rect -15130 3935 -15084 3973
rect -15130 3901 -15124 3935
rect -15090 3901 -15084 3935
rect -15130 3863 -15084 3901
rect -15130 3829 -15124 3863
rect -15090 3829 -15084 3863
rect -15130 3791 -15084 3829
rect -15130 3757 -15124 3791
rect -15090 3757 -15084 3791
rect -15130 3719 -15084 3757
rect -15130 3685 -15124 3719
rect -15090 3685 -15084 3719
rect -15130 3647 -15084 3685
rect -15130 3613 -15124 3647
rect -15090 3613 -15084 3647
rect -15130 3575 -15084 3613
rect -15130 3541 -15124 3575
rect -15090 3541 -15084 3575
rect -15130 3503 -15084 3541
rect -15130 3469 -15124 3503
rect -15090 3469 -15084 3503
rect -15130 3454 -15084 3469
rect -15034 4439 -14988 4454
rect -15034 4405 -15028 4439
rect -14994 4405 -14988 4439
rect -15034 4367 -14988 4405
rect -15034 4333 -15028 4367
rect -14994 4333 -14988 4367
rect -15034 4295 -14988 4333
rect -15034 4261 -15028 4295
rect -14994 4261 -14988 4295
rect -15034 4223 -14988 4261
rect -15034 4189 -15028 4223
rect -14994 4189 -14988 4223
rect -15034 4151 -14988 4189
rect -15034 4117 -15028 4151
rect -14994 4117 -14988 4151
rect -15034 4079 -14988 4117
rect -15034 4045 -15028 4079
rect -14994 4045 -14988 4079
rect -15034 4007 -14988 4045
rect -15034 3973 -15028 4007
rect -14994 3973 -14988 4007
rect -15034 3935 -14988 3973
rect -15034 3901 -15028 3935
rect -14994 3901 -14988 3935
rect -15034 3863 -14988 3901
rect -15034 3829 -15028 3863
rect -14994 3829 -14988 3863
rect -15034 3791 -14988 3829
rect -15034 3757 -15028 3791
rect -14994 3757 -14988 3791
rect -15034 3719 -14988 3757
rect -15034 3685 -15028 3719
rect -14994 3685 -14988 3719
rect -15034 3647 -14988 3685
rect -15034 3613 -15028 3647
rect -14994 3613 -14988 3647
rect -15034 3575 -14988 3613
rect -15034 3541 -15028 3575
rect -14994 3541 -14988 3575
rect -15034 3503 -14988 3541
rect -15034 3469 -15028 3503
rect -14994 3469 -14988 3503
rect -15034 3454 -14988 3469
rect -14938 4439 -14892 4454
rect -14938 4405 -14932 4439
rect -14898 4405 -14892 4439
rect -14938 4367 -14892 4405
rect -14938 4333 -14932 4367
rect -14898 4333 -14892 4367
rect -14938 4295 -14892 4333
rect -14938 4261 -14932 4295
rect -14898 4261 -14892 4295
rect -14938 4223 -14892 4261
rect -14938 4189 -14932 4223
rect -14898 4189 -14892 4223
rect -14938 4151 -14892 4189
rect -14938 4117 -14932 4151
rect -14898 4117 -14892 4151
rect -14938 4079 -14892 4117
rect -14938 4045 -14932 4079
rect -14898 4045 -14892 4079
rect -14938 4007 -14892 4045
rect -14938 3973 -14932 4007
rect -14898 3973 -14892 4007
rect -14938 3935 -14892 3973
rect -14938 3901 -14932 3935
rect -14898 3901 -14892 3935
rect -14938 3863 -14892 3901
rect -14938 3829 -14932 3863
rect -14898 3829 -14892 3863
rect -14938 3791 -14892 3829
rect -14938 3757 -14932 3791
rect -14898 3757 -14892 3791
rect -14938 3719 -14892 3757
rect -14938 3685 -14932 3719
rect -14898 3685 -14892 3719
rect -14938 3647 -14892 3685
rect -14938 3613 -14932 3647
rect -14898 3613 -14892 3647
rect -14938 3575 -14892 3613
rect -14938 3541 -14932 3575
rect -14898 3541 -14892 3575
rect -14938 3503 -14892 3541
rect -14938 3469 -14932 3503
rect -14898 3469 -14892 3503
rect -14938 3454 -14892 3469
rect -14842 4439 -14796 4454
rect -14842 4405 -14836 4439
rect -14802 4405 -14796 4439
rect -14842 4367 -14796 4405
rect -14842 4333 -14836 4367
rect -14802 4333 -14796 4367
rect -14842 4295 -14796 4333
rect -14842 4261 -14836 4295
rect -14802 4261 -14796 4295
rect -14842 4223 -14796 4261
rect -14842 4189 -14836 4223
rect -14802 4189 -14796 4223
rect -14842 4151 -14796 4189
rect -14842 4117 -14836 4151
rect -14802 4117 -14796 4151
rect -14842 4079 -14796 4117
rect -14842 4045 -14836 4079
rect -14802 4045 -14796 4079
rect -14842 4007 -14796 4045
rect -14842 3973 -14836 4007
rect -14802 3973 -14796 4007
rect -14842 3935 -14796 3973
rect -14842 3901 -14836 3935
rect -14802 3901 -14796 3935
rect -14842 3863 -14796 3901
rect -14842 3829 -14836 3863
rect -14802 3829 -14796 3863
rect -14842 3791 -14796 3829
rect -14842 3757 -14836 3791
rect -14802 3757 -14796 3791
rect -14842 3719 -14796 3757
rect -14842 3685 -14836 3719
rect -14802 3685 -14796 3719
rect -14842 3647 -14796 3685
rect -14842 3613 -14836 3647
rect -14802 3613 -14796 3647
rect -14842 3575 -14796 3613
rect -14842 3541 -14836 3575
rect -14802 3541 -14796 3575
rect -14842 3503 -14796 3541
rect -14842 3469 -14836 3503
rect -14802 3469 -14796 3503
rect -14842 3454 -14796 3469
rect -14618 4445 -14572 4460
rect -14618 4411 -14612 4445
rect -14578 4411 -14572 4445
rect -14618 4373 -14572 4411
rect -14618 4339 -14612 4373
rect -14578 4339 -14572 4373
rect -14618 4301 -14572 4339
rect -14618 4267 -14612 4301
rect -14578 4267 -14572 4301
rect -14618 4229 -14572 4267
rect -14618 4195 -14612 4229
rect -14578 4195 -14572 4229
rect -14618 4157 -14572 4195
rect -14618 4123 -14612 4157
rect -14578 4123 -14572 4157
rect -14618 4085 -14572 4123
rect -14618 4051 -14612 4085
rect -14578 4051 -14572 4085
rect -14618 4013 -14572 4051
rect -14618 3979 -14612 4013
rect -14578 3979 -14572 4013
rect -14618 3941 -14572 3979
rect -14618 3907 -14612 3941
rect -14578 3907 -14572 3941
rect -14618 3869 -14572 3907
rect -14618 3835 -14612 3869
rect -14578 3835 -14572 3869
rect -14618 3797 -14572 3835
rect -14618 3763 -14612 3797
rect -14578 3763 -14572 3797
rect -14618 3725 -14572 3763
rect -14618 3691 -14612 3725
rect -14578 3691 -14572 3725
rect -14618 3653 -14572 3691
rect -14618 3619 -14612 3653
rect -14578 3619 -14572 3653
rect -14618 3581 -14572 3619
rect -14618 3547 -14612 3581
rect -14578 3547 -14572 3581
rect -14618 3509 -14572 3547
rect -14618 3475 -14612 3509
rect -14578 3475 -14572 3509
rect -14618 3460 -14572 3475
rect -14522 4445 -14476 4460
rect -14522 4411 -14516 4445
rect -14482 4411 -14476 4445
rect -14522 4373 -14476 4411
rect -14522 4339 -14516 4373
rect -14482 4339 -14476 4373
rect -14522 4301 -14476 4339
rect -14522 4267 -14516 4301
rect -14482 4267 -14476 4301
rect -14522 4229 -14476 4267
rect -14522 4195 -14516 4229
rect -14482 4195 -14476 4229
rect -14522 4157 -14476 4195
rect -14522 4123 -14516 4157
rect -14482 4123 -14476 4157
rect -14522 4085 -14476 4123
rect -14522 4051 -14516 4085
rect -14482 4051 -14476 4085
rect -14522 4013 -14476 4051
rect -14522 3979 -14516 4013
rect -14482 3979 -14476 4013
rect -14522 3941 -14476 3979
rect -14522 3907 -14516 3941
rect -14482 3907 -14476 3941
rect -14522 3869 -14476 3907
rect -14522 3835 -14516 3869
rect -14482 3835 -14476 3869
rect -14522 3797 -14476 3835
rect -14522 3763 -14516 3797
rect -14482 3763 -14476 3797
rect -14522 3725 -14476 3763
rect -14522 3691 -14516 3725
rect -14482 3691 -14476 3725
rect -14522 3653 -14476 3691
rect -14522 3619 -14516 3653
rect -14482 3619 -14476 3653
rect -14522 3581 -14476 3619
rect -14522 3547 -14516 3581
rect -14482 3547 -14476 3581
rect -14522 3509 -14476 3547
rect -14522 3475 -14516 3509
rect -14482 3475 -14476 3509
rect -14522 3460 -14476 3475
rect -14426 4445 -14380 4460
rect -14426 4411 -14420 4445
rect -14386 4411 -14380 4445
rect -14426 4373 -14380 4411
rect -14426 4339 -14420 4373
rect -14386 4339 -14380 4373
rect -14426 4301 -14380 4339
rect -14426 4267 -14420 4301
rect -14386 4267 -14380 4301
rect -14426 4229 -14380 4267
rect -14426 4195 -14420 4229
rect -14386 4195 -14380 4229
rect -14426 4157 -14380 4195
rect -14426 4123 -14420 4157
rect -14386 4123 -14380 4157
rect -14426 4085 -14380 4123
rect -14426 4051 -14420 4085
rect -14386 4051 -14380 4085
rect -14426 4013 -14380 4051
rect -14426 3979 -14420 4013
rect -14386 3979 -14380 4013
rect -14426 3941 -14380 3979
rect -14426 3907 -14420 3941
rect -14386 3907 -14380 3941
rect -14426 3869 -14380 3907
rect -14426 3835 -14420 3869
rect -14386 3835 -14380 3869
rect -14426 3797 -14380 3835
rect -14426 3763 -14420 3797
rect -14386 3763 -14380 3797
rect -14426 3725 -14380 3763
rect -14426 3691 -14420 3725
rect -14386 3691 -14380 3725
rect -14426 3653 -14380 3691
rect -14426 3619 -14420 3653
rect -14386 3619 -14380 3653
rect -14426 3581 -14380 3619
rect -14426 3547 -14420 3581
rect -14386 3547 -14380 3581
rect -14426 3509 -14380 3547
rect -14426 3475 -14420 3509
rect -14386 3475 -14380 3509
rect -14426 3460 -14380 3475
rect -14330 4445 -14284 4460
rect -14330 4411 -14324 4445
rect -14290 4411 -14284 4445
rect -14330 4373 -14284 4411
rect -14330 4339 -14324 4373
rect -14290 4339 -14284 4373
rect -14330 4301 -14284 4339
rect -14330 4267 -14324 4301
rect -14290 4267 -14284 4301
rect -14330 4229 -14284 4267
rect -14330 4195 -14324 4229
rect -14290 4195 -14284 4229
rect -14330 4157 -14284 4195
rect -14330 4123 -14324 4157
rect -14290 4123 -14284 4157
rect -14330 4085 -14284 4123
rect -14330 4051 -14324 4085
rect -14290 4051 -14284 4085
rect -14330 4013 -14284 4051
rect -14330 3979 -14324 4013
rect -14290 3979 -14284 4013
rect -14330 3941 -14284 3979
rect -14330 3907 -14324 3941
rect -14290 3907 -14284 3941
rect -14330 3869 -14284 3907
rect -14330 3835 -14324 3869
rect -14290 3835 -14284 3869
rect -14330 3797 -14284 3835
rect -14330 3763 -14324 3797
rect -14290 3763 -14284 3797
rect -14330 3725 -14284 3763
rect -14330 3691 -14324 3725
rect -14290 3691 -14284 3725
rect -14330 3653 -14284 3691
rect -14330 3619 -14324 3653
rect -14290 3619 -14284 3653
rect -14330 3581 -14284 3619
rect -14330 3547 -14324 3581
rect -14290 3547 -14284 3581
rect -14330 3509 -14284 3547
rect -14330 3475 -14324 3509
rect -14290 3475 -14284 3509
rect -14330 3460 -14284 3475
rect -14234 4445 -14188 4460
rect -14234 4411 -14228 4445
rect -14194 4411 -14188 4445
rect -14234 4373 -14188 4411
rect -14234 4339 -14228 4373
rect -14194 4339 -14188 4373
rect -14234 4301 -14188 4339
rect -14234 4267 -14228 4301
rect -14194 4267 -14188 4301
rect -14234 4229 -14188 4267
rect -14234 4195 -14228 4229
rect -14194 4195 -14188 4229
rect -14234 4157 -14188 4195
rect -14234 4123 -14228 4157
rect -14194 4123 -14188 4157
rect -14234 4085 -14188 4123
rect -14234 4051 -14228 4085
rect -14194 4051 -14188 4085
rect -14234 4013 -14188 4051
rect -14234 3979 -14228 4013
rect -14194 3979 -14188 4013
rect -14234 3941 -14188 3979
rect -14234 3907 -14228 3941
rect -14194 3907 -14188 3941
rect -14234 3869 -14188 3907
rect -14234 3835 -14228 3869
rect -14194 3835 -14188 3869
rect -14234 3797 -14188 3835
rect -14234 3763 -14228 3797
rect -14194 3763 -14188 3797
rect -14234 3725 -14188 3763
rect -14234 3691 -14228 3725
rect -14194 3691 -14188 3725
rect -14234 3653 -14188 3691
rect -14234 3619 -14228 3653
rect -14194 3619 -14188 3653
rect -14234 3581 -14188 3619
rect -14234 3547 -14228 3581
rect -14194 3547 -14188 3581
rect -14234 3509 -14188 3547
rect -14234 3475 -14228 3509
rect -14194 3475 -14188 3509
rect -14234 3460 -14188 3475
rect -14138 4445 -14092 4460
rect -14138 4411 -14132 4445
rect -14098 4411 -14092 4445
rect -14138 4373 -14092 4411
rect -14138 4339 -14132 4373
rect -14098 4339 -14092 4373
rect -14138 4301 -14092 4339
rect -14138 4267 -14132 4301
rect -14098 4267 -14092 4301
rect -14138 4229 -14092 4267
rect -14138 4195 -14132 4229
rect -14098 4195 -14092 4229
rect -14138 4157 -14092 4195
rect -14138 4123 -14132 4157
rect -14098 4123 -14092 4157
rect -14138 4085 -14092 4123
rect -14138 4051 -14132 4085
rect -14098 4051 -14092 4085
rect -14138 4013 -14092 4051
rect -14138 3979 -14132 4013
rect -14098 3979 -14092 4013
rect -14138 3941 -14092 3979
rect -14138 3907 -14132 3941
rect -14098 3907 -14092 3941
rect -14138 3869 -14092 3907
rect -14138 3835 -14132 3869
rect -14098 3835 -14092 3869
rect -14138 3797 -14092 3835
rect -14138 3763 -14132 3797
rect -14098 3763 -14092 3797
rect -14138 3725 -14092 3763
rect -14138 3691 -14132 3725
rect -14098 3691 -14092 3725
rect -14138 3653 -14092 3691
rect -14138 3619 -14132 3653
rect -14098 3619 -14092 3653
rect -14138 3581 -14092 3619
rect -14138 3547 -14132 3581
rect -14098 3547 -14092 3581
rect -14138 3509 -14092 3547
rect -14138 3475 -14132 3509
rect -14098 3475 -14092 3509
rect -14138 3460 -14092 3475
rect -14042 4445 -13996 4460
rect -14042 4411 -14036 4445
rect -14002 4411 -13996 4445
rect -14042 4373 -13996 4411
rect -14042 4339 -14036 4373
rect -14002 4339 -13996 4373
rect -14042 4301 -13996 4339
rect -14042 4267 -14036 4301
rect -14002 4267 -13996 4301
rect -14042 4229 -13996 4267
rect -14042 4195 -14036 4229
rect -14002 4195 -13996 4229
rect -14042 4157 -13996 4195
rect -14042 4123 -14036 4157
rect -14002 4123 -13996 4157
rect -14042 4085 -13996 4123
rect -14042 4051 -14036 4085
rect -14002 4051 -13996 4085
rect -14042 4013 -13996 4051
rect -14042 3979 -14036 4013
rect -14002 3979 -13996 4013
rect -14042 3941 -13996 3979
rect -14042 3907 -14036 3941
rect -14002 3907 -13996 3941
rect -14042 3869 -13996 3907
rect -14042 3835 -14036 3869
rect -14002 3835 -13996 3869
rect -14042 3797 -13996 3835
rect -14042 3763 -14036 3797
rect -14002 3763 -13996 3797
rect -14042 3725 -13996 3763
rect -14042 3691 -14036 3725
rect -14002 3691 -13996 3725
rect -14042 3653 -13996 3691
rect -14042 3619 -14036 3653
rect -14002 3619 -13996 3653
rect -14042 3581 -13996 3619
rect -14042 3547 -14036 3581
rect -14002 3547 -13996 3581
rect -14042 3509 -13996 3547
rect -14042 3475 -14036 3509
rect -14002 3475 -13996 3509
rect -14042 3460 -13996 3475
rect -13946 4445 -13900 4460
rect -13946 4411 -13940 4445
rect -13906 4411 -13900 4445
rect -13946 4373 -13900 4411
rect -13946 4339 -13940 4373
rect -13906 4339 -13900 4373
rect -13946 4301 -13900 4339
rect -13946 4267 -13940 4301
rect -13906 4267 -13900 4301
rect -13946 4229 -13900 4267
rect -13946 4195 -13940 4229
rect -13906 4195 -13900 4229
rect -13946 4157 -13900 4195
rect -13946 4123 -13940 4157
rect -13906 4123 -13900 4157
rect -13946 4085 -13900 4123
rect -13946 4051 -13940 4085
rect -13906 4051 -13900 4085
rect -13946 4013 -13900 4051
rect -13946 3979 -13940 4013
rect -13906 3979 -13900 4013
rect -13946 3941 -13900 3979
rect -13946 3907 -13940 3941
rect -13906 3907 -13900 3941
rect -13946 3869 -13900 3907
rect -13946 3835 -13940 3869
rect -13906 3835 -13900 3869
rect -13946 3797 -13900 3835
rect -13946 3763 -13940 3797
rect -13906 3763 -13900 3797
rect -13946 3725 -13900 3763
rect -13946 3691 -13940 3725
rect -13906 3691 -13900 3725
rect -13946 3653 -13900 3691
rect -13946 3619 -13940 3653
rect -13906 3619 -13900 3653
rect -13946 3581 -13900 3619
rect -13946 3547 -13940 3581
rect -13906 3547 -13900 3581
rect -13946 3509 -13900 3547
rect -13946 3475 -13940 3509
rect -13906 3475 -13900 3509
rect -13946 3460 -13900 3475
rect -13850 4445 -13804 4460
rect -13850 4411 -13844 4445
rect -13810 4411 -13804 4445
rect -13850 4373 -13804 4411
rect -13850 4339 -13844 4373
rect -13810 4339 -13804 4373
rect -13850 4301 -13804 4339
rect -13850 4267 -13844 4301
rect -13810 4267 -13804 4301
rect -13850 4229 -13804 4267
rect -13850 4195 -13844 4229
rect -13810 4195 -13804 4229
rect -13850 4157 -13804 4195
rect -13850 4123 -13844 4157
rect -13810 4123 -13804 4157
rect -13850 4085 -13804 4123
rect -13850 4051 -13844 4085
rect -13810 4051 -13804 4085
rect -13850 4013 -13804 4051
rect -13850 3979 -13844 4013
rect -13810 3979 -13804 4013
rect -13850 3941 -13804 3979
rect -13850 3907 -13844 3941
rect -13810 3907 -13804 3941
rect -13850 3869 -13804 3907
rect -13850 3835 -13844 3869
rect -13810 3835 -13804 3869
rect -13850 3797 -13804 3835
rect -13850 3763 -13844 3797
rect -13810 3763 -13804 3797
rect -13850 3725 -13804 3763
rect -13850 3691 -13844 3725
rect -13810 3691 -13804 3725
rect -13850 3653 -13804 3691
rect -13850 3619 -13844 3653
rect -13810 3619 -13804 3653
rect -13850 3581 -13804 3619
rect -13850 3547 -13844 3581
rect -13810 3547 -13804 3581
rect -13850 3509 -13804 3547
rect -13850 3475 -13844 3509
rect -13810 3475 -13804 3509
rect -13850 3460 -13804 3475
rect -13754 4445 -13708 4460
rect -13754 4411 -13748 4445
rect -13714 4411 -13708 4445
rect -13754 4373 -13708 4411
rect -13754 4339 -13748 4373
rect -13714 4339 -13708 4373
rect -13754 4301 -13708 4339
rect -13754 4267 -13748 4301
rect -13714 4267 -13708 4301
rect -13754 4229 -13708 4267
rect -13754 4195 -13748 4229
rect -13714 4195 -13708 4229
rect -13754 4157 -13708 4195
rect -13754 4123 -13748 4157
rect -13714 4123 -13708 4157
rect -13754 4085 -13708 4123
rect -13754 4051 -13748 4085
rect -13714 4051 -13708 4085
rect -13754 4013 -13708 4051
rect -13754 3979 -13748 4013
rect -13714 3979 -13708 4013
rect -13754 3941 -13708 3979
rect -13754 3907 -13748 3941
rect -13714 3907 -13708 3941
rect -13754 3869 -13708 3907
rect -13754 3835 -13748 3869
rect -13714 3835 -13708 3869
rect -13754 3797 -13708 3835
rect -13754 3763 -13748 3797
rect -13714 3763 -13708 3797
rect -13754 3725 -13708 3763
rect -13754 3691 -13748 3725
rect -13714 3691 -13708 3725
rect -13754 3653 -13708 3691
rect -13754 3619 -13748 3653
rect -13714 3619 -13708 3653
rect -13754 3581 -13708 3619
rect -13754 3547 -13748 3581
rect -13714 3547 -13708 3581
rect -13754 3509 -13708 3547
rect -13754 3475 -13748 3509
rect -13714 3475 -13708 3509
rect -13754 3460 -13708 3475
rect -13658 4445 -13612 4460
rect -13658 4411 -13652 4445
rect -13618 4411 -13612 4445
rect -13658 4373 -13612 4411
rect -13658 4339 -13652 4373
rect -13618 4339 -13612 4373
rect -13658 4301 -13612 4339
rect -13658 4267 -13652 4301
rect -13618 4267 -13612 4301
rect -13658 4229 -13612 4267
rect -13658 4195 -13652 4229
rect -13618 4195 -13612 4229
rect -13658 4157 -13612 4195
rect -13658 4123 -13652 4157
rect -13618 4123 -13612 4157
rect -13658 4085 -13612 4123
rect -13658 4051 -13652 4085
rect -13618 4051 -13612 4085
rect -13658 4013 -13612 4051
rect -13658 3979 -13652 4013
rect -13618 3979 -13612 4013
rect -13658 3941 -13612 3979
rect -13658 3907 -13652 3941
rect -13618 3907 -13612 3941
rect -13658 3869 -13612 3907
rect -13658 3835 -13652 3869
rect -13618 3835 -13612 3869
rect -13658 3797 -13612 3835
rect -13658 3763 -13652 3797
rect -13618 3763 -13612 3797
rect -13658 3725 -13612 3763
rect -13658 3691 -13652 3725
rect -13618 3691 -13612 3725
rect -13658 3653 -13612 3691
rect -13658 3619 -13652 3653
rect -13618 3619 -13612 3653
rect -13658 3581 -13612 3619
rect -13658 3547 -13652 3581
rect -13618 3547 -13612 3581
rect -13658 3509 -13612 3547
rect -13658 3475 -13652 3509
rect -13618 3475 -13612 3509
rect -13658 3460 -13612 3475
rect -13562 4445 -13516 4460
rect -13562 4411 -13556 4445
rect -13522 4411 -13516 4445
rect -13562 4373 -13516 4411
rect -13562 4339 -13556 4373
rect -13522 4339 -13516 4373
rect -13562 4301 -13516 4339
rect -13562 4267 -13556 4301
rect -13522 4267 -13516 4301
rect -13562 4229 -13516 4267
rect -13562 4195 -13556 4229
rect -13522 4195 -13516 4229
rect -13562 4157 -13516 4195
rect -13562 4123 -13556 4157
rect -13522 4123 -13516 4157
rect -13562 4085 -13516 4123
rect -13562 4051 -13556 4085
rect -13522 4051 -13516 4085
rect -13562 4013 -13516 4051
rect -13562 3979 -13556 4013
rect -13522 3979 -13516 4013
rect -13562 3941 -13516 3979
rect -13562 3907 -13556 3941
rect -13522 3907 -13516 3941
rect -13562 3869 -13516 3907
rect -13562 3835 -13556 3869
rect -13522 3835 -13516 3869
rect -13562 3797 -13516 3835
rect -13562 3763 -13556 3797
rect -13522 3763 -13516 3797
rect -13562 3725 -13516 3763
rect -13562 3691 -13556 3725
rect -13522 3691 -13516 3725
rect -13562 3653 -13516 3691
rect -13562 3619 -13556 3653
rect -13522 3619 -13516 3653
rect -13562 3581 -13516 3619
rect -13562 3547 -13556 3581
rect -13522 3547 -13516 3581
rect -13562 3509 -13516 3547
rect -13562 3475 -13556 3509
rect -13522 3475 -13516 3509
rect -13562 3460 -13516 3475
rect -13466 4445 -13420 4460
rect -13466 4411 -13460 4445
rect -13426 4411 -13420 4445
rect -13466 4373 -13420 4411
rect -13466 4339 -13460 4373
rect -13426 4339 -13420 4373
rect -13466 4301 -13420 4339
rect -13466 4267 -13460 4301
rect -13426 4267 -13420 4301
rect -13466 4229 -13420 4267
rect -13466 4195 -13460 4229
rect -13426 4195 -13420 4229
rect -13466 4157 -13420 4195
rect -13466 4123 -13460 4157
rect -13426 4123 -13420 4157
rect -13466 4085 -13420 4123
rect -13466 4051 -13460 4085
rect -13426 4051 -13420 4085
rect -13466 4013 -13420 4051
rect -13466 3979 -13460 4013
rect -13426 3979 -13420 4013
rect -13466 3941 -13420 3979
rect -13466 3907 -13460 3941
rect -13426 3907 -13420 3941
rect -13466 3869 -13420 3907
rect -13466 3835 -13460 3869
rect -13426 3835 -13420 3869
rect -13466 3797 -13420 3835
rect -13466 3763 -13460 3797
rect -13426 3763 -13420 3797
rect -13466 3725 -13420 3763
rect -13466 3691 -13460 3725
rect -13426 3691 -13420 3725
rect -13466 3653 -13420 3691
rect -13466 3619 -13460 3653
rect -13426 3619 -13420 3653
rect -13466 3581 -13420 3619
rect -13466 3547 -13460 3581
rect -13426 3547 -13420 3581
rect -13466 3509 -13420 3547
rect -13466 3475 -13460 3509
rect -13426 3475 -13420 3509
rect -13466 3460 -13420 3475
rect -13370 4445 -13324 4460
rect -13370 4411 -13364 4445
rect -13330 4411 -13324 4445
rect -13370 4373 -13324 4411
rect -13370 4339 -13364 4373
rect -13330 4339 -13324 4373
rect -13370 4301 -13324 4339
rect -13370 4267 -13364 4301
rect -13330 4267 -13324 4301
rect -13370 4229 -13324 4267
rect -13370 4195 -13364 4229
rect -13330 4195 -13324 4229
rect -13370 4157 -13324 4195
rect -13370 4123 -13364 4157
rect -13330 4123 -13324 4157
rect -13370 4085 -13324 4123
rect -13370 4051 -13364 4085
rect -13330 4051 -13324 4085
rect -13370 4013 -13324 4051
rect -13370 3979 -13364 4013
rect -13330 3979 -13324 4013
rect -13370 3941 -13324 3979
rect -13370 3907 -13364 3941
rect -13330 3907 -13324 3941
rect -13370 3869 -13324 3907
rect -13370 3835 -13364 3869
rect -13330 3835 -13324 3869
rect -13370 3797 -13324 3835
rect -13370 3763 -13364 3797
rect -13330 3763 -13324 3797
rect -13370 3725 -13324 3763
rect -13370 3691 -13364 3725
rect -13330 3691 -13324 3725
rect -13370 3653 -13324 3691
rect -13370 3619 -13364 3653
rect -13330 3619 -13324 3653
rect -13370 3581 -13324 3619
rect -13370 3547 -13364 3581
rect -13330 3547 -13324 3581
rect -13370 3509 -13324 3547
rect -13370 3475 -13364 3509
rect -13330 3475 -13324 3509
rect -13370 3460 -13324 3475
rect -13274 4445 -13228 4460
rect -13274 4411 -13268 4445
rect -13234 4411 -13228 4445
rect -13274 4373 -13228 4411
rect -13274 4339 -13268 4373
rect -13234 4339 -13228 4373
rect -13274 4301 -13228 4339
rect -13274 4267 -13268 4301
rect -13234 4267 -13228 4301
rect -13274 4229 -13228 4267
rect -13274 4195 -13268 4229
rect -13234 4195 -13228 4229
rect -13274 4157 -13228 4195
rect -13274 4123 -13268 4157
rect -13234 4123 -13228 4157
rect -13274 4085 -13228 4123
rect -13274 4051 -13268 4085
rect -13234 4051 -13228 4085
rect -13274 4013 -13228 4051
rect -13274 3979 -13268 4013
rect -13234 3979 -13228 4013
rect -13274 3941 -13228 3979
rect -13274 3907 -13268 3941
rect -13234 3907 -13228 3941
rect -13274 3869 -13228 3907
rect -13274 3835 -13268 3869
rect -13234 3835 -13228 3869
rect -13274 3797 -13228 3835
rect -13274 3763 -13268 3797
rect -13234 3763 -13228 3797
rect -13274 3725 -13228 3763
rect -13274 3691 -13268 3725
rect -13234 3691 -13228 3725
rect -13274 3653 -13228 3691
rect -13274 3619 -13268 3653
rect -13234 3619 -13228 3653
rect -13274 3581 -13228 3619
rect -13274 3547 -13268 3581
rect -13234 3547 -13228 3581
rect -13274 3509 -13228 3547
rect -13274 3475 -13268 3509
rect -13234 3475 -13228 3509
rect -13274 3460 -13228 3475
rect -13178 4445 -13132 4460
rect -13178 4411 -13172 4445
rect -13138 4411 -13132 4445
rect -13178 4373 -13132 4411
rect -13178 4339 -13172 4373
rect -13138 4339 -13132 4373
rect -13178 4301 -13132 4339
rect -13178 4267 -13172 4301
rect -13138 4267 -13132 4301
rect -13178 4229 -13132 4267
rect -13178 4195 -13172 4229
rect -13138 4195 -13132 4229
rect -13178 4157 -13132 4195
rect -13178 4123 -13172 4157
rect -13138 4123 -13132 4157
rect -13178 4085 -13132 4123
rect -13178 4051 -13172 4085
rect -13138 4051 -13132 4085
rect -13178 4013 -13132 4051
rect -13178 3979 -13172 4013
rect -13138 3979 -13132 4013
rect -13178 3941 -13132 3979
rect -13178 3907 -13172 3941
rect -13138 3907 -13132 3941
rect -13178 3869 -13132 3907
rect -13178 3835 -13172 3869
rect -13138 3835 -13132 3869
rect -13178 3797 -13132 3835
rect -13178 3763 -13172 3797
rect -13138 3763 -13132 3797
rect -13178 3725 -13132 3763
rect -13178 3691 -13172 3725
rect -13138 3691 -13132 3725
rect -13178 3653 -13132 3691
rect -13178 3619 -13172 3653
rect -13138 3619 -13132 3653
rect -13178 3581 -13132 3619
rect -13178 3547 -13172 3581
rect -13138 3547 -13132 3581
rect -13178 3509 -13132 3547
rect -13178 3475 -13172 3509
rect -13138 3475 -13132 3509
rect -13178 3460 -13132 3475
rect -12934 4451 -12888 4466
rect -12934 4417 -12928 4451
rect -12894 4417 -12888 4451
rect -12934 4379 -12888 4417
rect -12934 4345 -12928 4379
rect -12894 4345 -12888 4379
rect -12934 4307 -12888 4345
rect -12934 4273 -12928 4307
rect -12894 4273 -12888 4307
rect -12934 4235 -12888 4273
rect -12934 4201 -12928 4235
rect -12894 4201 -12888 4235
rect -12934 4163 -12888 4201
rect -12934 4129 -12928 4163
rect -12894 4129 -12888 4163
rect -12934 4091 -12888 4129
rect -12934 4057 -12928 4091
rect -12894 4057 -12888 4091
rect -12934 4019 -12888 4057
rect -12934 3985 -12928 4019
rect -12894 3985 -12888 4019
rect -12934 3947 -12888 3985
rect -12934 3913 -12928 3947
rect -12894 3913 -12888 3947
rect -12934 3875 -12888 3913
rect -12934 3841 -12928 3875
rect -12894 3841 -12888 3875
rect -12934 3803 -12888 3841
rect -12934 3769 -12928 3803
rect -12894 3769 -12888 3803
rect -12934 3731 -12888 3769
rect -12934 3697 -12928 3731
rect -12894 3697 -12888 3731
rect -12934 3659 -12888 3697
rect -12934 3625 -12928 3659
rect -12894 3625 -12888 3659
rect -12934 3587 -12888 3625
rect -12934 3553 -12928 3587
rect -12894 3553 -12888 3587
rect -12934 3515 -12888 3553
rect -12934 3481 -12928 3515
rect -12894 3481 -12888 3515
rect -12934 3466 -12888 3481
rect -12838 4451 -12792 4466
rect -12838 4417 -12832 4451
rect -12798 4417 -12792 4451
rect -12838 4379 -12792 4417
rect -12838 4345 -12832 4379
rect -12798 4345 -12792 4379
rect -12838 4307 -12792 4345
rect -12838 4273 -12832 4307
rect -12798 4273 -12792 4307
rect -12838 4235 -12792 4273
rect -12838 4201 -12832 4235
rect -12798 4201 -12792 4235
rect -12838 4163 -12792 4201
rect -12838 4129 -12832 4163
rect -12798 4129 -12792 4163
rect -12838 4091 -12792 4129
rect -12838 4057 -12832 4091
rect -12798 4057 -12792 4091
rect -12838 4019 -12792 4057
rect -12838 3985 -12832 4019
rect -12798 3985 -12792 4019
rect -12838 3947 -12792 3985
rect -12838 3913 -12832 3947
rect -12798 3913 -12792 3947
rect -12838 3875 -12792 3913
rect -12838 3841 -12832 3875
rect -12798 3841 -12792 3875
rect -12838 3803 -12792 3841
rect -12838 3769 -12832 3803
rect -12798 3769 -12792 3803
rect -12838 3731 -12792 3769
rect -12838 3697 -12832 3731
rect -12798 3697 -12792 3731
rect -12838 3659 -12792 3697
rect -12838 3625 -12832 3659
rect -12798 3625 -12792 3659
rect -12838 3587 -12792 3625
rect -12838 3553 -12832 3587
rect -12798 3553 -12792 3587
rect -12838 3515 -12792 3553
rect -12838 3481 -12832 3515
rect -12798 3481 -12792 3515
rect -12838 3466 -12792 3481
rect -12742 4451 -12696 4466
rect -12742 4417 -12736 4451
rect -12702 4417 -12696 4451
rect -12742 4379 -12696 4417
rect -12742 4345 -12736 4379
rect -12702 4345 -12696 4379
rect -12742 4307 -12696 4345
rect -12742 4273 -12736 4307
rect -12702 4273 -12696 4307
rect -12742 4235 -12696 4273
rect -12742 4201 -12736 4235
rect -12702 4201 -12696 4235
rect -12742 4163 -12696 4201
rect -12742 4129 -12736 4163
rect -12702 4129 -12696 4163
rect -12742 4091 -12696 4129
rect -12742 4057 -12736 4091
rect -12702 4057 -12696 4091
rect -12742 4019 -12696 4057
rect -12742 3985 -12736 4019
rect -12702 3985 -12696 4019
rect -12742 3947 -12696 3985
rect -12742 3913 -12736 3947
rect -12702 3913 -12696 3947
rect -12742 3875 -12696 3913
rect -12742 3841 -12736 3875
rect -12702 3841 -12696 3875
rect -12742 3803 -12696 3841
rect -12742 3769 -12736 3803
rect -12702 3769 -12696 3803
rect -12742 3731 -12696 3769
rect -12742 3697 -12736 3731
rect -12702 3697 -12696 3731
rect -12742 3659 -12696 3697
rect -12742 3625 -12736 3659
rect -12702 3625 -12696 3659
rect -12742 3587 -12696 3625
rect -12742 3553 -12736 3587
rect -12702 3553 -12696 3587
rect -12742 3515 -12696 3553
rect -12742 3481 -12736 3515
rect -12702 3481 -12696 3515
rect -12742 3466 -12696 3481
rect -12646 4451 -12600 4466
rect -12646 4417 -12640 4451
rect -12606 4417 -12600 4451
rect -12646 4379 -12600 4417
rect -12646 4345 -12640 4379
rect -12606 4345 -12600 4379
rect -12646 4307 -12600 4345
rect -12646 4273 -12640 4307
rect -12606 4273 -12600 4307
rect -12646 4235 -12600 4273
rect -12646 4201 -12640 4235
rect -12606 4201 -12600 4235
rect -12646 4163 -12600 4201
rect -12646 4129 -12640 4163
rect -12606 4129 -12600 4163
rect -12646 4091 -12600 4129
rect -12646 4057 -12640 4091
rect -12606 4057 -12600 4091
rect -12646 4019 -12600 4057
rect -12646 3985 -12640 4019
rect -12606 3985 -12600 4019
rect -12646 3947 -12600 3985
rect -12646 3913 -12640 3947
rect -12606 3913 -12600 3947
rect -12646 3875 -12600 3913
rect -12646 3841 -12640 3875
rect -12606 3841 -12600 3875
rect -12646 3803 -12600 3841
rect -12646 3769 -12640 3803
rect -12606 3769 -12600 3803
rect -12646 3731 -12600 3769
rect -12646 3697 -12640 3731
rect -12606 3697 -12600 3731
rect -12646 3659 -12600 3697
rect -12646 3625 -12640 3659
rect -12606 3625 -12600 3659
rect -12646 3587 -12600 3625
rect -12646 3553 -12640 3587
rect -12606 3553 -12600 3587
rect -12646 3515 -12600 3553
rect -12646 3481 -12640 3515
rect -12606 3481 -12600 3515
rect -12646 3466 -12600 3481
rect -12550 4451 -12504 4466
rect -12550 4417 -12544 4451
rect -12510 4417 -12504 4451
rect -12550 4379 -12504 4417
rect -12550 4345 -12544 4379
rect -12510 4345 -12504 4379
rect -12550 4307 -12504 4345
rect -12550 4273 -12544 4307
rect -12510 4273 -12504 4307
rect -12550 4235 -12504 4273
rect -12550 4201 -12544 4235
rect -12510 4201 -12504 4235
rect -12550 4163 -12504 4201
rect -12550 4129 -12544 4163
rect -12510 4129 -12504 4163
rect -12550 4091 -12504 4129
rect -12550 4057 -12544 4091
rect -12510 4057 -12504 4091
rect -12550 4019 -12504 4057
rect -12550 3985 -12544 4019
rect -12510 3985 -12504 4019
rect -12550 3947 -12504 3985
rect -12550 3913 -12544 3947
rect -12510 3913 -12504 3947
rect -12550 3875 -12504 3913
rect -12550 3841 -12544 3875
rect -12510 3841 -12504 3875
rect -12550 3803 -12504 3841
rect -12550 3769 -12544 3803
rect -12510 3769 -12504 3803
rect -12550 3731 -12504 3769
rect -12550 3697 -12544 3731
rect -12510 3697 -12504 3731
rect -12550 3659 -12504 3697
rect -12550 3625 -12544 3659
rect -12510 3625 -12504 3659
rect -12550 3587 -12504 3625
rect -12550 3553 -12544 3587
rect -12510 3553 -12504 3587
rect -12550 3515 -12504 3553
rect -12550 3481 -12544 3515
rect -12510 3481 -12504 3515
rect -12550 3466 -12504 3481
rect -12454 4451 -12408 4466
rect -12454 4417 -12448 4451
rect -12414 4417 -12408 4451
rect -12454 4379 -12408 4417
rect -12454 4345 -12448 4379
rect -12414 4345 -12408 4379
rect -12454 4307 -12408 4345
rect -12454 4273 -12448 4307
rect -12414 4273 -12408 4307
rect -12454 4235 -12408 4273
rect -12454 4201 -12448 4235
rect -12414 4201 -12408 4235
rect -12454 4163 -12408 4201
rect -12454 4129 -12448 4163
rect -12414 4129 -12408 4163
rect -12454 4091 -12408 4129
rect -12454 4057 -12448 4091
rect -12414 4057 -12408 4091
rect -12454 4019 -12408 4057
rect -12454 3985 -12448 4019
rect -12414 3985 -12408 4019
rect -12454 3947 -12408 3985
rect -12454 3913 -12448 3947
rect -12414 3913 -12408 3947
rect -12454 3875 -12408 3913
rect -12454 3841 -12448 3875
rect -12414 3841 -12408 3875
rect -12454 3803 -12408 3841
rect -12454 3769 -12448 3803
rect -12414 3769 -12408 3803
rect -12454 3731 -12408 3769
rect -12454 3697 -12448 3731
rect -12414 3697 -12408 3731
rect -12454 3659 -12408 3697
rect -12454 3625 -12448 3659
rect -12414 3625 -12408 3659
rect -12454 3587 -12408 3625
rect -12454 3553 -12448 3587
rect -12414 3553 -12408 3587
rect -12454 3515 -12408 3553
rect -12454 3481 -12448 3515
rect -12414 3481 -12408 3515
rect -12454 3466 -12408 3481
rect -12358 4451 -12312 4466
rect -12358 4417 -12352 4451
rect -12318 4417 -12312 4451
rect -12358 4379 -12312 4417
rect -12358 4345 -12352 4379
rect -12318 4345 -12312 4379
rect -12358 4307 -12312 4345
rect -12358 4273 -12352 4307
rect -12318 4273 -12312 4307
rect -12358 4235 -12312 4273
rect -12358 4201 -12352 4235
rect -12318 4201 -12312 4235
rect -12358 4163 -12312 4201
rect -12358 4129 -12352 4163
rect -12318 4129 -12312 4163
rect -12358 4091 -12312 4129
rect -12358 4057 -12352 4091
rect -12318 4057 -12312 4091
rect -12358 4019 -12312 4057
rect -12358 3985 -12352 4019
rect -12318 3985 -12312 4019
rect -12358 3947 -12312 3985
rect -12358 3913 -12352 3947
rect -12318 3913 -12312 3947
rect -12358 3875 -12312 3913
rect -12358 3841 -12352 3875
rect -12318 3841 -12312 3875
rect -12358 3803 -12312 3841
rect -12358 3769 -12352 3803
rect -12318 3769 -12312 3803
rect -12358 3731 -12312 3769
rect -12358 3697 -12352 3731
rect -12318 3697 -12312 3731
rect -12358 3659 -12312 3697
rect -12358 3625 -12352 3659
rect -12318 3625 -12312 3659
rect -12358 3587 -12312 3625
rect -12358 3553 -12352 3587
rect -12318 3553 -12312 3587
rect -12358 3515 -12312 3553
rect -12358 3481 -12352 3515
rect -12318 3481 -12312 3515
rect -12358 3466 -12312 3481
rect -12262 4451 -12216 4466
rect -12262 4417 -12256 4451
rect -12222 4417 -12216 4451
rect -12262 4379 -12216 4417
rect -12262 4345 -12256 4379
rect -12222 4345 -12216 4379
rect -12262 4307 -12216 4345
rect -12262 4273 -12256 4307
rect -12222 4273 -12216 4307
rect -12262 4235 -12216 4273
rect -12262 4201 -12256 4235
rect -12222 4201 -12216 4235
rect -12262 4163 -12216 4201
rect -12262 4129 -12256 4163
rect -12222 4129 -12216 4163
rect -12262 4091 -12216 4129
rect -12262 4057 -12256 4091
rect -12222 4057 -12216 4091
rect -12262 4019 -12216 4057
rect -12262 3985 -12256 4019
rect -12222 3985 -12216 4019
rect -12262 3947 -12216 3985
rect -12262 3913 -12256 3947
rect -12222 3913 -12216 3947
rect -12262 3875 -12216 3913
rect -12262 3841 -12256 3875
rect -12222 3841 -12216 3875
rect -12262 3803 -12216 3841
rect -12262 3769 -12256 3803
rect -12222 3769 -12216 3803
rect -12262 3731 -12216 3769
rect -12262 3697 -12256 3731
rect -12222 3697 -12216 3731
rect -12262 3659 -12216 3697
rect -12262 3625 -12256 3659
rect -12222 3625 -12216 3659
rect -12262 3587 -12216 3625
rect -12262 3553 -12256 3587
rect -12222 3553 -12216 3587
rect -12262 3515 -12216 3553
rect -12262 3481 -12256 3515
rect -12222 3481 -12216 3515
rect -12262 3466 -12216 3481
rect -12166 4451 -12120 4466
rect -12166 4417 -12160 4451
rect -12126 4417 -12120 4451
rect -12166 4379 -12120 4417
rect -12166 4345 -12160 4379
rect -12126 4345 -12120 4379
rect -12166 4307 -12120 4345
rect -12166 4273 -12160 4307
rect -12126 4273 -12120 4307
rect -12166 4235 -12120 4273
rect -12166 4201 -12160 4235
rect -12126 4201 -12120 4235
rect -12166 4163 -12120 4201
rect -12166 4129 -12160 4163
rect -12126 4129 -12120 4163
rect -12166 4091 -12120 4129
rect -12166 4057 -12160 4091
rect -12126 4057 -12120 4091
rect -12166 4019 -12120 4057
rect -12166 3985 -12160 4019
rect -12126 3985 -12120 4019
rect -12166 3947 -12120 3985
rect -12166 3913 -12160 3947
rect -12126 3913 -12120 3947
rect -12166 3875 -12120 3913
rect -12166 3841 -12160 3875
rect -12126 3841 -12120 3875
rect -12166 3803 -12120 3841
rect -12166 3769 -12160 3803
rect -12126 3769 -12120 3803
rect -12166 3731 -12120 3769
rect -12166 3697 -12160 3731
rect -12126 3697 -12120 3731
rect -12166 3659 -12120 3697
rect -12166 3625 -12160 3659
rect -12126 3625 -12120 3659
rect -12166 3587 -12120 3625
rect -12166 3553 -12160 3587
rect -12126 3553 -12120 3587
rect -12166 3515 -12120 3553
rect -12166 3481 -12160 3515
rect -12126 3481 -12120 3515
rect -12166 3466 -12120 3481
rect -12070 4451 -12024 4466
rect -12070 4417 -12064 4451
rect -12030 4417 -12024 4451
rect -12070 4379 -12024 4417
rect -12070 4345 -12064 4379
rect -12030 4345 -12024 4379
rect -12070 4307 -12024 4345
rect -12070 4273 -12064 4307
rect -12030 4273 -12024 4307
rect -12070 4235 -12024 4273
rect -12070 4201 -12064 4235
rect -12030 4201 -12024 4235
rect -12070 4163 -12024 4201
rect -12070 4129 -12064 4163
rect -12030 4129 -12024 4163
rect -12070 4091 -12024 4129
rect -12070 4057 -12064 4091
rect -12030 4057 -12024 4091
rect -12070 4019 -12024 4057
rect -12070 3985 -12064 4019
rect -12030 3985 -12024 4019
rect -12070 3947 -12024 3985
rect -12070 3913 -12064 3947
rect -12030 3913 -12024 3947
rect -12070 3875 -12024 3913
rect -12070 3841 -12064 3875
rect -12030 3841 -12024 3875
rect -12070 3803 -12024 3841
rect -12070 3769 -12064 3803
rect -12030 3769 -12024 3803
rect -12070 3731 -12024 3769
rect -12070 3697 -12064 3731
rect -12030 3697 -12024 3731
rect -12070 3659 -12024 3697
rect -12070 3625 -12064 3659
rect -12030 3625 -12024 3659
rect -12070 3587 -12024 3625
rect -12070 3553 -12064 3587
rect -12030 3553 -12024 3587
rect -12070 3515 -12024 3553
rect -12070 3481 -12064 3515
rect -12030 3481 -12024 3515
rect -12070 3466 -12024 3481
rect -11974 4451 -11928 4466
rect -11974 4417 -11968 4451
rect -11934 4417 -11928 4451
rect -11974 4379 -11928 4417
rect -11974 4345 -11968 4379
rect -11934 4345 -11928 4379
rect -11974 4307 -11928 4345
rect -11974 4273 -11968 4307
rect -11934 4273 -11928 4307
rect -11974 4235 -11928 4273
rect -11974 4201 -11968 4235
rect -11934 4201 -11928 4235
rect -11974 4163 -11928 4201
rect -11974 4129 -11968 4163
rect -11934 4129 -11928 4163
rect -11974 4091 -11928 4129
rect -11974 4057 -11968 4091
rect -11934 4057 -11928 4091
rect -11974 4019 -11928 4057
rect -11974 3985 -11968 4019
rect -11934 3985 -11928 4019
rect -11974 3947 -11928 3985
rect -11974 3913 -11968 3947
rect -11934 3913 -11928 3947
rect -11974 3875 -11928 3913
rect -11974 3841 -11968 3875
rect -11934 3841 -11928 3875
rect -11974 3803 -11928 3841
rect -11974 3769 -11968 3803
rect -11934 3769 -11928 3803
rect -11974 3731 -11928 3769
rect -11974 3697 -11968 3731
rect -11934 3697 -11928 3731
rect -11974 3659 -11928 3697
rect -11974 3625 -11968 3659
rect -11934 3625 -11928 3659
rect -11974 3587 -11928 3625
rect -11974 3553 -11968 3587
rect -11934 3553 -11928 3587
rect -11974 3515 -11928 3553
rect -11974 3481 -11968 3515
rect -11934 3481 -11928 3515
rect -11974 3466 -11928 3481
rect -11766 4453 -11720 4468
rect -11766 4419 -11760 4453
rect -11726 4419 -11720 4453
rect -11766 4381 -11720 4419
rect -11766 4347 -11760 4381
rect -11726 4347 -11720 4381
rect -11766 4309 -11720 4347
rect -11766 4275 -11760 4309
rect -11726 4275 -11720 4309
rect -11766 4237 -11720 4275
rect -11766 4203 -11760 4237
rect -11726 4203 -11720 4237
rect -11766 4165 -11720 4203
rect -11766 4131 -11760 4165
rect -11726 4131 -11720 4165
rect -11766 4093 -11720 4131
rect -11766 4059 -11760 4093
rect -11726 4059 -11720 4093
rect -11766 4021 -11720 4059
rect -11766 3987 -11760 4021
rect -11726 3987 -11720 4021
rect -11766 3949 -11720 3987
rect -11766 3915 -11760 3949
rect -11726 3915 -11720 3949
rect -11766 3877 -11720 3915
rect -11766 3843 -11760 3877
rect -11726 3843 -11720 3877
rect -11766 3805 -11720 3843
rect -11766 3771 -11760 3805
rect -11726 3771 -11720 3805
rect -11766 3733 -11720 3771
rect -11766 3699 -11760 3733
rect -11726 3699 -11720 3733
rect -11766 3661 -11720 3699
rect -11766 3627 -11760 3661
rect -11726 3627 -11720 3661
rect -11766 3589 -11720 3627
rect -11766 3555 -11760 3589
rect -11726 3555 -11720 3589
rect -11766 3517 -11720 3555
rect -11766 3483 -11760 3517
rect -11726 3483 -11720 3517
rect -11766 3468 -11720 3483
rect -11670 4453 -11624 4468
rect -11670 4419 -11664 4453
rect -11630 4419 -11624 4453
rect -11670 4381 -11624 4419
rect -11670 4347 -11664 4381
rect -11630 4347 -11624 4381
rect -11670 4309 -11624 4347
rect -11670 4275 -11664 4309
rect -11630 4275 -11624 4309
rect -11670 4237 -11624 4275
rect -11670 4203 -11664 4237
rect -11630 4203 -11624 4237
rect -11670 4165 -11624 4203
rect -11670 4131 -11664 4165
rect -11630 4131 -11624 4165
rect -11670 4093 -11624 4131
rect -11670 4059 -11664 4093
rect -11630 4059 -11624 4093
rect -11670 4021 -11624 4059
rect -11670 3987 -11664 4021
rect -11630 3987 -11624 4021
rect -11670 3949 -11624 3987
rect -11670 3915 -11664 3949
rect -11630 3915 -11624 3949
rect -11670 3877 -11624 3915
rect -11670 3843 -11664 3877
rect -11630 3843 -11624 3877
rect -11670 3805 -11624 3843
rect -11670 3771 -11664 3805
rect -11630 3771 -11624 3805
rect -11670 3733 -11624 3771
rect -11670 3699 -11664 3733
rect -11630 3699 -11624 3733
rect -11670 3661 -11624 3699
rect -11670 3627 -11664 3661
rect -11630 3627 -11624 3661
rect -11670 3589 -11624 3627
rect -11670 3555 -11664 3589
rect -11630 3555 -11624 3589
rect -11670 3517 -11624 3555
rect -11670 3483 -11664 3517
rect -11630 3483 -11624 3517
rect -11670 3468 -11624 3483
rect -11574 4453 -11528 4468
rect -11574 4419 -11568 4453
rect -11534 4419 -11528 4453
rect -11574 4381 -11528 4419
rect -11574 4347 -11568 4381
rect -11534 4347 -11528 4381
rect -11574 4309 -11528 4347
rect -11574 4275 -11568 4309
rect -11534 4275 -11528 4309
rect -11574 4237 -11528 4275
rect -11574 4203 -11568 4237
rect -11534 4203 -11528 4237
rect -11574 4165 -11528 4203
rect -11574 4131 -11568 4165
rect -11534 4131 -11528 4165
rect -11574 4093 -11528 4131
rect -11574 4059 -11568 4093
rect -11534 4059 -11528 4093
rect -11574 4021 -11528 4059
rect -11574 3987 -11568 4021
rect -11534 3987 -11528 4021
rect -11574 3949 -11528 3987
rect -11574 3915 -11568 3949
rect -11534 3915 -11528 3949
rect -11574 3877 -11528 3915
rect -11574 3843 -11568 3877
rect -11534 3843 -11528 3877
rect -11574 3805 -11528 3843
rect -11574 3771 -11568 3805
rect -11534 3771 -11528 3805
rect -11574 3733 -11528 3771
rect -11574 3699 -11568 3733
rect -11534 3699 -11528 3733
rect -11574 3661 -11528 3699
rect -11574 3627 -11568 3661
rect -11534 3627 -11528 3661
rect -11574 3589 -11528 3627
rect -11574 3555 -11568 3589
rect -11534 3555 -11528 3589
rect -11574 3517 -11528 3555
rect -11574 3483 -11568 3517
rect -11534 3483 -11528 3517
rect -11574 3468 -11528 3483
rect -11478 4453 -11432 4468
rect -11478 4419 -11472 4453
rect -11438 4419 -11432 4453
rect -11478 4381 -11432 4419
rect -11478 4347 -11472 4381
rect -11438 4347 -11432 4381
rect -11478 4309 -11432 4347
rect -11478 4275 -11472 4309
rect -11438 4275 -11432 4309
rect -11478 4237 -11432 4275
rect -11478 4203 -11472 4237
rect -11438 4203 -11432 4237
rect -11478 4165 -11432 4203
rect -11478 4131 -11472 4165
rect -11438 4131 -11432 4165
rect -11478 4093 -11432 4131
rect -11478 4059 -11472 4093
rect -11438 4059 -11432 4093
rect -11478 4021 -11432 4059
rect -11478 3987 -11472 4021
rect -11438 3987 -11432 4021
rect -11478 3949 -11432 3987
rect -11478 3915 -11472 3949
rect -11438 3915 -11432 3949
rect -11478 3877 -11432 3915
rect -11478 3843 -11472 3877
rect -11438 3843 -11432 3877
rect -11478 3805 -11432 3843
rect -11478 3771 -11472 3805
rect -11438 3771 -11432 3805
rect -11478 3733 -11432 3771
rect -11478 3699 -11472 3733
rect -11438 3699 -11432 3733
rect -11478 3661 -11432 3699
rect -11478 3627 -11472 3661
rect -11438 3627 -11432 3661
rect -11478 3589 -11432 3627
rect -11478 3555 -11472 3589
rect -11438 3555 -11432 3589
rect -11478 3517 -11432 3555
rect -11478 3483 -11472 3517
rect -11438 3483 -11432 3517
rect -11478 3468 -11432 3483
rect -11382 4453 -11336 4468
rect -11382 4419 -11376 4453
rect -11342 4419 -11336 4453
rect -11382 4381 -11336 4419
rect -11382 4347 -11376 4381
rect -11342 4347 -11336 4381
rect -11382 4309 -11336 4347
rect -11382 4275 -11376 4309
rect -11342 4275 -11336 4309
rect -11382 4237 -11336 4275
rect -11382 4203 -11376 4237
rect -11342 4203 -11336 4237
rect -11382 4165 -11336 4203
rect -11382 4131 -11376 4165
rect -11342 4131 -11336 4165
rect -11382 4093 -11336 4131
rect -11382 4059 -11376 4093
rect -11342 4059 -11336 4093
rect -11382 4021 -11336 4059
rect -11382 3987 -11376 4021
rect -11342 3987 -11336 4021
rect -11382 3949 -11336 3987
rect -11382 3915 -11376 3949
rect -11342 3915 -11336 3949
rect -11382 3877 -11336 3915
rect -11382 3843 -11376 3877
rect -11342 3843 -11336 3877
rect -11382 3805 -11336 3843
rect -11382 3771 -11376 3805
rect -11342 3771 -11336 3805
rect -11382 3733 -11336 3771
rect -11382 3699 -11376 3733
rect -11342 3699 -11336 3733
rect -11382 3661 -11336 3699
rect -11382 3627 -11376 3661
rect -11342 3627 -11336 3661
rect -11382 3589 -11336 3627
rect -11382 3555 -11376 3589
rect -11342 3555 -11336 3589
rect -11382 3517 -11336 3555
rect -11382 3483 -11376 3517
rect -11342 3483 -11336 3517
rect -11382 3468 -11336 3483
rect -11286 4453 -11240 4468
rect -11286 4419 -11280 4453
rect -11246 4419 -11240 4453
rect -11286 4381 -11240 4419
rect -11286 4347 -11280 4381
rect -11246 4347 -11240 4381
rect -11286 4309 -11240 4347
rect -11286 4275 -11280 4309
rect -11246 4275 -11240 4309
rect -11286 4237 -11240 4275
rect -11286 4203 -11280 4237
rect -11246 4203 -11240 4237
rect -11286 4165 -11240 4203
rect -11286 4131 -11280 4165
rect -11246 4131 -11240 4165
rect -11286 4093 -11240 4131
rect -11286 4059 -11280 4093
rect -11246 4059 -11240 4093
rect -11286 4021 -11240 4059
rect -11286 3987 -11280 4021
rect -11246 3987 -11240 4021
rect -11286 3949 -11240 3987
rect -11286 3915 -11280 3949
rect -11246 3915 -11240 3949
rect -11286 3877 -11240 3915
rect -11286 3843 -11280 3877
rect -11246 3843 -11240 3877
rect -11286 3805 -11240 3843
rect -11286 3771 -11280 3805
rect -11246 3771 -11240 3805
rect -11286 3733 -11240 3771
rect -11286 3699 -11280 3733
rect -11246 3699 -11240 3733
rect -11286 3661 -11240 3699
rect -11286 3627 -11280 3661
rect -11246 3627 -11240 3661
rect -11286 3589 -11240 3627
rect -11286 3555 -11280 3589
rect -11246 3555 -11240 3589
rect -11286 3517 -11240 3555
rect -11286 3483 -11280 3517
rect -11246 3483 -11240 3517
rect -11286 3468 -11240 3483
rect -10296 4437 -10250 4452
rect -10296 4403 -10290 4437
rect -10256 4403 -10250 4437
rect -10296 4365 -10250 4403
rect -10296 4331 -10290 4365
rect -10256 4331 -10250 4365
rect -10296 4293 -10250 4331
rect -10296 4259 -10290 4293
rect -10256 4259 -10250 4293
rect -10296 4221 -10250 4259
rect -10296 4187 -10290 4221
rect -10256 4187 -10250 4221
rect -10296 4149 -10250 4187
rect -10296 4115 -10290 4149
rect -10256 4115 -10250 4149
rect -10296 4077 -10250 4115
rect -10296 4043 -10290 4077
rect -10256 4043 -10250 4077
rect -10296 4005 -10250 4043
rect -10296 3971 -10290 4005
rect -10256 3971 -10250 4005
rect -10296 3933 -10250 3971
rect -10296 3899 -10290 3933
rect -10256 3899 -10250 3933
rect -10296 3861 -10250 3899
rect -10296 3827 -10290 3861
rect -10256 3827 -10250 3861
rect -10296 3789 -10250 3827
rect -10296 3755 -10290 3789
rect -10256 3755 -10250 3789
rect -10296 3717 -10250 3755
rect -10296 3683 -10290 3717
rect -10256 3683 -10250 3717
rect -10296 3645 -10250 3683
rect -10296 3611 -10290 3645
rect -10256 3611 -10250 3645
rect -10296 3573 -10250 3611
rect -10296 3539 -10290 3573
rect -10256 3539 -10250 3573
rect -10296 3501 -10250 3539
rect -10296 3467 -10290 3501
rect -10256 3467 -10250 3501
rect -10296 3452 -10250 3467
rect -10200 4437 -10154 4452
rect -10200 4403 -10194 4437
rect -10160 4403 -10154 4437
rect -10200 4365 -10154 4403
rect -10200 4331 -10194 4365
rect -10160 4331 -10154 4365
rect -10200 4293 -10154 4331
rect -10200 4259 -10194 4293
rect -10160 4259 -10154 4293
rect -10200 4221 -10154 4259
rect -10200 4187 -10194 4221
rect -10160 4187 -10154 4221
rect -10200 4149 -10154 4187
rect -10200 4115 -10194 4149
rect -10160 4115 -10154 4149
rect -10200 4077 -10154 4115
rect -10200 4043 -10194 4077
rect -10160 4043 -10154 4077
rect -10200 4005 -10154 4043
rect -10200 3971 -10194 4005
rect -10160 3971 -10154 4005
rect -10200 3933 -10154 3971
rect -10200 3899 -10194 3933
rect -10160 3899 -10154 3933
rect -10200 3861 -10154 3899
rect -10200 3827 -10194 3861
rect -10160 3827 -10154 3861
rect -10200 3789 -10154 3827
rect -10200 3755 -10194 3789
rect -10160 3755 -10154 3789
rect -10200 3717 -10154 3755
rect -10200 3683 -10194 3717
rect -10160 3683 -10154 3717
rect -10200 3645 -10154 3683
rect -10200 3611 -10194 3645
rect -10160 3611 -10154 3645
rect -10200 3573 -10154 3611
rect -10200 3539 -10194 3573
rect -10160 3539 -10154 3573
rect -10200 3501 -10154 3539
rect -10200 3467 -10194 3501
rect -10160 3467 -10154 3501
rect -10200 3452 -10154 3467
rect -10104 4437 -10058 4452
rect -10104 4403 -10098 4437
rect -10064 4403 -10058 4437
rect -10104 4365 -10058 4403
rect -10104 4331 -10098 4365
rect -10064 4331 -10058 4365
rect -10104 4293 -10058 4331
rect -10104 4259 -10098 4293
rect -10064 4259 -10058 4293
rect -10104 4221 -10058 4259
rect -10104 4187 -10098 4221
rect -10064 4187 -10058 4221
rect -10104 4149 -10058 4187
rect -10104 4115 -10098 4149
rect -10064 4115 -10058 4149
rect -10104 4077 -10058 4115
rect -10104 4043 -10098 4077
rect -10064 4043 -10058 4077
rect -10104 4005 -10058 4043
rect -10104 3971 -10098 4005
rect -10064 3971 -10058 4005
rect -10104 3933 -10058 3971
rect -10104 3899 -10098 3933
rect -10064 3899 -10058 3933
rect -10104 3861 -10058 3899
rect -10104 3827 -10098 3861
rect -10064 3827 -10058 3861
rect -10104 3789 -10058 3827
rect -10104 3755 -10098 3789
rect -10064 3755 -10058 3789
rect -10104 3717 -10058 3755
rect -10104 3683 -10098 3717
rect -10064 3683 -10058 3717
rect -10104 3645 -10058 3683
rect -10104 3611 -10098 3645
rect -10064 3611 -10058 3645
rect -10104 3573 -10058 3611
rect -10104 3539 -10098 3573
rect -10064 3539 -10058 3573
rect -10104 3501 -10058 3539
rect -10104 3467 -10098 3501
rect -10064 3467 -10058 3501
rect -10104 3452 -10058 3467
rect -10008 4437 -9962 4452
rect -10008 4403 -10002 4437
rect -9968 4403 -9962 4437
rect -10008 4365 -9962 4403
rect -10008 4331 -10002 4365
rect -9968 4331 -9962 4365
rect -10008 4293 -9962 4331
rect -10008 4259 -10002 4293
rect -9968 4259 -9962 4293
rect -10008 4221 -9962 4259
rect -10008 4187 -10002 4221
rect -9968 4187 -9962 4221
rect -10008 4149 -9962 4187
rect -10008 4115 -10002 4149
rect -9968 4115 -9962 4149
rect -10008 4077 -9962 4115
rect -10008 4043 -10002 4077
rect -9968 4043 -9962 4077
rect -10008 4005 -9962 4043
rect -10008 3971 -10002 4005
rect -9968 3971 -9962 4005
rect -10008 3933 -9962 3971
rect -10008 3899 -10002 3933
rect -9968 3899 -9962 3933
rect -10008 3861 -9962 3899
rect -10008 3827 -10002 3861
rect -9968 3827 -9962 3861
rect -10008 3789 -9962 3827
rect -10008 3755 -10002 3789
rect -9968 3755 -9962 3789
rect -10008 3717 -9962 3755
rect -10008 3683 -10002 3717
rect -9968 3683 -9962 3717
rect -10008 3645 -9962 3683
rect -10008 3611 -10002 3645
rect -9968 3611 -9962 3645
rect -10008 3573 -9962 3611
rect -10008 3539 -10002 3573
rect -9968 3539 -9962 3573
rect -10008 3501 -9962 3539
rect -10008 3467 -10002 3501
rect -9968 3467 -9962 3501
rect -10008 3452 -9962 3467
rect -9912 4437 -9866 4452
rect -9912 4403 -9906 4437
rect -9872 4403 -9866 4437
rect -9912 4365 -9866 4403
rect -9912 4331 -9906 4365
rect -9872 4331 -9866 4365
rect -9912 4293 -9866 4331
rect -9912 4259 -9906 4293
rect -9872 4259 -9866 4293
rect -9912 4221 -9866 4259
rect -9912 4187 -9906 4221
rect -9872 4187 -9866 4221
rect -9912 4149 -9866 4187
rect -9912 4115 -9906 4149
rect -9872 4115 -9866 4149
rect -9912 4077 -9866 4115
rect -9912 4043 -9906 4077
rect -9872 4043 -9866 4077
rect -9912 4005 -9866 4043
rect -9912 3971 -9906 4005
rect -9872 3971 -9866 4005
rect -9912 3933 -9866 3971
rect -9912 3899 -9906 3933
rect -9872 3899 -9866 3933
rect -9912 3861 -9866 3899
rect -9912 3827 -9906 3861
rect -9872 3827 -9866 3861
rect -9912 3789 -9866 3827
rect -9912 3755 -9906 3789
rect -9872 3755 -9866 3789
rect -9912 3717 -9866 3755
rect -9912 3683 -9906 3717
rect -9872 3683 -9866 3717
rect -9912 3645 -9866 3683
rect -9912 3611 -9906 3645
rect -9872 3611 -9866 3645
rect -9912 3573 -9866 3611
rect -9912 3539 -9906 3573
rect -9872 3539 -9866 3573
rect -9912 3501 -9866 3539
rect -9912 3467 -9906 3501
rect -9872 3467 -9866 3501
rect -9912 3452 -9866 3467
rect -9816 4437 -9770 4452
rect -9816 4403 -9810 4437
rect -9776 4403 -9770 4437
rect -9816 4365 -9770 4403
rect -9816 4331 -9810 4365
rect -9776 4331 -9770 4365
rect -9816 4293 -9770 4331
rect -9816 4259 -9810 4293
rect -9776 4259 -9770 4293
rect -9816 4221 -9770 4259
rect -9816 4187 -9810 4221
rect -9776 4187 -9770 4221
rect -9816 4149 -9770 4187
rect -9816 4115 -9810 4149
rect -9776 4115 -9770 4149
rect -9816 4077 -9770 4115
rect -9816 4043 -9810 4077
rect -9776 4043 -9770 4077
rect -9816 4005 -9770 4043
rect -9816 3971 -9810 4005
rect -9776 3971 -9770 4005
rect -9816 3933 -9770 3971
rect -9816 3899 -9810 3933
rect -9776 3899 -9770 3933
rect -9816 3861 -9770 3899
rect -9816 3827 -9810 3861
rect -9776 3827 -9770 3861
rect -9816 3789 -9770 3827
rect -9816 3755 -9810 3789
rect -9776 3755 -9770 3789
rect -9816 3717 -9770 3755
rect -9816 3683 -9810 3717
rect -9776 3683 -9770 3717
rect -9816 3645 -9770 3683
rect -9816 3611 -9810 3645
rect -9776 3611 -9770 3645
rect -9816 3573 -9770 3611
rect -9816 3539 -9810 3573
rect -9776 3539 -9770 3573
rect -9816 3501 -9770 3539
rect -9816 3467 -9810 3501
rect -9776 3467 -9770 3501
rect -9816 3452 -9770 3467
rect -9720 4437 -9674 4452
rect -9720 4403 -9714 4437
rect -9680 4403 -9674 4437
rect -9720 4365 -9674 4403
rect -9720 4331 -9714 4365
rect -9680 4331 -9674 4365
rect -9720 4293 -9674 4331
rect -9720 4259 -9714 4293
rect -9680 4259 -9674 4293
rect -9720 4221 -9674 4259
rect -9720 4187 -9714 4221
rect -9680 4187 -9674 4221
rect -9720 4149 -9674 4187
rect -9720 4115 -9714 4149
rect -9680 4115 -9674 4149
rect -9720 4077 -9674 4115
rect -9720 4043 -9714 4077
rect -9680 4043 -9674 4077
rect -9720 4005 -9674 4043
rect -9720 3971 -9714 4005
rect -9680 3971 -9674 4005
rect -9720 3933 -9674 3971
rect -9720 3899 -9714 3933
rect -9680 3899 -9674 3933
rect -9720 3861 -9674 3899
rect -9720 3827 -9714 3861
rect -9680 3827 -9674 3861
rect -9720 3789 -9674 3827
rect -9720 3755 -9714 3789
rect -9680 3755 -9674 3789
rect -9720 3717 -9674 3755
rect -9720 3683 -9714 3717
rect -9680 3683 -9674 3717
rect -9720 3645 -9674 3683
rect -9720 3611 -9714 3645
rect -9680 3611 -9674 3645
rect -9720 3573 -9674 3611
rect -9720 3539 -9714 3573
rect -9680 3539 -9674 3573
rect -9720 3501 -9674 3539
rect -9720 3467 -9714 3501
rect -9680 3467 -9674 3501
rect -9720 3452 -9674 3467
rect -9624 4437 -9578 4452
rect -9624 4403 -9618 4437
rect -9584 4403 -9578 4437
rect -9624 4365 -9578 4403
rect -9624 4331 -9618 4365
rect -9584 4331 -9578 4365
rect -9624 4293 -9578 4331
rect -9624 4259 -9618 4293
rect -9584 4259 -9578 4293
rect -9624 4221 -9578 4259
rect -9624 4187 -9618 4221
rect -9584 4187 -9578 4221
rect -9624 4149 -9578 4187
rect -9624 4115 -9618 4149
rect -9584 4115 -9578 4149
rect -9624 4077 -9578 4115
rect -9624 4043 -9618 4077
rect -9584 4043 -9578 4077
rect -9624 4005 -9578 4043
rect -9624 3971 -9618 4005
rect -9584 3971 -9578 4005
rect -9624 3933 -9578 3971
rect -9624 3899 -9618 3933
rect -9584 3899 -9578 3933
rect -9624 3861 -9578 3899
rect -9624 3827 -9618 3861
rect -9584 3827 -9578 3861
rect -9624 3789 -9578 3827
rect -9624 3755 -9618 3789
rect -9584 3755 -9578 3789
rect -9624 3717 -9578 3755
rect -9624 3683 -9618 3717
rect -9584 3683 -9578 3717
rect -9624 3645 -9578 3683
rect -9624 3611 -9618 3645
rect -9584 3611 -9578 3645
rect -9624 3573 -9578 3611
rect -9624 3539 -9618 3573
rect -9584 3539 -9578 3573
rect -9624 3501 -9578 3539
rect -9624 3467 -9618 3501
rect -9584 3467 -9578 3501
rect -9624 3452 -9578 3467
rect -9528 4437 -9482 4452
rect -9528 4403 -9522 4437
rect -9488 4403 -9482 4437
rect -9528 4365 -9482 4403
rect -9528 4331 -9522 4365
rect -9488 4331 -9482 4365
rect -9528 4293 -9482 4331
rect -9528 4259 -9522 4293
rect -9488 4259 -9482 4293
rect -9528 4221 -9482 4259
rect -9528 4187 -9522 4221
rect -9488 4187 -9482 4221
rect -9528 4149 -9482 4187
rect -9528 4115 -9522 4149
rect -9488 4115 -9482 4149
rect -9528 4077 -9482 4115
rect -9528 4043 -9522 4077
rect -9488 4043 -9482 4077
rect -9528 4005 -9482 4043
rect -9528 3971 -9522 4005
rect -9488 3971 -9482 4005
rect -9528 3933 -9482 3971
rect -9528 3899 -9522 3933
rect -9488 3899 -9482 3933
rect -9528 3861 -9482 3899
rect -9528 3827 -9522 3861
rect -9488 3827 -9482 3861
rect -9528 3789 -9482 3827
rect -9528 3755 -9522 3789
rect -9488 3755 -9482 3789
rect -9528 3717 -9482 3755
rect -9528 3683 -9522 3717
rect -9488 3683 -9482 3717
rect -9528 3645 -9482 3683
rect -9528 3611 -9522 3645
rect -9488 3611 -9482 3645
rect -9528 3573 -9482 3611
rect -9528 3539 -9522 3573
rect -9488 3539 -9482 3573
rect -9528 3501 -9482 3539
rect -9528 3467 -9522 3501
rect -9488 3467 -9482 3501
rect -9528 3452 -9482 3467
rect -9432 4437 -9386 4452
rect -9432 4403 -9426 4437
rect -9392 4403 -9386 4437
rect -9432 4365 -9386 4403
rect -9432 4331 -9426 4365
rect -9392 4331 -9386 4365
rect -9432 4293 -9386 4331
rect -9432 4259 -9426 4293
rect -9392 4259 -9386 4293
rect -9432 4221 -9386 4259
rect -9432 4187 -9426 4221
rect -9392 4187 -9386 4221
rect -9432 4149 -9386 4187
rect -9432 4115 -9426 4149
rect -9392 4115 -9386 4149
rect -9432 4077 -9386 4115
rect -9432 4043 -9426 4077
rect -9392 4043 -9386 4077
rect -9432 4005 -9386 4043
rect -9432 3971 -9426 4005
rect -9392 3971 -9386 4005
rect -9432 3933 -9386 3971
rect -9432 3899 -9426 3933
rect -9392 3899 -9386 3933
rect -9432 3861 -9386 3899
rect -9432 3827 -9426 3861
rect -9392 3827 -9386 3861
rect -9432 3789 -9386 3827
rect -9432 3755 -9426 3789
rect -9392 3755 -9386 3789
rect -9432 3717 -9386 3755
rect -9432 3683 -9426 3717
rect -9392 3683 -9386 3717
rect -9432 3645 -9386 3683
rect -9432 3611 -9426 3645
rect -9392 3611 -9386 3645
rect -9432 3573 -9386 3611
rect -9432 3539 -9426 3573
rect -9392 3539 -9386 3573
rect -9432 3501 -9386 3539
rect -9432 3467 -9426 3501
rect -9392 3467 -9386 3501
rect -9432 3452 -9386 3467
rect -9336 4437 -9290 4452
rect -9336 4403 -9330 4437
rect -9296 4403 -9290 4437
rect -9336 4365 -9290 4403
rect -9336 4331 -9330 4365
rect -9296 4331 -9290 4365
rect -9336 4293 -9290 4331
rect -9336 4259 -9330 4293
rect -9296 4259 -9290 4293
rect -9336 4221 -9290 4259
rect -9336 4187 -9330 4221
rect -9296 4187 -9290 4221
rect -9336 4149 -9290 4187
rect -9336 4115 -9330 4149
rect -9296 4115 -9290 4149
rect -9336 4077 -9290 4115
rect -9336 4043 -9330 4077
rect -9296 4043 -9290 4077
rect -9336 4005 -9290 4043
rect -9336 3971 -9330 4005
rect -9296 3971 -9290 4005
rect -9336 3933 -9290 3971
rect -9336 3899 -9330 3933
rect -9296 3899 -9290 3933
rect -9336 3861 -9290 3899
rect -9336 3827 -9330 3861
rect -9296 3827 -9290 3861
rect -9336 3789 -9290 3827
rect -9336 3755 -9330 3789
rect -9296 3755 -9290 3789
rect -9336 3717 -9290 3755
rect -9336 3683 -9330 3717
rect -9296 3683 -9290 3717
rect -9336 3645 -9290 3683
rect -9336 3611 -9330 3645
rect -9296 3611 -9290 3645
rect -9336 3573 -9290 3611
rect -9336 3539 -9330 3573
rect -9296 3539 -9290 3573
rect -9336 3501 -9290 3539
rect -9336 3467 -9330 3501
rect -9296 3467 -9290 3501
rect -9336 3452 -9290 3467
rect -9240 4437 -9194 4452
rect -9240 4403 -9234 4437
rect -9200 4403 -9194 4437
rect -9240 4365 -9194 4403
rect -9240 4331 -9234 4365
rect -9200 4331 -9194 4365
rect -9240 4293 -9194 4331
rect -9240 4259 -9234 4293
rect -9200 4259 -9194 4293
rect -9240 4221 -9194 4259
rect -9240 4187 -9234 4221
rect -9200 4187 -9194 4221
rect -9240 4149 -9194 4187
rect -9240 4115 -9234 4149
rect -9200 4115 -9194 4149
rect -9240 4077 -9194 4115
rect -9240 4043 -9234 4077
rect -9200 4043 -9194 4077
rect -9240 4005 -9194 4043
rect -9240 3971 -9234 4005
rect -9200 3971 -9194 4005
rect -9240 3933 -9194 3971
rect -9240 3899 -9234 3933
rect -9200 3899 -9194 3933
rect -9240 3861 -9194 3899
rect -9240 3827 -9234 3861
rect -9200 3827 -9194 3861
rect -9240 3789 -9194 3827
rect -9240 3755 -9234 3789
rect -9200 3755 -9194 3789
rect -9240 3717 -9194 3755
rect -9240 3683 -9234 3717
rect -9200 3683 -9194 3717
rect -9240 3645 -9194 3683
rect -9240 3611 -9234 3645
rect -9200 3611 -9194 3645
rect -9240 3573 -9194 3611
rect -9240 3539 -9234 3573
rect -9200 3539 -9194 3573
rect -9240 3501 -9194 3539
rect -9240 3467 -9234 3501
rect -9200 3467 -9194 3501
rect -9240 3452 -9194 3467
rect -9144 4437 -9098 4452
rect -9144 4403 -9138 4437
rect -9104 4403 -9098 4437
rect -9144 4365 -9098 4403
rect -9144 4331 -9138 4365
rect -9104 4331 -9098 4365
rect -9144 4293 -9098 4331
rect -9144 4259 -9138 4293
rect -9104 4259 -9098 4293
rect -9144 4221 -9098 4259
rect -9144 4187 -9138 4221
rect -9104 4187 -9098 4221
rect -9144 4149 -9098 4187
rect -9144 4115 -9138 4149
rect -9104 4115 -9098 4149
rect -9144 4077 -9098 4115
rect -9144 4043 -9138 4077
rect -9104 4043 -9098 4077
rect -9144 4005 -9098 4043
rect -9144 3971 -9138 4005
rect -9104 3971 -9098 4005
rect -9144 3933 -9098 3971
rect -9144 3899 -9138 3933
rect -9104 3899 -9098 3933
rect -9144 3861 -9098 3899
rect -9144 3827 -9138 3861
rect -9104 3827 -9098 3861
rect -9144 3789 -9098 3827
rect -9144 3755 -9138 3789
rect -9104 3755 -9098 3789
rect -9144 3717 -9098 3755
rect -9144 3683 -9138 3717
rect -9104 3683 -9098 3717
rect -9144 3645 -9098 3683
rect -9144 3611 -9138 3645
rect -9104 3611 -9098 3645
rect -9144 3573 -9098 3611
rect -9144 3539 -9138 3573
rect -9104 3539 -9098 3573
rect -9144 3501 -9098 3539
rect -9144 3467 -9138 3501
rect -9104 3467 -9098 3501
rect -9144 3452 -9098 3467
rect -9048 4437 -9002 4452
rect -9048 4403 -9042 4437
rect -9008 4403 -9002 4437
rect -9048 4365 -9002 4403
rect -9048 4331 -9042 4365
rect -9008 4331 -9002 4365
rect -9048 4293 -9002 4331
rect -9048 4259 -9042 4293
rect -9008 4259 -9002 4293
rect -9048 4221 -9002 4259
rect -9048 4187 -9042 4221
rect -9008 4187 -9002 4221
rect -9048 4149 -9002 4187
rect -9048 4115 -9042 4149
rect -9008 4115 -9002 4149
rect -9048 4077 -9002 4115
rect -9048 4043 -9042 4077
rect -9008 4043 -9002 4077
rect -9048 4005 -9002 4043
rect -9048 3971 -9042 4005
rect -9008 3971 -9002 4005
rect -9048 3933 -9002 3971
rect -9048 3899 -9042 3933
rect -9008 3899 -9002 3933
rect -9048 3861 -9002 3899
rect -9048 3827 -9042 3861
rect -9008 3827 -9002 3861
rect -9048 3789 -9002 3827
rect -9048 3755 -9042 3789
rect -9008 3755 -9002 3789
rect -9048 3717 -9002 3755
rect -9048 3683 -9042 3717
rect -9008 3683 -9002 3717
rect -9048 3645 -9002 3683
rect -9048 3611 -9042 3645
rect -9008 3611 -9002 3645
rect -9048 3573 -9002 3611
rect -9048 3539 -9042 3573
rect -9008 3539 -9002 3573
rect -9048 3501 -9002 3539
rect -9048 3467 -9042 3501
rect -9008 3467 -9002 3501
rect -9048 3452 -9002 3467
rect -8952 4437 -8906 4452
rect -8952 4403 -8946 4437
rect -8912 4403 -8906 4437
rect -8952 4365 -8906 4403
rect -8952 4331 -8946 4365
rect -8912 4331 -8906 4365
rect -8952 4293 -8906 4331
rect -8952 4259 -8946 4293
rect -8912 4259 -8906 4293
rect -8952 4221 -8906 4259
rect -8952 4187 -8946 4221
rect -8912 4187 -8906 4221
rect -8952 4149 -8906 4187
rect -8952 4115 -8946 4149
rect -8912 4115 -8906 4149
rect -8952 4077 -8906 4115
rect -8952 4043 -8946 4077
rect -8912 4043 -8906 4077
rect -8952 4005 -8906 4043
rect -8952 3971 -8946 4005
rect -8912 3971 -8906 4005
rect -8952 3933 -8906 3971
rect -8952 3899 -8946 3933
rect -8912 3899 -8906 3933
rect -8952 3861 -8906 3899
rect -8952 3827 -8946 3861
rect -8912 3827 -8906 3861
rect -8952 3789 -8906 3827
rect -8952 3755 -8946 3789
rect -8912 3755 -8906 3789
rect -8952 3717 -8906 3755
rect -8952 3683 -8946 3717
rect -8912 3683 -8906 3717
rect -8952 3645 -8906 3683
rect -8952 3611 -8946 3645
rect -8912 3611 -8906 3645
rect -8952 3573 -8906 3611
rect -8952 3539 -8946 3573
rect -8912 3539 -8906 3573
rect -8952 3501 -8906 3539
rect -8952 3467 -8946 3501
rect -8912 3467 -8906 3501
rect -8952 3452 -8906 3467
rect -8856 4437 -8810 4452
rect -8856 4403 -8850 4437
rect -8816 4403 -8810 4437
rect -8856 4365 -8810 4403
rect -8856 4331 -8850 4365
rect -8816 4331 -8810 4365
rect -8856 4293 -8810 4331
rect -8856 4259 -8850 4293
rect -8816 4259 -8810 4293
rect -8856 4221 -8810 4259
rect -8856 4187 -8850 4221
rect -8816 4187 -8810 4221
rect -8856 4149 -8810 4187
rect -8856 4115 -8850 4149
rect -8816 4115 -8810 4149
rect -8856 4077 -8810 4115
rect -8856 4043 -8850 4077
rect -8816 4043 -8810 4077
rect -8856 4005 -8810 4043
rect -8856 3971 -8850 4005
rect -8816 3971 -8810 4005
rect -8856 3933 -8810 3971
rect -8856 3899 -8850 3933
rect -8816 3899 -8810 3933
rect -8856 3861 -8810 3899
rect -8856 3827 -8850 3861
rect -8816 3827 -8810 3861
rect -8856 3789 -8810 3827
rect -8856 3755 -8850 3789
rect -8816 3755 -8810 3789
rect -8856 3717 -8810 3755
rect -8856 3683 -8850 3717
rect -8816 3683 -8810 3717
rect -8856 3645 -8810 3683
rect -8856 3611 -8850 3645
rect -8816 3611 -8810 3645
rect -8856 3573 -8810 3611
rect -8856 3539 -8850 3573
rect -8816 3539 -8810 3573
rect -8856 3501 -8810 3539
rect -8856 3467 -8850 3501
rect -8816 3467 -8810 3501
rect -8856 3452 -8810 3467
rect -8760 4437 -8714 4452
rect -8760 4403 -8754 4437
rect -8720 4403 -8714 4437
rect -8760 4365 -8714 4403
rect -8760 4331 -8754 4365
rect -8720 4331 -8714 4365
rect -8760 4293 -8714 4331
rect -8760 4259 -8754 4293
rect -8720 4259 -8714 4293
rect -8760 4221 -8714 4259
rect -8760 4187 -8754 4221
rect -8720 4187 -8714 4221
rect -8760 4149 -8714 4187
rect -8760 4115 -8754 4149
rect -8720 4115 -8714 4149
rect -8760 4077 -8714 4115
rect -8760 4043 -8754 4077
rect -8720 4043 -8714 4077
rect -8760 4005 -8714 4043
rect -8760 3971 -8754 4005
rect -8720 3971 -8714 4005
rect -8760 3933 -8714 3971
rect -8760 3899 -8754 3933
rect -8720 3899 -8714 3933
rect -8760 3861 -8714 3899
rect -8760 3827 -8754 3861
rect -8720 3827 -8714 3861
rect -8760 3789 -8714 3827
rect -8760 3755 -8754 3789
rect -8720 3755 -8714 3789
rect -8760 3717 -8714 3755
rect -8760 3683 -8754 3717
rect -8720 3683 -8714 3717
rect -8760 3645 -8714 3683
rect -8760 3611 -8754 3645
rect -8720 3611 -8714 3645
rect -8760 3573 -8714 3611
rect -8760 3539 -8754 3573
rect -8720 3539 -8714 3573
rect -8760 3501 -8714 3539
rect -8760 3467 -8754 3501
rect -8720 3467 -8714 3501
rect -8760 3452 -8714 3467
rect -8664 4437 -8618 4452
rect -8664 4403 -8658 4437
rect -8624 4403 -8618 4437
rect -8664 4365 -8618 4403
rect -8664 4331 -8658 4365
rect -8624 4331 -8618 4365
rect -8664 4293 -8618 4331
rect -8664 4259 -8658 4293
rect -8624 4259 -8618 4293
rect -8664 4221 -8618 4259
rect -8664 4187 -8658 4221
rect -8624 4187 -8618 4221
rect -8664 4149 -8618 4187
rect -8664 4115 -8658 4149
rect -8624 4115 -8618 4149
rect -8664 4077 -8618 4115
rect -8664 4043 -8658 4077
rect -8624 4043 -8618 4077
rect -8664 4005 -8618 4043
rect -8664 3971 -8658 4005
rect -8624 3971 -8618 4005
rect -8664 3933 -8618 3971
rect -8664 3899 -8658 3933
rect -8624 3899 -8618 3933
rect -8664 3861 -8618 3899
rect -8664 3827 -8658 3861
rect -8624 3827 -8618 3861
rect -8664 3789 -8618 3827
rect -8664 3755 -8658 3789
rect -8624 3755 -8618 3789
rect -8664 3717 -8618 3755
rect -8664 3683 -8658 3717
rect -8624 3683 -8618 3717
rect -8664 3645 -8618 3683
rect -8664 3611 -8658 3645
rect -8624 3611 -8618 3645
rect -8664 3573 -8618 3611
rect -8664 3539 -8658 3573
rect -8624 3539 -8618 3573
rect -8664 3501 -8618 3539
rect -8664 3467 -8658 3501
rect -8624 3467 -8618 3501
rect -8664 3452 -8618 3467
rect -8568 4437 -8522 4452
rect -8568 4403 -8562 4437
rect -8528 4403 -8522 4437
rect -8568 4365 -8522 4403
rect -8568 4331 -8562 4365
rect -8528 4331 -8522 4365
rect -8568 4293 -8522 4331
rect -8568 4259 -8562 4293
rect -8528 4259 -8522 4293
rect -8568 4221 -8522 4259
rect -8568 4187 -8562 4221
rect -8528 4187 -8522 4221
rect -8568 4149 -8522 4187
rect -8568 4115 -8562 4149
rect -8528 4115 -8522 4149
rect -8568 4077 -8522 4115
rect -8568 4043 -8562 4077
rect -8528 4043 -8522 4077
rect -8568 4005 -8522 4043
rect -8568 3971 -8562 4005
rect -8528 3971 -8522 4005
rect -8568 3933 -8522 3971
rect -8568 3899 -8562 3933
rect -8528 3899 -8522 3933
rect -8568 3861 -8522 3899
rect -8568 3827 -8562 3861
rect -8528 3827 -8522 3861
rect -8568 3789 -8522 3827
rect -8568 3755 -8562 3789
rect -8528 3755 -8522 3789
rect -8568 3717 -8522 3755
rect -8568 3683 -8562 3717
rect -8528 3683 -8522 3717
rect -8568 3645 -8522 3683
rect -8568 3611 -8562 3645
rect -8528 3611 -8522 3645
rect -8568 3573 -8522 3611
rect -8568 3539 -8562 3573
rect -8528 3539 -8522 3573
rect -8568 3501 -8522 3539
rect -8568 3467 -8562 3501
rect -8528 3467 -8522 3501
rect -8568 3452 -8522 3467
rect -8472 4437 -8426 4452
rect -8472 4403 -8466 4437
rect -8432 4403 -8426 4437
rect -8472 4365 -8426 4403
rect -8472 4331 -8466 4365
rect -8432 4331 -8426 4365
rect -8472 4293 -8426 4331
rect -8472 4259 -8466 4293
rect -8432 4259 -8426 4293
rect -8472 4221 -8426 4259
rect -8472 4187 -8466 4221
rect -8432 4187 -8426 4221
rect -8472 4149 -8426 4187
rect -8472 4115 -8466 4149
rect -8432 4115 -8426 4149
rect -8472 4077 -8426 4115
rect -8472 4043 -8466 4077
rect -8432 4043 -8426 4077
rect -8472 4005 -8426 4043
rect -8472 3971 -8466 4005
rect -8432 3971 -8426 4005
rect -8472 3933 -8426 3971
rect -8472 3899 -8466 3933
rect -8432 3899 -8426 3933
rect -8472 3861 -8426 3899
rect -8472 3827 -8466 3861
rect -8432 3827 -8426 3861
rect -8472 3789 -8426 3827
rect -8472 3755 -8466 3789
rect -8432 3755 -8426 3789
rect -8472 3717 -8426 3755
rect -8472 3683 -8466 3717
rect -8432 3683 -8426 3717
rect -8472 3645 -8426 3683
rect -8472 3611 -8466 3645
rect -8432 3611 -8426 3645
rect -8472 3573 -8426 3611
rect -8472 3539 -8466 3573
rect -8432 3539 -8426 3573
rect -8472 3501 -8426 3539
rect -8472 3467 -8466 3501
rect -8432 3467 -8426 3501
rect -8472 3452 -8426 3467
rect -8376 4437 -8330 4452
rect -8376 4403 -8370 4437
rect -8336 4403 -8330 4437
rect -8376 4365 -8330 4403
rect -8376 4331 -8370 4365
rect -8336 4331 -8330 4365
rect -8376 4293 -8330 4331
rect -8376 4259 -8370 4293
rect -8336 4259 -8330 4293
rect -8376 4221 -8330 4259
rect -8376 4187 -8370 4221
rect -8336 4187 -8330 4221
rect -8376 4149 -8330 4187
rect -8376 4115 -8370 4149
rect -8336 4115 -8330 4149
rect -8376 4077 -8330 4115
rect -8376 4043 -8370 4077
rect -8336 4043 -8330 4077
rect -8376 4005 -8330 4043
rect -8376 3971 -8370 4005
rect -8336 3971 -8330 4005
rect -8376 3933 -8330 3971
rect -8376 3899 -8370 3933
rect -8336 3899 -8330 3933
rect -8376 3861 -8330 3899
rect -8376 3827 -8370 3861
rect -8336 3827 -8330 3861
rect -8376 3789 -8330 3827
rect -8376 3755 -8370 3789
rect -8336 3755 -8330 3789
rect -8376 3717 -8330 3755
rect -8376 3683 -8370 3717
rect -8336 3683 -8330 3717
rect -8376 3645 -8330 3683
rect -8376 3611 -8370 3645
rect -8336 3611 -8330 3645
rect -8376 3573 -8330 3611
rect -8376 3539 -8370 3573
rect -8336 3539 -8330 3573
rect -8376 3501 -8330 3539
rect -8376 3467 -8370 3501
rect -8336 3467 -8330 3501
rect -8376 3452 -8330 3467
rect -8152 4443 -8106 4458
rect -8152 4409 -8146 4443
rect -8112 4409 -8106 4443
rect -8152 4371 -8106 4409
rect -8152 4337 -8146 4371
rect -8112 4337 -8106 4371
rect -8152 4299 -8106 4337
rect -8152 4265 -8146 4299
rect -8112 4265 -8106 4299
rect -8152 4227 -8106 4265
rect -8152 4193 -8146 4227
rect -8112 4193 -8106 4227
rect -8152 4155 -8106 4193
rect -8152 4121 -8146 4155
rect -8112 4121 -8106 4155
rect -8152 4083 -8106 4121
rect -8152 4049 -8146 4083
rect -8112 4049 -8106 4083
rect -8152 4011 -8106 4049
rect -8152 3977 -8146 4011
rect -8112 3977 -8106 4011
rect -8152 3939 -8106 3977
rect -8152 3905 -8146 3939
rect -8112 3905 -8106 3939
rect -8152 3867 -8106 3905
rect -8152 3833 -8146 3867
rect -8112 3833 -8106 3867
rect -8152 3795 -8106 3833
rect -8152 3761 -8146 3795
rect -8112 3761 -8106 3795
rect -8152 3723 -8106 3761
rect -8152 3689 -8146 3723
rect -8112 3689 -8106 3723
rect -8152 3651 -8106 3689
rect -8152 3617 -8146 3651
rect -8112 3617 -8106 3651
rect -8152 3579 -8106 3617
rect -8152 3545 -8146 3579
rect -8112 3545 -8106 3579
rect -8152 3507 -8106 3545
rect -8152 3473 -8146 3507
rect -8112 3473 -8106 3507
rect -8152 3458 -8106 3473
rect -8056 4443 -8010 4458
rect -8056 4409 -8050 4443
rect -8016 4409 -8010 4443
rect -8056 4371 -8010 4409
rect -8056 4337 -8050 4371
rect -8016 4337 -8010 4371
rect -8056 4299 -8010 4337
rect -8056 4265 -8050 4299
rect -8016 4265 -8010 4299
rect -8056 4227 -8010 4265
rect -8056 4193 -8050 4227
rect -8016 4193 -8010 4227
rect -8056 4155 -8010 4193
rect -8056 4121 -8050 4155
rect -8016 4121 -8010 4155
rect -8056 4083 -8010 4121
rect -8056 4049 -8050 4083
rect -8016 4049 -8010 4083
rect -8056 4011 -8010 4049
rect -8056 3977 -8050 4011
rect -8016 3977 -8010 4011
rect -8056 3939 -8010 3977
rect -8056 3905 -8050 3939
rect -8016 3905 -8010 3939
rect -8056 3867 -8010 3905
rect -8056 3833 -8050 3867
rect -8016 3833 -8010 3867
rect -8056 3795 -8010 3833
rect -8056 3761 -8050 3795
rect -8016 3761 -8010 3795
rect -8056 3723 -8010 3761
rect -8056 3689 -8050 3723
rect -8016 3689 -8010 3723
rect -8056 3651 -8010 3689
rect -8056 3617 -8050 3651
rect -8016 3617 -8010 3651
rect -8056 3579 -8010 3617
rect -8056 3545 -8050 3579
rect -8016 3545 -8010 3579
rect -8056 3507 -8010 3545
rect -8056 3473 -8050 3507
rect -8016 3473 -8010 3507
rect -8056 3458 -8010 3473
rect -7960 4443 -7914 4458
rect -7960 4409 -7954 4443
rect -7920 4409 -7914 4443
rect -7960 4371 -7914 4409
rect -7960 4337 -7954 4371
rect -7920 4337 -7914 4371
rect -7960 4299 -7914 4337
rect -7960 4265 -7954 4299
rect -7920 4265 -7914 4299
rect -7960 4227 -7914 4265
rect -7960 4193 -7954 4227
rect -7920 4193 -7914 4227
rect -7960 4155 -7914 4193
rect -7960 4121 -7954 4155
rect -7920 4121 -7914 4155
rect -7960 4083 -7914 4121
rect -7960 4049 -7954 4083
rect -7920 4049 -7914 4083
rect -7960 4011 -7914 4049
rect -7960 3977 -7954 4011
rect -7920 3977 -7914 4011
rect -7960 3939 -7914 3977
rect -7960 3905 -7954 3939
rect -7920 3905 -7914 3939
rect -7960 3867 -7914 3905
rect -7960 3833 -7954 3867
rect -7920 3833 -7914 3867
rect -7960 3795 -7914 3833
rect -7960 3761 -7954 3795
rect -7920 3761 -7914 3795
rect -7960 3723 -7914 3761
rect -7960 3689 -7954 3723
rect -7920 3689 -7914 3723
rect -7960 3651 -7914 3689
rect -7960 3617 -7954 3651
rect -7920 3617 -7914 3651
rect -7960 3579 -7914 3617
rect -7960 3545 -7954 3579
rect -7920 3545 -7914 3579
rect -7960 3507 -7914 3545
rect -7960 3473 -7954 3507
rect -7920 3473 -7914 3507
rect -7960 3458 -7914 3473
rect -7864 4443 -7818 4458
rect -7864 4409 -7858 4443
rect -7824 4409 -7818 4443
rect -7864 4371 -7818 4409
rect -7864 4337 -7858 4371
rect -7824 4337 -7818 4371
rect -7864 4299 -7818 4337
rect -7864 4265 -7858 4299
rect -7824 4265 -7818 4299
rect -7864 4227 -7818 4265
rect -7864 4193 -7858 4227
rect -7824 4193 -7818 4227
rect -7864 4155 -7818 4193
rect -7864 4121 -7858 4155
rect -7824 4121 -7818 4155
rect -7864 4083 -7818 4121
rect -7864 4049 -7858 4083
rect -7824 4049 -7818 4083
rect -7864 4011 -7818 4049
rect -7864 3977 -7858 4011
rect -7824 3977 -7818 4011
rect -7864 3939 -7818 3977
rect -7864 3905 -7858 3939
rect -7824 3905 -7818 3939
rect -7864 3867 -7818 3905
rect -7864 3833 -7858 3867
rect -7824 3833 -7818 3867
rect -7864 3795 -7818 3833
rect -7864 3761 -7858 3795
rect -7824 3761 -7818 3795
rect -7864 3723 -7818 3761
rect -7864 3689 -7858 3723
rect -7824 3689 -7818 3723
rect -7864 3651 -7818 3689
rect -7864 3617 -7858 3651
rect -7824 3617 -7818 3651
rect -7864 3579 -7818 3617
rect -7864 3545 -7858 3579
rect -7824 3545 -7818 3579
rect -7864 3507 -7818 3545
rect -7864 3473 -7858 3507
rect -7824 3473 -7818 3507
rect -7864 3458 -7818 3473
rect -7768 4443 -7722 4458
rect -7768 4409 -7762 4443
rect -7728 4409 -7722 4443
rect -7768 4371 -7722 4409
rect -7768 4337 -7762 4371
rect -7728 4337 -7722 4371
rect -7768 4299 -7722 4337
rect -7768 4265 -7762 4299
rect -7728 4265 -7722 4299
rect -7768 4227 -7722 4265
rect -7768 4193 -7762 4227
rect -7728 4193 -7722 4227
rect -7768 4155 -7722 4193
rect -7768 4121 -7762 4155
rect -7728 4121 -7722 4155
rect -7768 4083 -7722 4121
rect -7768 4049 -7762 4083
rect -7728 4049 -7722 4083
rect -7768 4011 -7722 4049
rect -7768 3977 -7762 4011
rect -7728 3977 -7722 4011
rect -7768 3939 -7722 3977
rect -7768 3905 -7762 3939
rect -7728 3905 -7722 3939
rect -7768 3867 -7722 3905
rect -7768 3833 -7762 3867
rect -7728 3833 -7722 3867
rect -7768 3795 -7722 3833
rect -7768 3761 -7762 3795
rect -7728 3761 -7722 3795
rect -7768 3723 -7722 3761
rect -7768 3689 -7762 3723
rect -7728 3689 -7722 3723
rect -7768 3651 -7722 3689
rect -7768 3617 -7762 3651
rect -7728 3617 -7722 3651
rect -7768 3579 -7722 3617
rect -7768 3545 -7762 3579
rect -7728 3545 -7722 3579
rect -7768 3507 -7722 3545
rect -7768 3473 -7762 3507
rect -7728 3473 -7722 3507
rect -7768 3458 -7722 3473
rect -7672 4443 -7626 4458
rect -7672 4409 -7666 4443
rect -7632 4409 -7626 4443
rect -7672 4371 -7626 4409
rect -7672 4337 -7666 4371
rect -7632 4337 -7626 4371
rect -7672 4299 -7626 4337
rect -7672 4265 -7666 4299
rect -7632 4265 -7626 4299
rect -7672 4227 -7626 4265
rect -7672 4193 -7666 4227
rect -7632 4193 -7626 4227
rect -7672 4155 -7626 4193
rect -7672 4121 -7666 4155
rect -7632 4121 -7626 4155
rect -7672 4083 -7626 4121
rect -7672 4049 -7666 4083
rect -7632 4049 -7626 4083
rect -7672 4011 -7626 4049
rect -7672 3977 -7666 4011
rect -7632 3977 -7626 4011
rect -7672 3939 -7626 3977
rect -7672 3905 -7666 3939
rect -7632 3905 -7626 3939
rect -7672 3867 -7626 3905
rect -7672 3833 -7666 3867
rect -7632 3833 -7626 3867
rect -7672 3795 -7626 3833
rect -7672 3761 -7666 3795
rect -7632 3761 -7626 3795
rect -7672 3723 -7626 3761
rect -7672 3689 -7666 3723
rect -7632 3689 -7626 3723
rect -7672 3651 -7626 3689
rect -7672 3617 -7666 3651
rect -7632 3617 -7626 3651
rect -7672 3579 -7626 3617
rect -7672 3545 -7666 3579
rect -7632 3545 -7626 3579
rect -7672 3507 -7626 3545
rect -7672 3473 -7666 3507
rect -7632 3473 -7626 3507
rect -7672 3458 -7626 3473
rect -7576 4443 -7530 4458
rect -7576 4409 -7570 4443
rect -7536 4409 -7530 4443
rect -7576 4371 -7530 4409
rect -7576 4337 -7570 4371
rect -7536 4337 -7530 4371
rect -7576 4299 -7530 4337
rect -7576 4265 -7570 4299
rect -7536 4265 -7530 4299
rect -7576 4227 -7530 4265
rect -7576 4193 -7570 4227
rect -7536 4193 -7530 4227
rect -7576 4155 -7530 4193
rect -7576 4121 -7570 4155
rect -7536 4121 -7530 4155
rect -7576 4083 -7530 4121
rect -7576 4049 -7570 4083
rect -7536 4049 -7530 4083
rect -7576 4011 -7530 4049
rect -7576 3977 -7570 4011
rect -7536 3977 -7530 4011
rect -7576 3939 -7530 3977
rect -7576 3905 -7570 3939
rect -7536 3905 -7530 3939
rect -7576 3867 -7530 3905
rect -7576 3833 -7570 3867
rect -7536 3833 -7530 3867
rect -7576 3795 -7530 3833
rect -7576 3761 -7570 3795
rect -7536 3761 -7530 3795
rect -7576 3723 -7530 3761
rect -7576 3689 -7570 3723
rect -7536 3689 -7530 3723
rect -7576 3651 -7530 3689
rect -7576 3617 -7570 3651
rect -7536 3617 -7530 3651
rect -7576 3579 -7530 3617
rect -7576 3545 -7570 3579
rect -7536 3545 -7530 3579
rect -7576 3507 -7530 3545
rect -7576 3473 -7570 3507
rect -7536 3473 -7530 3507
rect -7576 3458 -7530 3473
rect -7480 4443 -7434 4458
rect -7480 4409 -7474 4443
rect -7440 4409 -7434 4443
rect -7480 4371 -7434 4409
rect -7480 4337 -7474 4371
rect -7440 4337 -7434 4371
rect -7480 4299 -7434 4337
rect -7480 4265 -7474 4299
rect -7440 4265 -7434 4299
rect -7480 4227 -7434 4265
rect -7480 4193 -7474 4227
rect -7440 4193 -7434 4227
rect -7480 4155 -7434 4193
rect -7480 4121 -7474 4155
rect -7440 4121 -7434 4155
rect -7480 4083 -7434 4121
rect -7480 4049 -7474 4083
rect -7440 4049 -7434 4083
rect -7480 4011 -7434 4049
rect -7480 3977 -7474 4011
rect -7440 3977 -7434 4011
rect -7480 3939 -7434 3977
rect -7480 3905 -7474 3939
rect -7440 3905 -7434 3939
rect -7480 3867 -7434 3905
rect -7480 3833 -7474 3867
rect -7440 3833 -7434 3867
rect -7480 3795 -7434 3833
rect -7480 3761 -7474 3795
rect -7440 3761 -7434 3795
rect -7480 3723 -7434 3761
rect -7480 3689 -7474 3723
rect -7440 3689 -7434 3723
rect -7480 3651 -7434 3689
rect -7480 3617 -7474 3651
rect -7440 3617 -7434 3651
rect -7480 3579 -7434 3617
rect -7480 3545 -7474 3579
rect -7440 3545 -7434 3579
rect -7480 3507 -7434 3545
rect -7480 3473 -7474 3507
rect -7440 3473 -7434 3507
rect -7480 3458 -7434 3473
rect -7384 4443 -7338 4458
rect -7384 4409 -7378 4443
rect -7344 4409 -7338 4443
rect -7384 4371 -7338 4409
rect -7384 4337 -7378 4371
rect -7344 4337 -7338 4371
rect -7384 4299 -7338 4337
rect -7384 4265 -7378 4299
rect -7344 4265 -7338 4299
rect -7384 4227 -7338 4265
rect -7384 4193 -7378 4227
rect -7344 4193 -7338 4227
rect -7384 4155 -7338 4193
rect -7384 4121 -7378 4155
rect -7344 4121 -7338 4155
rect -7384 4083 -7338 4121
rect -7384 4049 -7378 4083
rect -7344 4049 -7338 4083
rect -7384 4011 -7338 4049
rect -7384 3977 -7378 4011
rect -7344 3977 -7338 4011
rect -7384 3939 -7338 3977
rect -7384 3905 -7378 3939
rect -7344 3905 -7338 3939
rect -7384 3867 -7338 3905
rect -7384 3833 -7378 3867
rect -7344 3833 -7338 3867
rect -7384 3795 -7338 3833
rect -7384 3761 -7378 3795
rect -7344 3761 -7338 3795
rect -7384 3723 -7338 3761
rect -7384 3689 -7378 3723
rect -7344 3689 -7338 3723
rect -7384 3651 -7338 3689
rect -7384 3617 -7378 3651
rect -7344 3617 -7338 3651
rect -7384 3579 -7338 3617
rect -7384 3545 -7378 3579
rect -7344 3545 -7338 3579
rect -7384 3507 -7338 3545
rect -7384 3473 -7378 3507
rect -7344 3473 -7338 3507
rect -7384 3458 -7338 3473
rect -7288 4443 -7242 4458
rect -7288 4409 -7282 4443
rect -7248 4409 -7242 4443
rect -7288 4371 -7242 4409
rect -7288 4337 -7282 4371
rect -7248 4337 -7242 4371
rect -7288 4299 -7242 4337
rect -7288 4265 -7282 4299
rect -7248 4265 -7242 4299
rect -7288 4227 -7242 4265
rect -7288 4193 -7282 4227
rect -7248 4193 -7242 4227
rect -7288 4155 -7242 4193
rect -7288 4121 -7282 4155
rect -7248 4121 -7242 4155
rect -7288 4083 -7242 4121
rect -7288 4049 -7282 4083
rect -7248 4049 -7242 4083
rect -7288 4011 -7242 4049
rect -7288 3977 -7282 4011
rect -7248 3977 -7242 4011
rect -7288 3939 -7242 3977
rect -7288 3905 -7282 3939
rect -7248 3905 -7242 3939
rect -7288 3867 -7242 3905
rect -7288 3833 -7282 3867
rect -7248 3833 -7242 3867
rect -7288 3795 -7242 3833
rect -7288 3761 -7282 3795
rect -7248 3761 -7242 3795
rect -7288 3723 -7242 3761
rect -7288 3689 -7282 3723
rect -7248 3689 -7242 3723
rect -7288 3651 -7242 3689
rect -7288 3617 -7282 3651
rect -7248 3617 -7242 3651
rect -7288 3579 -7242 3617
rect -7288 3545 -7282 3579
rect -7248 3545 -7242 3579
rect -7288 3507 -7242 3545
rect -7288 3473 -7282 3507
rect -7248 3473 -7242 3507
rect -7288 3458 -7242 3473
rect -7192 4443 -7146 4458
rect -7192 4409 -7186 4443
rect -7152 4409 -7146 4443
rect -7192 4371 -7146 4409
rect -7192 4337 -7186 4371
rect -7152 4337 -7146 4371
rect -7192 4299 -7146 4337
rect -7192 4265 -7186 4299
rect -7152 4265 -7146 4299
rect -7192 4227 -7146 4265
rect -7192 4193 -7186 4227
rect -7152 4193 -7146 4227
rect -7192 4155 -7146 4193
rect -7192 4121 -7186 4155
rect -7152 4121 -7146 4155
rect -7192 4083 -7146 4121
rect -7192 4049 -7186 4083
rect -7152 4049 -7146 4083
rect -7192 4011 -7146 4049
rect -7192 3977 -7186 4011
rect -7152 3977 -7146 4011
rect -7192 3939 -7146 3977
rect -7192 3905 -7186 3939
rect -7152 3905 -7146 3939
rect -7192 3867 -7146 3905
rect -7192 3833 -7186 3867
rect -7152 3833 -7146 3867
rect -7192 3795 -7146 3833
rect -7192 3761 -7186 3795
rect -7152 3761 -7146 3795
rect -7192 3723 -7146 3761
rect -7192 3689 -7186 3723
rect -7152 3689 -7146 3723
rect -7192 3651 -7146 3689
rect -7192 3617 -7186 3651
rect -7152 3617 -7146 3651
rect -7192 3579 -7146 3617
rect -7192 3545 -7186 3579
rect -7152 3545 -7146 3579
rect -7192 3507 -7146 3545
rect -7192 3473 -7186 3507
rect -7152 3473 -7146 3507
rect -7192 3458 -7146 3473
rect -7096 4443 -7050 4458
rect -7096 4409 -7090 4443
rect -7056 4409 -7050 4443
rect -7096 4371 -7050 4409
rect -7096 4337 -7090 4371
rect -7056 4337 -7050 4371
rect -7096 4299 -7050 4337
rect -7096 4265 -7090 4299
rect -7056 4265 -7050 4299
rect -7096 4227 -7050 4265
rect -7096 4193 -7090 4227
rect -7056 4193 -7050 4227
rect -7096 4155 -7050 4193
rect -7096 4121 -7090 4155
rect -7056 4121 -7050 4155
rect -7096 4083 -7050 4121
rect -7096 4049 -7090 4083
rect -7056 4049 -7050 4083
rect -7096 4011 -7050 4049
rect -7096 3977 -7090 4011
rect -7056 3977 -7050 4011
rect -7096 3939 -7050 3977
rect -7096 3905 -7090 3939
rect -7056 3905 -7050 3939
rect -7096 3867 -7050 3905
rect -7096 3833 -7090 3867
rect -7056 3833 -7050 3867
rect -7096 3795 -7050 3833
rect -7096 3761 -7090 3795
rect -7056 3761 -7050 3795
rect -7096 3723 -7050 3761
rect -7096 3689 -7090 3723
rect -7056 3689 -7050 3723
rect -7096 3651 -7050 3689
rect -7096 3617 -7090 3651
rect -7056 3617 -7050 3651
rect -7096 3579 -7050 3617
rect -7096 3545 -7090 3579
rect -7056 3545 -7050 3579
rect -7096 3507 -7050 3545
rect -7096 3473 -7090 3507
rect -7056 3473 -7050 3507
rect -7096 3458 -7050 3473
rect -7000 4443 -6954 4458
rect -7000 4409 -6994 4443
rect -6960 4409 -6954 4443
rect -7000 4371 -6954 4409
rect -7000 4337 -6994 4371
rect -6960 4337 -6954 4371
rect -7000 4299 -6954 4337
rect -7000 4265 -6994 4299
rect -6960 4265 -6954 4299
rect -7000 4227 -6954 4265
rect -7000 4193 -6994 4227
rect -6960 4193 -6954 4227
rect -7000 4155 -6954 4193
rect -7000 4121 -6994 4155
rect -6960 4121 -6954 4155
rect -7000 4083 -6954 4121
rect -7000 4049 -6994 4083
rect -6960 4049 -6954 4083
rect -7000 4011 -6954 4049
rect -7000 3977 -6994 4011
rect -6960 3977 -6954 4011
rect -7000 3939 -6954 3977
rect -7000 3905 -6994 3939
rect -6960 3905 -6954 3939
rect -7000 3867 -6954 3905
rect -7000 3833 -6994 3867
rect -6960 3833 -6954 3867
rect -7000 3795 -6954 3833
rect -7000 3761 -6994 3795
rect -6960 3761 -6954 3795
rect -7000 3723 -6954 3761
rect -7000 3689 -6994 3723
rect -6960 3689 -6954 3723
rect -7000 3651 -6954 3689
rect -7000 3617 -6994 3651
rect -6960 3617 -6954 3651
rect -7000 3579 -6954 3617
rect -7000 3545 -6994 3579
rect -6960 3545 -6954 3579
rect -7000 3507 -6954 3545
rect -7000 3473 -6994 3507
rect -6960 3473 -6954 3507
rect -7000 3458 -6954 3473
rect -6904 4443 -6858 4458
rect -6904 4409 -6898 4443
rect -6864 4409 -6858 4443
rect -6904 4371 -6858 4409
rect -6904 4337 -6898 4371
rect -6864 4337 -6858 4371
rect -6904 4299 -6858 4337
rect -6904 4265 -6898 4299
rect -6864 4265 -6858 4299
rect -6904 4227 -6858 4265
rect -6904 4193 -6898 4227
rect -6864 4193 -6858 4227
rect -6904 4155 -6858 4193
rect -6904 4121 -6898 4155
rect -6864 4121 -6858 4155
rect -6904 4083 -6858 4121
rect -6904 4049 -6898 4083
rect -6864 4049 -6858 4083
rect -6904 4011 -6858 4049
rect -6904 3977 -6898 4011
rect -6864 3977 -6858 4011
rect -6904 3939 -6858 3977
rect -6904 3905 -6898 3939
rect -6864 3905 -6858 3939
rect -6904 3867 -6858 3905
rect -6904 3833 -6898 3867
rect -6864 3833 -6858 3867
rect -6904 3795 -6858 3833
rect -6904 3761 -6898 3795
rect -6864 3761 -6858 3795
rect -6904 3723 -6858 3761
rect -6904 3689 -6898 3723
rect -6864 3689 -6858 3723
rect -6904 3651 -6858 3689
rect -6904 3617 -6898 3651
rect -6864 3617 -6858 3651
rect -6904 3579 -6858 3617
rect -6904 3545 -6898 3579
rect -6864 3545 -6858 3579
rect -6904 3507 -6858 3545
rect -6904 3473 -6898 3507
rect -6864 3473 -6858 3507
rect -6904 3458 -6858 3473
rect -6808 4443 -6762 4458
rect -6808 4409 -6802 4443
rect -6768 4409 -6762 4443
rect -6808 4371 -6762 4409
rect -6808 4337 -6802 4371
rect -6768 4337 -6762 4371
rect -6808 4299 -6762 4337
rect -6808 4265 -6802 4299
rect -6768 4265 -6762 4299
rect -6808 4227 -6762 4265
rect -6808 4193 -6802 4227
rect -6768 4193 -6762 4227
rect -6808 4155 -6762 4193
rect -6808 4121 -6802 4155
rect -6768 4121 -6762 4155
rect -6808 4083 -6762 4121
rect -6808 4049 -6802 4083
rect -6768 4049 -6762 4083
rect -6808 4011 -6762 4049
rect -6808 3977 -6802 4011
rect -6768 3977 -6762 4011
rect -6808 3939 -6762 3977
rect -6808 3905 -6802 3939
rect -6768 3905 -6762 3939
rect -6808 3867 -6762 3905
rect -6808 3833 -6802 3867
rect -6768 3833 -6762 3867
rect -6808 3795 -6762 3833
rect -6808 3761 -6802 3795
rect -6768 3761 -6762 3795
rect -6808 3723 -6762 3761
rect -6808 3689 -6802 3723
rect -6768 3689 -6762 3723
rect -6808 3651 -6762 3689
rect -6808 3617 -6802 3651
rect -6768 3617 -6762 3651
rect -6808 3579 -6762 3617
rect -6808 3545 -6802 3579
rect -6768 3545 -6762 3579
rect -6808 3507 -6762 3545
rect -6808 3473 -6802 3507
rect -6768 3473 -6762 3507
rect -6808 3458 -6762 3473
rect -6712 4443 -6666 4458
rect -6712 4409 -6706 4443
rect -6672 4409 -6666 4443
rect -6712 4371 -6666 4409
rect -6712 4337 -6706 4371
rect -6672 4337 -6666 4371
rect -6712 4299 -6666 4337
rect -6712 4265 -6706 4299
rect -6672 4265 -6666 4299
rect -6712 4227 -6666 4265
rect -6712 4193 -6706 4227
rect -6672 4193 -6666 4227
rect -6712 4155 -6666 4193
rect -6712 4121 -6706 4155
rect -6672 4121 -6666 4155
rect -6712 4083 -6666 4121
rect -6712 4049 -6706 4083
rect -6672 4049 -6666 4083
rect -6712 4011 -6666 4049
rect -6712 3977 -6706 4011
rect -6672 3977 -6666 4011
rect -6712 3939 -6666 3977
rect -6712 3905 -6706 3939
rect -6672 3905 -6666 3939
rect -6712 3867 -6666 3905
rect -6712 3833 -6706 3867
rect -6672 3833 -6666 3867
rect -6712 3795 -6666 3833
rect -6712 3761 -6706 3795
rect -6672 3761 -6666 3795
rect -6712 3723 -6666 3761
rect -6712 3689 -6706 3723
rect -6672 3689 -6666 3723
rect -6712 3651 -6666 3689
rect -6712 3617 -6706 3651
rect -6672 3617 -6666 3651
rect -6712 3579 -6666 3617
rect -6712 3545 -6706 3579
rect -6672 3545 -6666 3579
rect -6712 3507 -6666 3545
rect -6712 3473 -6706 3507
rect -6672 3473 -6666 3507
rect -6712 3458 -6666 3473
rect -6468 4449 -6422 4464
rect -6468 4415 -6462 4449
rect -6428 4415 -6422 4449
rect -6468 4377 -6422 4415
rect -6468 4343 -6462 4377
rect -6428 4343 -6422 4377
rect -6468 4305 -6422 4343
rect -6468 4271 -6462 4305
rect -6428 4271 -6422 4305
rect -6468 4233 -6422 4271
rect -6468 4199 -6462 4233
rect -6428 4199 -6422 4233
rect -6468 4161 -6422 4199
rect -6468 4127 -6462 4161
rect -6428 4127 -6422 4161
rect -6468 4089 -6422 4127
rect -6468 4055 -6462 4089
rect -6428 4055 -6422 4089
rect -6468 4017 -6422 4055
rect -6468 3983 -6462 4017
rect -6428 3983 -6422 4017
rect -6468 3945 -6422 3983
rect -6468 3911 -6462 3945
rect -6428 3911 -6422 3945
rect -6468 3873 -6422 3911
rect -6468 3839 -6462 3873
rect -6428 3839 -6422 3873
rect -6468 3801 -6422 3839
rect -6468 3767 -6462 3801
rect -6428 3767 -6422 3801
rect -6468 3729 -6422 3767
rect -6468 3695 -6462 3729
rect -6428 3695 -6422 3729
rect -6468 3657 -6422 3695
rect -6468 3623 -6462 3657
rect -6428 3623 -6422 3657
rect -6468 3585 -6422 3623
rect -6468 3551 -6462 3585
rect -6428 3551 -6422 3585
rect -6468 3513 -6422 3551
rect -6468 3479 -6462 3513
rect -6428 3479 -6422 3513
rect -6468 3464 -6422 3479
rect -6372 4449 -6326 4464
rect -6372 4415 -6366 4449
rect -6332 4415 -6326 4449
rect -6372 4377 -6326 4415
rect -6372 4343 -6366 4377
rect -6332 4343 -6326 4377
rect -6372 4305 -6326 4343
rect -6372 4271 -6366 4305
rect -6332 4271 -6326 4305
rect -6372 4233 -6326 4271
rect -6372 4199 -6366 4233
rect -6332 4199 -6326 4233
rect -6372 4161 -6326 4199
rect -6372 4127 -6366 4161
rect -6332 4127 -6326 4161
rect -6372 4089 -6326 4127
rect -6372 4055 -6366 4089
rect -6332 4055 -6326 4089
rect -6372 4017 -6326 4055
rect -6372 3983 -6366 4017
rect -6332 3983 -6326 4017
rect -6372 3945 -6326 3983
rect -6372 3911 -6366 3945
rect -6332 3911 -6326 3945
rect -6372 3873 -6326 3911
rect -6372 3839 -6366 3873
rect -6332 3839 -6326 3873
rect -6372 3801 -6326 3839
rect -6372 3767 -6366 3801
rect -6332 3767 -6326 3801
rect -6372 3729 -6326 3767
rect -6372 3695 -6366 3729
rect -6332 3695 -6326 3729
rect -6372 3657 -6326 3695
rect -6372 3623 -6366 3657
rect -6332 3623 -6326 3657
rect -6372 3585 -6326 3623
rect -6372 3551 -6366 3585
rect -6332 3551 -6326 3585
rect -6372 3513 -6326 3551
rect -6372 3479 -6366 3513
rect -6332 3479 -6326 3513
rect -6372 3464 -6326 3479
rect -6276 4449 -6230 4464
rect -6276 4415 -6270 4449
rect -6236 4415 -6230 4449
rect -6276 4377 -6230 4415
rect -6276 4343 -6270 4377
rect -6236 4343 -6230 4377
rect -6276 4305 -6230 4343
rect -6276 4271 -6270 4305
rect -6236 4271 -6230 4305
rect -6276 4233 -6230 4271
rect -6276 4199 -6270 4233
rect -6236 4199 -6230 4233
rect -6276 4161 -6230 4199
rect -6276 4127 -6270 4161
rect -6236 4127 -6230 4161
rect -6276 4089 -6230 4127
rect -6276 4055 -6270 4089
rect -6236 4055 -6230 4089
rect -6276 4017 -6230 4055
rect -6276 3983 -6270 4017
rect -6236 3983 -6230 4017
rect -6276 3945 -6230 3983
rect -6276 3911 -6270 3945
rect -6236 3911 -6230 3945
rect -6276 3873 -6230 3911
rect -6276 3839 -6270 3873
rect -6236 3839 -6230 3873
rect -6276 3801 -6230 3839
rect -6276 3767 -6270 3801
rect -6236 3767 -6230 3801
rect -6276 3729 -6230 3767
rect -6276 3695 -6270 3729
rect -6236 3695 -6230 3729
rect -6276 3657 -6230 3695
rect -6276 3623 -6270 3657
rect -6236 3623 -6230 3657
rect -6276 3585 -6230 3623
rect -6276 3551 -6270 3585
rect -6236 3551 -6230 3585
rect -6276 3513 -6230 3551
rect -6276 3479 -6270 3513
rect -6236 3479 -6230 3513
rect -6276 3464 -6230 3479
rect -6180 4449 -6134 4464
rect -6180 4415 -6174 4449
rect -6140 4415 -6134 4449
rect -6180 4377 -6134 4415
rect -6180 4343 -6174 4377
rect -6140 4343 -6134 4377
rect -6180 4305 -6134 4343
rect -6180 4271 -6174 4305
rect -6140 4271 -6134 4305
rect -6180 4233 -6134 4271
rect -6180 4199 -6174 4233
rect -6140 4199 -6134 4233
rect -6180 4161 -6134 4199
rect -6180 4127 -6174 4161
rect -6140 4127 -6134 4161
rect -6180 4089 -6134 4127
rect -6180 4055 -6174 4089
rect -6140 4055 -6134 4089
rect -6180 4017 -6134 4055
rect -6180 3983 -6174 4017
rect -6140 3983 -6134 4017
rect -6180 3945 -6134 3983
rect -6180 3911 -6174 3945
rect -6140 3911 -6134 3945
rect -6180 3873 -6134 3911
rect -6180 3839 -6174 3873
rect -6140 3839 -6134 3873
rect -6180 3801 -6134 3839
rect -6180 3767 -6174 3801
rect -6140 3767 -6134 3801
rect -6180 3729 -6134 3767
rect -6180 3695 -6174 3729
rect -6140 3695 -6134 3729
rect -6180 3657 -6134 3695
rect -6180 3623 -6174 3657
rect -6140 3623 -6134 3657
rect -6180 3585 -6134 3623
rect -6180 3551 -6174 3585
rect -6140 3551 -6134 3585
rect -6180 3513 -6134 3551
rect -6180 3479 -6174 3513
rect -6140 3479 -6134 3513
rect -6180 3464 -6134 3479
rect -6084 4449 -6038 4464
rect -6084 4415 -6078 4449
rect -6044 4415 -6038 4449
rect -6084 4377 -6038 4415
rect -6084 4343 -6078 4377
rect -6044 4343 -6038 4377
rect -6084 4305 -6038 4343
rect -6084 4271 -6078 4305
rect -6044 4271 -6038 4305
rect -6084 4233 -6038 4271
rect -6084 4199 -6078 4233
rect -6044 4199 -6038 4233
rect -6084 4161 -6038 4199
rect -6084 4127 -6078 4161
rect -6044 4127 -6038 4161
rect -6084 4089 -6038 4127
rect -6084 4055 -6078 4089
rect -6044 4055 -6038 4089
rect -6084 4017 -6038 4055
rect -6084 3983 -6078 4017
rect -6044 3983 -6038 4017
rect -6084 3945 -6038 3983
rect -6084 3911 -6078 3945
rect -6044 3911 -6038 3945
rect -6084 3873 -6038 3911
rect -6084 3839 -6078 3873
rect -6044 3839 -6038 3873
rect -6084 3801 -6038 3839
rect -6084 3767 -6078 3801
rect -6044 3767 -6038 3801
rect -6084 3729 -6038 3767
rect -6084 3695 -6078 3729
rect -6044 3695 -6038 3729
rect -6084 3657 -6038 3695
rect -6084 3623 -6078 3657
rect -6044 3623 -6038 3657
rect -6084 3585 -6038 3623
rect -6084 3551 -6078 3585
rect -6044 3551 -6038 3585
rect -6084 3513 -6038 3551
rect -6084 3479 -6078 3513
rect -6044 3479 -6038 3513
rect -6084 3464 -6038 3479
rect -5988 4449 -5942 4464
rect -5988 4415 -5982 4449
rect -5948 4415 -5942 4449
rect -5988 4377 -5942 4415
rect -5988 4343 -5982 4377
rect -5948 4343 -5942 4377
rect -5988 4305 -5942 4343
rect -5988 4271 -5982 4305
rect -5948 4271 -5942 4305
rect -5988 4233 -5942 4271
rect -5988 4199 -5982 4233
rect -5948 4199 -5942 4233
rect -5988 4161 -5942 4199
rect -5988 4127 -5982 4161
rect -5948 4127 -5942 4161
rect -5988 4089 -5942 4127
rect -5988 4055 -5982 4089
rect -5948 4055 -5942 4089
rect -5988 4017 -5942 4055
rect -5988 3983 -5982 4017
rect -5948 3983 -5942 4017
rect -5988 3945 -5942 3983
rect -5988 3911 -5982 3945
rect -5948 3911 -5942 3945
rect -5988 3873 -5942 3911
rect -5988 3839 -5982 3873
rect -5948 3839 -5942 3873
rect -5988 3801 -5942 3839
rect -5988 3767 -5982 3801
rect -5948 3767 -5942 3801
rect -5988 3729 -5942 3767
rect -5988 3695 -5982 3729
rect -5948 3695 -5942 3729
rect -5988 3657 -5942 3695
rect -5988 3623 -5982 3657
rect -5948 3623 -5942 3657
rect -5988 3585 -5942 3623
rect -5988 3551 -5982 3585
rect -5948 3551 -5942 3585
rect -5988 3513 -5942 3551
rect -5988 3479 -5982 3513
rect -5948 3479 -5942 3513
rect -5988 3464 -5942 3479
rect -5892 4449 -5846 4464
rect -5892 4415 -5886 4449
rect -5852 4415 -5846 4449
rect -5892 4377 -5846 4415
rect -5892 4343 -5886 4377
rect -5852 4343 -5846 4377
rect -5892 4305 -5846 4343
rect -5892 4271 -5886 4305
rect -5852 4271 -5846 4305
rect -5892 4233 -5846 4271
rect -5892 4199 -5886 4233
rect -5852 4199 -5846 4233
rect -5892 4161 -5846 4199
rect -5892 4127 -5886 4161
rect -5852 4127 -5846 4161
rect -5892 4089 -5846 4127
rect -5892 4055 -5886 4089
rect -5852 4055 -5846 4089
rect -5892 4017 -5846 4055
rect -5892 3983 -5886 4017
rect -5852 3983 -5846 4017
rect -5892 3945 -5846 3983
rect -5892 3911 -5886 3945
rect -5852 3911 -5846 3945
rect -5892 3873 -5846 3911
rect -5892 3839 -5886 3873
rect -5852 3839 -5846 3873
rect -5892 3801 -5846 3839
rect -5892 3767 -5886 3801
rect -5852 3767 -5846 3801
rect -5892 3729 -5846 3767
rect -5892 3695 -5886 3729
rect -5852 3695 -5846 3729
rect -5892 3657 -5846 3695
rect -5892 3623 -5886 3657
rect -5852 3623 -5846 3657
rect -5892 3585 -5846 3623
rect -5892 3551 -5886 3585
rect -5852 3551 -5846 3585
rect -5892 3513 -5846 3551
rect -5892 3479 -5886 3513
rect -5852 3479 -5846 3513
rect -5892 3464 -5846 3479
rect -5796 4449 -5750 4464
rect -5796 4415 -5790 4449
rect -5756 4415 -5750 4449
rect -5796 4377 -5750 4415
rect -5796 4343 -5790 4377
rect -5756 4343 -5750 4377
rect -5796 4305 -5750 4343
rect -5796 4271 -5790 4305
rect -5756 4271 -5750 4305
rect -5796 4233 -5750 4271
rect -5796 4199 -5790 4233
rect -5756 4199 -5750 4233
rect -5796 4161 -5750 4199
rect -5796 4127 -5790 4161
rect -5756 4127 -5750 4161
rect -5796 4089 -5750 4127
rect -5796 4055 -5790 4089
rect -5756 4055 -5750 4089
rect -5796 4017 -5750 4055
rect -5796 3983 -5790 4017
rect -5756 3983 -5750 4017
rect -5796 3945 -5750 3983
rect -5796 3911 -5790 3945
rect -5756 3911 -5750 3945
rect -5796 3873 -5750 3911
rect -5796 3839 -5790 3873
rect -5756 3839 -5750 3873
rect -5796 3801 -5750 3839
rect -5796 3767 -5790 3801
rect -5756 3767 -5750 3801
rect -5796 3729 -5750 3767
rect -5796 3695 -5790 3729
rect -5756 3695 -5750 3729
rect -5796 3657 -5750 3695
rect -5796 3623 -5790 3657
rect -5756 3623 -5750 3657
rect -5796 3585 -5750 3623
rect -5796 3551 -5790 3585
rect -5756 3551 -5750 3585
rect -5796 3513 -5750 3551
rect -5796 3479 -5790 3513
rect -5756 3479 -5750 3513
rect -5796 3464 -5750 3479
rect -5700 4449 -5654 4464
rect -5700 4415 -5694 4449
rect -5660 4415 -5654 4449
rect -5700 4377 -5654 4415
rect -5700 4343 -5694 4377
rect -5660 4343 -5654 4377
rect -5700 4305 -5654 4343
rect -5700 4271 -5694 4305
rect -5660 4271 -5654 4305
rect -5700 4233 -5654 4271
rect -5700 4199 -5694 4233
rect -5660 4199 -5654 4233
rect -5700 4161 -5654 4199
rect -5700 4127 -5694 4161
rect -5660 4127 -5654 4161
rect -5700 4089 -5654 4127
rect -5700 4055 -5694 4089
rect -5660 4055 -5654 4089
rect -5700 4017 -5654 4055
rect -5700 3983 -5694 4017
rect -5660 3983 -5654 4017
rect -5700 3945 -5654 3983
rect -5700 3911 -5694 3945
rect -5660 3911 -5654 3945
rect -5700 3873 -5654 3911
rect -5700 3839 -5694 3873
rect -5660 3839 -5654 3873
rect -5700 3801 -5654 3839
rect -5700 3767 -5694 3801
rect -5660 3767 -5654 3801
rect -5700 3729 -5654 3767
rect -5700 3695 -5694 3729
rect -5660 3695 -5654 3729
rect -5700 3657 -5654 3695
rect -5700 3623 -5694 3657
rect -5660 3623 -5654 3657
rect -5700 3585 -5654 3623
rect -5700 3551 -5694 3585
rect -5660 3551 -5654 3585
rect -5700 3513 -5654 3551
rect -5700 3479 -5694 3513
rect -5660 3479 -5654 3513
rect -5700 3464 -5654 3479
rect -5604 4449 -5558 4464
rect -5604 4415 -5598 4449
rect -5564 4415 -5558 4449
rect -5604 4377 -5558 4415
rect -5604 4343 -5598 4377
rect -5564 4343 -5558 4377
rect -5604 4305 -5558 4343
rect -5604 4271 -5598 4305
rect -5564 4271 -5558 4305
rect -5604 4233 -5558 4271
rect -5604 4199 -5598 4233
rect -5564 4199 -5558 4233
rect -5604 4161 -5558 4199
rect -5604 4127 -5598 4161
rect -5564 4127 -5558 4161
rect -5604 4089 -5558 4127
rect -5604 4055 -5598 4089
rect -5564 4055 -5558 4089
rect -5604 4017 -5558 4055
rect -5604 3983 -5598 4017
rect -5564 3983 -5558 4017
rect -5604 3945 -5558 3983
rect -5604 3911 -5598 3945
rect -5564 3911 -5558 3945
rect -5604 3873 -5558 3911
rect -5604 3839 -5598 3873
rect -5564 3839 -5558 3873
rect -5604 3801 -5558 3839
rect -5604 3767 -5598 3801
rect -5564 3767 -5558 3801
rect -5604 3729 -5558 3767
rect -5604 3695 -5598 3729
rect -5564 3695 -5558 3729
rect -5604 3657 -5558 3695
rect -5604 3623 -5598 3657
rect -5564 3623 -5558 3657
rect -5604 3585 -5558 3623
rect -5604 3551 -5598 3585
rect -5564 3551 -5558 3585
rect -5604 3513 -5558 3551
rect -5604 3479 -5598 3513
rect -5564 3479 -5558 3513
rect -5604 3464 -5558 3479
rect -5508 4449 -5462 4464
rect -5508 4415 -5502 4449
rect -5468 4415 -5462 4449
rect -5508 4377 -5462 4415
rect -5508 4343 -5502 4377
rect -5468 4343 -5462 4377
rect -5508 4305 -5462 4343
rect -5508 4271 -5502 4305
rect -5468 4271 -5462 4305
rect -5508 4233 -5462 4271
rect -5508 4199 -5502 4233
rect -5468 4199 -5462 4233
rect -5508 4161 -5462 4199
rect -5508 4127 -5502 4161
rect -5468 4127 -5462 4161
rect -5508 4089 -5462 4127
rect -5508 4055 -5502 4089
rect -5468 4055 -5462 4089
rect -5508 4017 -5462 4055
rect -5508 3983 -5502 4017
rect -5468 3983 -5462 4017
rect -5508 3945 -5462 3983
rect -5508 3911 -5502 3945
rect -5468 3911 -5462 3945
rect -5508 3873 -5462 3911
rect -5508 3839 -5502 3873
rect -5468 3839 -5462 3873
rect -5508 3801 -5462 3839
rect -5508 3767 -5502 3801
rect -5468 3767 -5462 3801
rect -5508 3729 -5462 3767
rect -5508 3695 -5502 3729
rect -5468 3695 -5462 3729
rect -5508 3657 -5462 3695
rect -5508 3623 -5502 3657
rect -5468 3623 -5462 3657
rect -5508 3585 -5462 3623
rect -5508 3551 -5502 3585
rect -5468 3551 -5462 3585
rect -5508 3513 -5462 3551
rect -5508 3479 -5502 3513
rect -5468 3479 -5462 3513
rect -5508 3464 -5462 3479
rect -5300 4451 -5254 4466
rect -5300 4417 -5294 4451
rect -5260 4417 -5254 4451
rect -5300 4379 -5254 4417
rect -5300 4345 -5294 4379
rect -5260 4345 -5254 4379
rect -5300 4307 -5254 4345
rect -5300 4273 -5294 4307
rect -5260 4273 -5254 4307
rect -5300 4235 -5254 4273
rect -5300 4201 -5294 4235
rect -5260 4201 -5254 4235
rect -5300 4163 -5254 4201
rect -5300 4129 -5294 4163
rect -5260 4129 -5254 4163
rect -5300 4091 -5254 4129
rect -5300 4057 -5294 4091
rect -5260 4057 -5254 4091
rect -5300 4019 -5254 4057
rect -5300 3985 -5294 4019
rect -5260 3985 -5254 4019
rect -5300 3947 -5254 3985
rect -5300 3913 -5294 3947
rect -5260 3913 -5254 3947
rect -5300 3875 -5254 3913
rect -5300 3841 -5294 3875
rect -5260 3841 -5254 3875
rect -5300 3803 -5254 3841
rect -5300 3769 -5294 3803
rect -5260 3769 -5254 3803
rect -5300 3731 -5254 3769
rect -5300 3697 -5294 3731
rect -5260 3697 -5254 3731
rect -5300 3659 -5254 3697
rect -5300 3625 -5294 3659
rect -5260 3625 -5254 3659
rect -5300 3587 -5254 3625
rect -5300 3553 -5294 3587
rect -5260 3553 -5254 3587
rect -5300 3515 -5254 3553
rect -5300 3481 -5294 3515
rect -5260 3481 -5254 3515
rect -5300 3466 -5254 3481
rect -5204 4451 -5158 4466
rect -5204 4417 -5198 4451
rect -5164 4417 -5158 4451
rect -5204 4379 -5158 4417
rect -5204 4345 -5198 4379
rect -5164 4345 -5158 4379
rect -5204 4307 -5158 4345
rect -5204 4273 -5198 4307
rect -5164 4273 -5158 4307
rect -5204 4235 -5158 4273
rect -5204 4201 -5198 4235
rect -5164 4201 -5158 4235
rect -5204 4163 -5158 4201
rect -5204 4129 -5198 4163
rect -5164 4129 -5158 4163
rect -5204 4091 -5158 4129
rect -5204 4057 -5198 4091
rect -5164 4057 -5158 4091
rect -5204 4019 -5158 4057
rect -5204 3985 -5198 4019
rect -5164 3985 -5158 4019
rect -5204 3947 -5158 3985
rect -5204 3913 -5198 3947
rect -5164 3913 -5158 3947
rect -5204 3875 -5158 3913
rect -5204 3841 -5198 3875
rect -5164 3841 -5158 3875
rect -5204 3803 -5158 3841
rect -5204 3769 -5198 3803
rect -5164 3769 -5158 3803
rect -5204 3731 -5158 3769
rect -5204 3697 -5198 3731
rect -5164 3697 -5158 3731
rect -5204 3659 -5158 3697
rect -5204 3625 -5198 3659
rect -5164 3625 -5158 3659
rect -5204 3587 -5158 3625
rect -5204 3553 -5198 3587
rect -5164 3553 -5158 3587
rect -5204 3515 -5158 3553
rect -5204 3481 -5198 3515
rect -5164 3481 -5158 3515
rect -5204 3466 -5158 3481
rect -5108 4451 -5062 4466
rect -5108 4417 -5102 4451
rect -5068 4417 -5062 4451
rect -5108 4379 -5062 4417
rect -5108 4345 -5102 4379
rect -5068 4345 -5062 4379
rect -5108 4307 -5062 4345
rect -5108 4273 -5102 4307
rect -5068 4273 -5062 4307
rect -5108 4235 -5062 4273
rect -5108 4201 -5102 4235
rect -5068 4201 -5062 4235
rect -5108 4163 -5062 4201
rect -5108 4129 -5102 4163
rect -5068 4129 -5062 4163
rect -5108 4091 -5062 4129
rect -5108 4057 -5102 4091
rect -5068 4057 -5062 4091
rect -5108 4019 -5062 4057
rect -5108 3985 -5102 4019
rect -5068 3985 -5062 4019
rect -5108 3947 -5062 3985
rect -5108 3913 -5102 3947
rect -5068 3913 -5062 3947
rect -5108 3875 -5062 3913
rect -5108 3841 -5102 3875
rect -5068 3841 -5062 3875
rect -5108 3803 -5062 3841
rect -5108 3769 -5102 3803
rect -5068 3769 -5062 3803
rect -5108 3731 -5062 3769
rect -5108 3697 -5102 3731
rect -5068 3697 -5062 3731
rect -5108 3659 -5062 3697
rect -5108 3625 -5102 3659
rect -5068 3625 -5062 3659
rect -5108 3587 -5062 3625
rect -5108 3553 -5102 3587
rect -5068 3553 -5062 3587
rect -5108 3515 -5062 3553
rect -5108 3481 -5102 3515
rect -5068 3481 -5062 3515
rect -5108 3466 -5062 3481
rect -5012 4451 -4966 4466
rect -5012 4417 -5006 4451
rect -4972 4417 -4966 4451
rect -5012 4379 -4966 4417
rect -5012 4345 -5006 4379
rect -4972 4345 -4966 4379
rect -5012 4307 -4966 4345
rect -5012 4273 -5006 4307
rect -4972 4273 -4966 4307
rect -5012 4235 -4966 4273
rect -5012 4201 -5006 4235
rect -4972 4201 -4966 4235
rect -5012 4163 -4966 4201
rect -5012 4129 -5006 4163
rect -4972 4129 -4966 4163
rect -5012 4091 -4966 4129
rect -5012 4057 -5006 4091
rect -4972 4057 -4966 4091
rect -5012 4019 -4966 4057
rect -5012 3985 -5006 4019
rect -4972 3985 -4966 4019
rect -5012 3947 -4966 3985
rect -5012 3913 -5006 3947
rect -4972 3913 -4966 3947
rect -5012 3875 -4966 3913
rect -5012 3841 -5006 3875
rect -4972 3841 -4966 3875
rect -5012 3803 -4966 3841
rect -5012 3769 -5006 3803
rect -4972 3769 -4966 3803
rect -5012 3731 -4966 3769
rect -5012 3697 -5006 3731
rect -4972 3697 -4966 3731
rect -5012 3659 -4966 3697
rect -5012 3625 -5006 3659
rect -4972 3625 -4966 3659
rect -5012 3587 -4966 3625
rect -5012 3553 -5006 3587
rect -4972 3553 -4966 3587
rect -5012 3515 -4966 3553
rect -5012 3481 -5006 3515
rect -4972 3481 -4966 3515
rect -5012 3466 -4966 3481
rect -4916 4451 -4870 4466
rect -4916 4417 -4910 4451
rect -4876 4417 -4870 4451
rect -4916 4379 -4870 4417
rect -4916 4345 -4910 4379
rect -4876 4345 -4870 4379
rect -4916 4307 -4870 4345
rect -4916 4273 -4910 4307
rect -4876 4273 -4870 4307
rect -4916 4235 -4870 4273
rect -4916 4201 -4910 4235
rect -4876 4201 -4870 4235
rect -4916 4163 -4870 4201
rect -4916 4129 -4910 4163
rect -4876 4129 -4870 4163
rect -4916 4091 -4870 4129
rect -4916 4057 -4910 4091
rect -4876 4057 -4870 4091
rect -4916 4019 -4870 4057
rect -4916 3985 -4910 4019
rect -4876 3985 -4870 4019
rect -4916 3947 -4870 3985
rect -4916 3913 -4910 3947
rect -4876 3913 -4870 3947
rect -4916 3875 -4870 3913
rect -4916 3841 -4910 3875
rect -4876 3841 -4870 3875
rect -4916 3803 -4870 3841
rect -4916 3769 -4910 3803
rect -4876 3769 -4870 3803
rect -4916 3731 -4870 3769
rect -4916 3697 -4910 3731
rect -4876 3697 -4870 3731
rect -4916 3659 -4870 3697
rect -4916 3625 -4910 3659
rect -4876 3625 -4870 3659
rect -4916 3587 -4870 3625
rect -4916 3553 -4910 3587
rect -4876 3553 -4870 3587
rect -4916 3515 -4870 3553
rect -4916 3481 -4910 3515
rect -4876 3481 -4870 3515
rect -4916 3466 -4870 3481
rect -4820 4451 -4774 4466
rect -4820 4417 -4814 4451
rect -4780 4417 -4774 4451
rect -4820 4379 -4774 4417
rect -4820 4345 -4814 4379
rect -4780 4345 -4774 4379
rect -4820 4307 -4774 4345
rect -4820 4273 -4814 4307
rect -4780 4273 -4774 4307
rect -4820 4235 -4774 4273
rect -4820 4201 -4814 4235
rect -4780 4201 -4774 4235
rect -4820 4163 -4774 4201
rect -4820 4129 -4814 4163
rect -4780 4129 -4774 4163
rect -4820 4091 -4774 4129
rect -4820 4057 -4814 4091
rect -4780 4057 -4774 4091
rect -4820 4019 -4774 4057
rect -4820 3985 -4814 4019
rect -4780 3985 -4774 4019
rect -4820 3947 -4774 3985
rect -4820 3913 -4814 3947
rect -4780 3913 -4774 3947
rect -4820 3875 -4774 3913
rect -4820 3841 -4814 3875
rect -4780 3841 -4774 3875
rect -4820 3803 -4774 3841
rect -4820 3769 -4814 3803
rect -4780 3769 -4774 3803
rect -4820 3731 -4774 3769
rect -4820 3697 -4814 3731
rect -4780 3697 -4774 3731
rect -4820 3659 -4774 3697
rect -4820 3625 -4814 3659
rect -4780 3625 -4774 3659
rect -4820 3587 -4774 3625
rect -4820 3553 -4814 3587
rect -4780 3553 -4774 3587
rect -4820 3515 -4774 3553
rect -4820 3481 -4814 3515
rect -4780 3481 -4774 3515
rect -4820 3466 -4774 3481
rect -1932 3434 -1546 3442
rect -1932 3428 -1544 3434
rect -1932 3394 -1590 3428
rect -1556 3394 -1544 3428
rect -1932 3388 -1544 3394
rect -1932 3380 -1546 3388
rect -1932 3372 -1590 3380
rect -21754 3275 -21642 3320
rect -21754 3241 -21714 3275
rect -21680 3241 -21642 3275
rect -21754 3158 -21642 3241
rect -20082 3281 -19982 3312
rect -20082 3247 -20050 3281
rect -20016 3247 -19982 3281
rect -20082 3176 -19982 3247
rect -18872 3287 -18792 3318
rect -18872 3253 -18846 3287
rect -18812 3253 -18792 3287
rect -24838 3130 -22884 3150
rect -24838 3096 -22974 3130
rect -22940 3096 -22884 3130
rect -24838 3078 -22884 3096
rect -21754 3132 -20684 3158
rect -21754 3098 -20771 3132
rect -20737 3098 -20684 3132
rect -24838 -5898 -24532 3078
rect -21754 3074 -20684 3098
rect -20082 3145 -19030 3176
rect -20082 3111 -19118 3145
rect -19084 3111 -19030 3145
rect -20082 3080 -19030 3111
rect -18872 3166 -18792 3253
rect -18188 3269 -18090 3296
rect -18188 3235 -18158 3269
rect -18124 3235 -18090 3269
rect -18188 3172 -18090 3235
rect -14924 3287 -14812 3332
rect -14924 3253 -14884 3287
rect -14850 3253 -14812 3287
rect -18872 3147 -18240 3166
rect -18872 3113 -18302 3147
rect -18268 3113 -18240 3147
rect -18872 3096 -18240 3113
rect -18188 3150 -17754 3172
rect -14924 3170 -14812 3253
rect -13252 3293 -13152 3324
rect -13252 3259 -13220 3293
rect -13186 3259 -13152 3293
rect -13252 3188 -13152 3259
rect -12042 3299 -11962 3330
rect -12042 3265 -12016 3299
rect -11982 3265 -11962 3299
rect -18188 3140 -17744 3150
rect -21754 3016 -21642 3074
rect -21754 2982 -21716 3016
rect -21682 2982 -21642 3016
rect -21754 2942 -21642 2982
rect -20082 3018 -19982 3080
rect -20082 2984 -20048 3018
rect -20014 2984 -19982 3018
rect -18872 3062 -18792 3096
rect -18872 3028 -18850 3062
rect -18816 3028 -18792 3062
rect -18872 3006 -18792 3028
rect -18188 3088 -17870 3140
rect -17818 3088 -17806 3140
rect -17754 3088 -17744 3140
rect -18188 3078 -17744 3088
rect -17380 3142 -16054 3162
rect -17380 3108 -16144 3142
rect -16110 3108 -16054 3142
rect -17380 3090 -16054 3108
rect -14924 3144 -13854 3170
rect -14924 3110 -13941 3144
rect -13907 3110 -13854 3144
rect -18188 3068 -17754 3078
rect -18188 3032 -18090 3068
rect -20082 2958 -19982 2984
rect -18188 2998 -18158 3032
rect -18124 2998 -18090 3032
rect -18188 2972 -18090 2998
rect -23498 2839 -23452 2854
rect -23498 2805 -23492 2839
rect -23458 2805 -23452 2839
rect -23498 2767 -23452 2805
rect -23498 2733 -23492 2767
rect -23458 2733 -23452 2767
rect -23498 2695 -23452 2733
rect -23498 2661 -23492 2695
rect -23458 2661 -23452 2695
rect -23498 2623 -23452 2661
rect -23498 2589 -23492 2623
rect -23458 2589 -23452 2623
rect -23498 2551 -23452 2589
rect -23498 2517 -23492 2551
rect -23458 2517 -23452 2551
rect -23498 2479 -23452 2517
rect -23498 2445 -23492 2479
rect -23458 2445 -23452 2479
rect -23498 2407 -23452 2445
rect -23498 2373 -23492 2407
rect -23458 2373 -23452 2407
rect -23498 2335 -23452 2373
rect -23498 2301 -23492 2335
rect -23458 2301 -23452 2335
rect -23498 2263 -23452 2301
rect -23498 2229 -23492 2263
rect -23458 2229 -23452 2263
rect -23498 2191 -23452 2229
rect -23498 2157 -23492 2191
rect -23458 2157 -23452 2191
rect -23498 2119 -23452 2157
rect -23498 2085 -23492 2119
rect -23458 2085 -23452 2119
rect -23498 2047 -23452 2085
rect -23498 2013 -23492 2047
rect -23458 2013 -23452 2047
rect -23498 1975 -23452 2013
rect -23498 1941 -23492 1975
rect -23458 1941 -23452 1975
rect -23498 1903 -23452 1941
rect -23498 1869 -23492 1903
rect -23458 1869 -23452 1903
rect -23498 1854 -23452 1869
rect -23402 2839 -23356 2854
rect -23402 2805 -23396 2839
rect -23362 2805 -23356 2839
rect -23402 2767 -23356 2805
rect -23402 2733 -23396 2767
rect -23362 2733 -23356 2767
rect -23402 2695 -23356 2733
rect -23402 2661 -23396 2695
rect -23362 2661 -23356 2695
rect -23402 2623 -23356 2661
rect -23402 2589 -23396 2623
rect -23362 2589 -23356 2623
rect -23402 2551 -23356 2589
rect -23402 2517 -23396 2551
rect -23362 2517 -23356 2551
rect -23402 2479 -23356 2517
rect -23402 2445 -23396 2479
rect -23362 2445 -23356 2479
rect -23402 2407 -23356 2445
rect -23402 2373 -23396 2407
rect -23362 2373 -23356 2407
rect -23402 2335 -23356 2373
rect -23402 2301 -23396 2335
rect -23362 2301 -23356 2335
rect -23402 2263 -23356 2301
rect -23402 2229 -23396 2263
rect -23362 2229 -23356 2263
rect -23402 2191 -23356 2229
rect -23402 2157 -23396 2191
rect -23362 2157 -23356 2191
rect -23402 2119 -23356 2157
rect -23402 2085 -23396 2119
rect -23362 2085 -23356 2119
rect -23402 2047 -23356 2085
rect -23402 2013 -23396 2047
rect -23362 2013 -23356 2047
rect -23402 1975 -23356 2013
rect -23402 1941 -23396 1975
rect -23362 1941 -23356 1975
rect -23402 1903 -23356 1941
rect -23402 1869 -23396 1903
rect -23362 1869 -23356 1903
rect -23402 1854 -23356 1869
rect -23306 2839 -23260 2854
rect -23306 2805 -23300 2839
rect -23266 2805 -23260 2839
rect -23306 2767 -23260 2805
rect -23306 2733 -23300 2767
rect -23266 2733 -23260 2767
rect -23306 2695 -23260 2733
rect -23306 2661 -23300 2695
rect -23266 2661 -23260 2695
rect -23306 2623 -23260 2661
rect -23306 2589 -23300 2623
rect -23266 2589 -23260 2623
rect -23306 2551 -23260 2589
rect -23306 2517 -23300 2551
rect -23266 2517 -23260 2551
rect -23306 2479 -23260 2517
rect -23306 2445 -23300 2479
rect -23266 2445 -23260 2479
rect -23306 2407 -23260 2445
rect -23306 2373 -23300 2407
rect -23266 2373 -23260 2407
rect -23306 2335 -23260 2373
rect -23306 2301 -23300 2335
rect -23266 2301 -23260 2335
rect -23306 2263 -23260 2301
rect -23306 2229 -23300 2263
rect -23266 2229 -23260 2263
rect -23306 2191 -23260 2229
rect -23306 2157 -23300 2191
rect -23266 2157 -23260 2191
rect -23306 2119 -23260 2157
rect -23306 2085 -23300 2119
rect -23266 2085 -23260 2119
rect -23306 2047 -23260 2085
rect -23306 2013 -23300 2047
rect -23266 2013 -23260 2047
rect -23306 1975 -23260 2013
rect -23306 1941 -23300 1975
rect -23266 1941 -23260 1975
rect -23306 1903 -23260 1941
rect -23306 1869 -23300 1903
rect -23266 1869 -23260 1903
rect -23306 1854 -23260 1869
rect -23210 2839 -23164 2854
rect -23210 2805 -23204 2839
rect -23170 2805 -23164 2839
rect -23210 2767 -23164 2805
rect -23210 2733 -23204 2767
rect -23170 2733 -23164 2767
rect -23210 2695 -23164 2733
rect -23210 2661 -23204 2695
rect -23170 2661 -23164 2695
rect -23210 2623 -23164 2661
rect -23210 2589 -23204 2623
rect -23170 2589 -23164 2623
rect -23210 2551 -23164 2589
rect -23210 2517 -23204 2551
rect -23170 2517 -23164 2551
rect -23210 2479 -23164 2517
rect -23210 2445 -23204 2479
rect -23170 2445 -23164 2479
rect -23210 2407 -23164 2445
rect -23210 2373 -23204 2407
rect -23170 2373 -23164 2407
rect -23210 2335 -23164 2373
rect -23210 2301 -23204 2335
rect -23170 2301 -23164 2335
rect -23210 2263 -23164 2301
rect -23210 2229 -23204 2263
rect -23170 2229 -23164 2263
rect -23210 2191 -23164 2229
rect -23210 2157 -23204 2191
rect -23170 2157 -23164 2191
rect -23210 2119 -23164 2157
rect -23210 2085 -23204 2119
rect -23170 2085 -23164 2119
rect -23210 2047 -23164 2085
rect -23210 2013 -23204 2047
rect -23170 2013 -23164 2047
rect -23210 1975 -23164 2013
rect -23210 1941 -23204 1975
rect -23170 1941 -23164 1975
rect -23210 1903 -23164 1941
rect -23210 1869 -23204 1903
rect -23170 1869 -23164 1903
rect -23210 1854 -23164 1869
rect -23114 2839 -23068 2854
rect -23114 2805 -23108 2839
rect -23074 2805 -23068 2839
rect -23114 2767 -23068 2805
rect -23114 2733 -23108 2767
rect -23074 2733 -23068 2767
rect -23114 2695 -23068 2733
rect -23114 2661 -23108 2695
rect -23074 2661 -23068 2695
rect -23114 2623 -23068 2661
rect -23114 2589 -23108 2623
rect -23074 2589 -23068 2623
rect -23114 2551 -23068 2589
rect -23114 2517 -23108 2551
rect -23074 2517 -23068 2551
rect -23114 2479 -23068 2517
rect -23114 2445 -23108 2479
rect -23074 2445 -23068 2479
rect -23114 2407 -23068 2445
rect -23114 2373 -23108 2407
rect -23074 2373 -23068 2407
rect -23114 2335 -23068 2373
rect -23114 2301 -23108 2335
rect -23074 2301 -23068 2335
rect -23114 2263 -23068 2301
rect -23114 2229 -23108 2263
rect -23074 2229 -23068 2263
rect -23114 2191 -23068 2229
rect -23114 2157 -23108 2191
rect -23074 2157 -23068 2191
rect -23114 2119 -23068 2157
rect -23114 2085 -23108 2119
rect -23074 2085 -23068 2119
rect -23114 2047 -23068 2085
rect -23114 2013 -23108 2047
rect -23074 2013 -23068 2047
rect -23114 1975 -23068 2013
rect -23114 1941 -23108 1975
rect -23074 1941 -23068 1975
rect -23114 1903 -23068 1941
rect -23114 1869 -23108 1903
rect -23074 1869 -23068 1903
rect -23114 1854 -23068 1869
rect -23018 2839 -22972 2854
rect -23018 2805 -23012 2839
rect -22978 2805 -22972 2839
rect -23018 2767 -22972 2805
rect -23018 2733 -23012 2767
rect -22978 2733 -22972 2767
rect -23018 2695 -22972 2733
rect -23018 2661 -23012 2695
rect -22978 2661 -22972 2695
rect -23018 2623 -22972 2661
rect -23018 2589 -23012 2623
rect -22978 2589 -22972 2623
rect -23018 2551 -22972 2589
rect -23018 2517 -23012 2551
rect -22978 2517 -22972 2551
rect -23018 2479 -22972 2517
rect -23018 2445 -23012 2479
rect -22978 2445 -22972 2479
rect -23018 2407 -22972 2445
rect -23018 2373 -23012 2407
rect -22978 2373 -22972 2407
rect -23018 2335 -22972 2373
rect -23018 2301 -23012 2335
rect -22978 2301 -22972 2335
rect -23018 2263 -22972 2301
rect -23018 2229 -23012 2263
rect -22978 2229 -22972 2263
rect -23018 2191 -22972 2229
rect -23018 2157 -23012 2191
rect -22978 2157 -22972 2191
rect -23018 2119 -22972 2157
rect -23018 2085 -23012 2119
rect -22978 2085 -22972 2119
rect -23018 2047 -22972 2085
rect -23018 2013 -23012 2047
rect -22978 2013 -22972 2047
rect -23018 1975 -22972 2013
rect -23018 1941 -23012 1975
rect -22978 1941 -22972 1975
rect -23018 1903 -22972 1941
rect -23018 1869 -23012 1903
rect -22978 1869 -22972 1903
rect -23018 1854 -22972 1869
rect -22922 2839 -22876 2854
rect -22922 2805 -22916 2839
rect -22882 2805 -22876 2839
rect -22922 2767 -22876 2805
rect -22922 2733 -22916 2767
rect -22882 2733 -22876 2767
rect -22922 2695 -22876 2733
rect -22922 2661 -22916 2695
rect -22882 2661 -22876 2695
rect -22922 2623 -22876 2661
rect -22922 2589 -22916 2623
rect -22882 2589 -22876 2623
rect -22922 2551 -22876 2589
rect -22922 2517 -22916 2551
rect -22882 2517 -22876 2551
rect -22922 2479 -22876 2517
rect -22922 2445 -22916 2479
rect -22882 2445 -22876 2479
rect -22922 2407 -22876 2445
rect -22922 2373 -22916 2407
rect -22882 2373 -22876 2407
rect -22922 2335 -22876 2373
rect -22922 2301 -22916 2335
rect -22882 2301 -22876 2335
rect -22922 2263 -22876 2301
rect -22922 2229 -22916 2263
rect -22882 2229 -22876 2263
rect -22922 2191 -22876 2229
rect -22922 2157 -22916 2191
rect -22882 2157 -22876 2191
rect -22922 2119 -22876 2157
rect -22922 2085 -22916 2119
rect -22882 2085 -22876 2119
rect -22922 2047 -22876 2085
rect -22922 2013 -22916 2047
rect -22882 2013 -22876 2047
rect -22922 1975 -22876 2013
rect -22922 1941 -22916 1975
rect -22882 1941 -22876 1975
rect -22922 1903 -22876 1941
rect -22922 1869 -22916 1903
rect -22882 1869 -22876 1903
rect -22922 1854 -22876 1869
rect -22826 2839 -22780 2854
rect -22826 2805 -22820 2839
rect -22786 2805 -22780 2839
rect -22826 2767 -22780 2805
rect -22826 2733 -22820 2767
rect -22786 2733 -22780 2767
rect -22826 2695 -22780 2733
rect -22826 2661 -22820 2695
rect -22786 2661 -22780 2695
rect -22826 2623 -22780 2661
rect -22826 2589 -22820 2623
rect -22786 2589 -22780 2623
rect -22826 2551 -22780 2589
rect -22826 2517 -22820 2551
rect -22786 2517 -22780 2551
rect -22826 2479 -22780 2517
rect -22826 2445 -22820 2479
rect -22786 2445 -22780 2479
rect -22826 2407 -22780 2445
rect -22826 2373 -22820 2407
rect -22786 2373 -22780 2407
rect -22826 2335 -22780 2373
rect -22826 2301 -22820 2335
rect -22786 2301 -22780 2335
rect -22826 2263 -22780 2301
rect -22826 2229 -22820 2263
rect -22786 2229 -22780 2263
rect -22826 2191 -22780 2229
rect -22826 2157 -22820 2191
rect -22786 2157 -22780 2191
rect -22826 2119 -22780 2157
rect -22826 2085 -22820 2119
rect -22786 2085 -22780 2119
rect -22826 2047 -22780 2085
rect -22826 2013 -22820 2047
rect -22786 2013 -22780 2047
rect -22826 1975 -22780 2013
rect -22826 1941 -22820 1975
rect -22786 1941 -22780 1975
rect -22826 1903 -22780 1941
rect -22826 1869 -22820 1903
rect -22786 1869 -22780 1903
rect -22826 1854 -22780 1869
rect -22730 2839 -22684 2854
rect -22730 2805 -22724 2839
rect -22690 2805 -22684 2839
rect -22730 2767 -22684 2805
rect -22730 2733 -22724 2767
rect -22690 2733 -22684 2767
rect -22730 2695 -22684 2733
rect -22730 2661 -22724 2695
rect -22690 2661 -22684 2695
rect -22730 2623 -22684 2661
rect -22730 2589 -22724 2623
rect -22690 2589 -22684 2623
rect -22730 2551 -22684 2589
rect -22730 2517 -22724 2551
rect -22690 2517 -22684 2551
rect -22730 2479 -22684 2517
rect -22730 2445 -22724 2479
rect -22690 2445 -22684 2479
rect -22730 2407 -22684 2445
rect -22730 2373 -22724 2407
rect -22690 2373 -22684 2407
rect -22730 2335 -22684 2373
rect -22730 2301 -22724 2335
rect -22690 2301 -22684 2335
rect -22730 2263 -22684 2301
rect -22730 2229 -22724 2263
rect -22690 2229 -22684 2263
rect -22730 2191 -22684 2229
rect -22730 2157 -22724 2191
rect -22690 2157 -22684 2191
rect -22730 2119 -22684 2157
rect -22730 2085 -22724 2119
rect -22690 2085 -22684 2119
rect -22730 2047 -22684 2085
rect -22730 2013 -22724 2047
rect -22690 2013 -22684 2047
rect -22730 1975 -22684 2013
rect -22730 1941 -22724 1975
rect -22690 1941 -22684 1975
rect -22730 1903 -22684 1941
rect -22730 1869 -22724 1903
rect -22690 1869 -22684 1903
rect -22730 1854 -22684 1869
rect -22634 2839 -22588 2854
rect -22634 2805 -22628 2839
rect -22594 2805 -22588 2839
rect -22634 2767 -22588 2805
rect -22634 2733 -22628 2767
rect -22594 2733 -22588 2767
rect -22634 2695 -22588 2733
rect -22634 2661 -22628 2695
rect -22594 2661 -22588 2695
rect -22634 2623 -22588 2661
rect -22634 2589 -22628 2623
rect -22594 2589 -22588 2623
rect -22634 2551 -22588 2589
rect -22634 2517 -22628 2551
rect -22594 2517 -22588 2551
rect -22634 2479 -22588 2517
rect -22634 2445 -22628 2479
rect -22594 2445 -22588 2479
rect -22634 2407 -22588 2445
rect -22634 2373 -22628 2407
rect -22594 2373 -22588 2407
rect -22634 2335 -22588 2373
rect -22634 2301 -22628 2335
rect -22594 2301 -22588 2335
rect -22634 2263 -22588 2301
rect -22634 2229 -22628 2263
rect -22594 2229 -22588 2263
rect -22634 2191 -22588 2229
rect -22634 2157 -22628 2191
rect -22594 2157 -22588 2191
rect -22634 2119 -22588 2157
rect -22634 2085 -22628 2119
rect -22594 2085 -22588 2119
rect -22634 2047 -22588 2085
rect -22634 2013 -22628 2047
rect -22594 2013 -22588 2047
rect -22634 1975 -22588 2013
rect -22634 1941 -22628 1975
rect -22594 1941 -22588 1975
rect -22634 1903 -22588 1941
rect -22634 1869 -22628 1903
rect -22594 1869 -22588 1903
rect -22634 1854 -22588 1869
rect -22538 2839 -22492 2854
rect -22538 2805 -22532 2839
rect -22498 2805 -22492 2839
rect -22538 2767 -22492 2805
rect -22538 2733 -22532 2767
rect -22498 2733 -22492 2767
rect -22538 2695 -22492 2733
rect -22538 2661 -22532 2695
rect -22498 2661 -22492 2695
rect -22538 2623 -22492 2661
rect -22538 2589 -22532 2623
rect -22498 2589 -22492 2623
rect -22538 2551 -22492 2589
rect -22538 2517 -22532 2551
rect -22498 2517 -22492 2551
rect -22538 2479 -22492 2517
rect -22538 2445 -22532 2479
rect -22498 2445 -22492 2479
rect -22538 2407 -22492 2445
rect -22538 2373 -22532 2407
rect -22498 2373 -22492 2407
rect -22538 2335 -22492 2373
rect -22538 2301 -22532 2335
rect -22498 2301 -22492 2335
rect -22538 2263 -22492 2301
rect -22538 2229 -22532 2263
rect -22498 2229 -22492 2263
rect -22538 2191 -22492 2229
rect -22538 2157 -22532 2191
rect -22498 2157 -22492 2191
rect -22538 2119 -22492 2157
rect -22538 2085 -22532 2119
rect -22498 2085 -22492 2119
rect -22538 2047 -22492 2085
rect -22538 2013 -22532 2047
rect -22498 2013 -22492 2047
rect -22538 1975 -22492 2013
rect -22538 1941 -22532 1975
rect -22498 1941 -22492 1975
rect -22538 1903 -22492 1941
rect -22538 1869 -22532 1903
rect -22498 1869 -22492 1903
rect -22538 1854 -22492 1869
rect -22442 2839 -22396 2854
rect -22442 2805 -22436 2839
rect -22402 2805 -22396 2839
rect -22442 2767 -22396 2805
rect -22442 2733 -22436 2767
rect -22402 2733 -22396 2767
rect -22442 2695 -22396 2733
rect -22442 2661 -22436 2695
rect -22402 2661 -22396 2695
rect -22442 2623 -22396 2661
rect -22442 2589 -22436 2623
rect -22402 2589 -22396 2623
rect -22442 2551 -22396 2589
rect -22442 2517 -22436 2551
rect -22402 2517 -22396 2551
rect -22442 2479 -22396 2517
rect -22442 2445 -22436 2479
rect -22402 2445 -22396 2479
rect -22442 2407 -22396 2445
rect -22442 2373 -22436 2407
rect -22402 2373 -22396 2407
rect -22442 2335 -22396 2373
rect -22442 2301 -22436 2335
rect -22402 2301 -22396 2335
rect -22442 2263 -22396 2301
rect -22442 2229 -22436 2263
rect -22402 2229 -22396 2263
rect -22442 2191 -22396 2229
rect -22442 2157 -22436 2191
rect -22402 2157 -22396 2191
rect -22442 2119 -22396 2157
rect -22442 2085 -22436 2119
rect -22402 2085 -22396 2119
rect -22442 2047 -22396 2085
rect -22442 2013 -22436 2047
rect -22402 2013 -22396 2047
rect -22442 1975 -22396 2013
rect -22442 1941 -22436 1975
rect -22402 1941 -22396 1975
rect -22442 1903 -22396 1941
rect -22442 1869 -22436 1903
rect -22402 1869 -22396 1903
rect -22442 1854 -22396 1869
rect -22346 2839 -22300 2854
rect -22346 2805 -22340 2839
rect -22306 2805 -22300 2839
rect -22346 2767 -22300 2805
rect -22346 2733 -22340 2767
rect -22306 2733 -22300 2767
rect -22346 2695 -22300 2733
rect -22346 2661 -22340 2695
rect -22306 2661 -22300 2695
rect -22346 2623 -22300 2661
rect -22346 2589 -22340 2623
rect -22306 2589 -22300 2623
rect -22346 2551 -22300 2589
rect -22346 2517 -22340 2551
rect -22306 2517 -22300 2551
rect -22346 2479 -22300 2517
rect -22346 2445 -22340 2479
rect -22306 2445 -22300 2479
rect -22346 2407 -22300 2445
rect -22346 2373 -22340 2407
rect -22306 2373 -22300 2407
rect -22346 2335 -22300 2373
rect -22346 2301 -22340 2335
rect -22306 2301 -22300 2335
rect -22346 2263 -22300 2301
rect -22346 2229 -22340 2263
rect -22306 2229 -22300 2263
rect -22346 2191 -22300 2229
rect -22346 2157 -22340 2191
rect -22306 2157 -22300 2191
rect -22346 2119 -22300 2157
rect -22346 2085 -22340 2119
rect -22306 2085 -22300 2119
rect -22346 2047 -22300 2085
rect -22346 2013 -22340 2047
rect -22306 2013 -22300 2047
rect -22346 1975 -22300 2013
rect -22346 1941 -22340 1975
rect -22306 1941 -22300 1975
rect -22346 1903 -22300 1941
rect -22346 1869 -22340 1903
rect -22306 1869 -22300 1903
rect -22346 1854 -22300 1869
rect -22250 2839 -22204 2854
rect -22250 2805 -22244 2839
rect -22210 2805 -22204 2839
rect -22250 2767 -22204 2805
rect -22250 2733 -22244 2767
rect -22210 2733 -22204 2767
rect -22250 2695 -22204 2733
rect -22250 2661 -22244 2695
rect -22210 2661 -22204 2695
rect -22250 2623 -22204 2661
rect -22250 2589 -22244 2623
rect -22210 2589 -22204 2623
rect -22250 2551 -22204 2589
rect -22250 2517 -22244 2551
rect -22210 2517 -22204 2551
rect -22250 2479 -22204 2517
rect -22250 2445 -22244 2479
rect -22210 2445 -22204 2479
rect -22250 2407 -22204 2445
rect -22250 2373 -22244 2407
rect -22210 2373 -22204 2407
rect -22250 2335 -22204 2373
rect -22250 2301 -22244 2335
rect -22210 2301 -22204 2335
rect -22250 2263 -22204 2301
rect -22250 2229 -22244 2263
rect -22210 2229 -22204 2263
rect -22250 2191 -22204 2229
rect -22250 2157 -22244 2191
rect -22210 2157 -22204 2191
rect -22250 2119 -22204 2157
rect -22250 2085 -22244 2119
rect -22210 2085 -22204 2119
rect -22250 2047 -22204 2085
rect -22250 2013 -22244 2047
rect -22210 2013 -22204 2047
rect -22250 1975 -22204 2013
rect -22250 1941 -22244 1975
rect -22210 1941 -22204 1975
rect -22250 1903 -22204 1941
rect -22250 1869 -22244 1903
rect -22210 1869 -22204 1903
rect -22250 1854 -22204 1869
rect -22154 2839 -22108 2854
rect -22154 2805 -22148 2839
rect -22114 2805 -22108 2839
rect -22154 2767 -22108 2805
rect -22154 2733 -22148 2767
rect -22114 2733 -22108 2767
rect -22154 2695 -22108 2733
rect -22154 2661 -22148 2695
rect -22114 2661 -22108 2695
rect -22154 2623 -22108 2661
rect -22154 2589 -22148 2623
rect -22114 2589 -22108 2623
rect -22154 2551 -22108 2589
rect -22154 2517 -22148 2551
rect -22114 2517 -22108 2551
rect -22154 2479 -22108 2517
rect -22154 2445 -22148 2479
rect -22114 2445 -22108 2479
rect -22154 2407 -22108 2445
rect -22154 2373 -22148 2407
rect -22114 2373 -22108 2407
rect -22154 2335 -22108 2373
rect -22154 2301 -22148 2335
rect -22114 2301 -22108 2335
rect -22154 2263 -22108 2301
rect -22154 2229 -22148 2263
rect -22114 2229 -22108 2263
rect -22154 2191 -22108 2229
rect -22154 2157 -22148 2191
rect -22114 2157 -22108 2191
rect -22154 2119 -22108 2157
rect -22154 2085 -22148 2119
rect -22114 2085 -22108 2119
rect -22154 2047 -22108 2085
rect -22154 2013 -22148 2047
rect -22114 2013 -22108 2047
rect -22154 1975 -22108 2013
rect -22154 1941 -22148 1975
rect -22114 1941 -22108 1975
rect -22154 1903 -22108 1941
rect -22154 1869 -22148 1903
rect -22114 1869 -22108 1903
rect -22154 1854 -22108 1869
rect -22058 2839 -22012 2854
rect -22058 2805 -22052 2839
rect -22018 2805 -22012 2839
rect -22058 2767 -22012 2805
rect -22058 2733 -22052 2767
rect -22018 2733 -22012 2767
rect -22058 2695 -22012 2733
rect -22058 2661 -22052 2695
rect -22018 2661 -22012 2695
rect -22058 2623 -22012 2661
rect -22058 2589 -22052 2623
rect -22018 2589 -22012 2623
rect -22058 2551 -22012 2589
rect -22058 2517 -22052 2551
rect -22018 2517 -22012 2551
rect -22058 2479 -22012 2517
rect -22058 2445 -22052 2479
rect -22018 2445 -22012 2479
rect -22058 2407 -22012 2445
rect -22058 2373 -22052 2407
rect -22018 2373 -22012 2407
rect -22058 2335 -22012 2373
rect -22058 2301 -22052 2335
rect -22018 2301 -22012 2335
rect -22058 2263 -22012 2301
rect -22058 2229 -22052 2263
rect -22018 2229 -22012 2263
rect -22058 2191 -22012 2229
rect -22058 2157 -22052 2191
rect -22018 2157 -22012 2191
rect -22058 2119 -22012 2157
rect -22058 2085 -22052 2119
rect -22018 2085 -22012 2119
rect -22058 2047 -22012 2085
rect -22058 2013 -22052 2047
rect -22018 2013 -22012 2047
rect -22058 1975 -22012 2013
rect -22058 1941 -22052 1975
rect -22018 1941 -22012 1975
rect -22058 1903 -22012 1941
rect -22058 1869 -22052 1903
rect -22018 1869 -22012 1903
rect -22058 1854 -22012 1869
rect -21962 2839 -21916 2854
rect -21962 2805 -21956 2839
rect -21922 2805 -21916 2839
rect -21962 2767 -21916 2805
rect -21962 2733 -21956 2767
rect -21922 2733 -21916 2767
rect -21962 2695 -21916 2733
rect -21962 2661 -21956 2695
rect -21922 2661 -21916 2695
rect -21962 2623 -21916 2661
rect -21962 2589 -21956 2623
rect -21922 2589 -21916 2623
rect -21962 2551 -21916 2589
rect -21962 2517 -21956 2551
rect -21922 2517 -21916 2551
rect -21962 2479 -21916 2517
rect -21962 2445 -21956 2479
rect -21922 2445 -21916 2479
rect -21962 2407 -21916 2445
rect -21962 2373 -21956 2407
rect -21922 2373 -21916 2407
rect -21962 2335 -21916 2373
rect -21962 2301 -21956 2335
rect -21922 2301 -21916 2335
rect -21962 2263 -21916 2301
rect -21962 2229 -21956 2263
rect -21922 2229 -21916 2263
rect -21962 2191 -21916 2229
rect -21962 2157 -21956 2191
rect -21922 2157 -21916 2191
rect -21962 2119 -21916 2157
rect -21962 2085 -21956 2119
rect -21922 2085 -21916 2119
rect -21962 2047 -21916 2085
rect -21962 2013 -21956 2047
rect -21922 2013 -21916 2047
rect -21962 1975 -21916 2013
rect -21962 1941 -21956 1975
rect -21922 1941 -21916 1975
rect -21962 1903 -21916 1941
rect -21962 1869 -21956 1903
rect -21922 1869 -21916 1903
rect -21962 1854 -21916 1869
rect -21866 2839 -21820 2854
rect -21866 2805 -21860 2839
rect -21826 2805 -21820 2839
rect -21866 2767 -21820 2805
rect -21866 2733 -21860 2767
rect -21826 2733 -21820 2767
rect -21866 2695 -21820 2733
rect -21866 2661 -21860 2695
rect -21826 2661 -21820 2695
rect -21866 2623 -21820 2661
rect -21866 2589 -21860 2623
rect -21826 2589 -21820 2623
rect -21866 2551 -21820 2589
rect -21866 2517 -21860 2551
rect -21826 2517 -21820 2551
rect -21866 2479 -21820 2517
rect -21866 2445 -21860 2479
rect -21826 2445 -21820 2479
rect -21866 2407 -21820 2445
rect -21866 2373 -21860 2407
rect -21826 2373 -21820 2407
rect -21866 2335 -21820 2373
rect -21866 2301 -21860 2335
rect -21826 2301 -21820 2335
rect -21866 2263 -21820 2301
rect -21866 2229 -21860 2263
rect -21826 2229 -21820 2263
rect -21866 2191 -21820 2229
rect -21866 2157 -21860 2191
rect -21826 2157 -21820 2191
rect -21866 2119 -21820 2157
rect -21866 2085 -21860 2119
rect -21826 2085 -21820 2119
rect -21866 2047 -21820 2085
rect -21866 2013 -21860 2047
rect -21826 2013 -21820 2047
rect -21866 1975 -21820 2013
rect -21866 1941 -21860 1975
rect -21826 1941 -21820 1975
rect -21866 1903 -21820 1941
rect -21866 1869 -21860 1903
rect -21826 1869 -21820 1903
rect -21866 1854 -21820 1869
rect -21770 2839 -21724 2854
rect -21770 2805 -21764 2839
rect -21730 2805 -21724 2839
rect -21770 2767 -21724 2805
rect -21770 2733 -21764 2767
rect -21730 2733 -21724 2767
rect -21770 2695 -21724 2733
rect -21770 2661 -21764 2695
rect -21730 2661 -21724 2695
rect -21770 2623 -21724 2661
rect -21770 2589 -21764 2623
rect -21730 2589 -21724 2623
rect -21770 2551 -21724 2589
rect -21770 2517 -21764 2551
rect -21730 2517 -21724 2551
rect -21770 2479 -21724 2517
rect -21770 2445 -21764 2479
rect -21730 2445 -21724 2479
rect -21770 2407 -21724 2445
rect -21770 2373 -21764 2407
rect -21730 2373 -21724 2407
rect -21770 2335 -21724 2373
rect -21770 2301 -21764 2335
rect -21730 2301 -21724 2335
rect -21770 2263 -21724 2301
rect -21770 2229 -21764 2263
rect -21730 2229 -21724 2263
rect -21770 2191 -21724 2229
rect -21770 2157 -21764 2191
rect -21730 2157 -21724 2191
rect -21770 2119 -21724 2157
rect -21770 2085 -21764 2119
rect -21730 2085 -21724 2119
rect -21770 2047 -21724 2085
rect -21770 2013 -21764 2047
rect -21730 2013 -21724 2047
rect -21770 1975 -21724 2013
rect -21770 1941 -21764 1975
rect -21730 1941 -21724 1975
rect -21770 1903 -21724 1941
rect -21770 1869 -21764 1903
rect -21730 1869 -21724 1903
rect -21770 1854 -21724 1869
rect -21674 2839 -21628 2854
rect -21674 2805 -21668 2839
rect -21634 2805 -21628 2839
rect -21674 2767 -21628 2805
rect -21674 2733 -21668 2767
rect -21634 2733 -21628 2767
rect -21674 2695 -21628 2733
rect -21674 2661 -21668 2695
rect -21634 2661 -21628 2695
rect -21674 2623 -21628 2661
rect -21674 2589 -21668 2623
rect -21634 2589 -21628 2623
rect -21674 2551 -21628 2589
rect -21674 2517 -21668 2551
rect -21634 2517 -21628 2551
rect -21674 2479 -21628 2517
rect -21674 2445 -21668 2479
rect -21634 2445 -21628 2479
rect -21674 2407 -21628 2445
rect -21674 2373 -21668 2407
rect -21634 2373 -21628 2407
rect -21674 2335 -21628 2373
rect -21674 2301 -21668 2335
rect -21634 2301 -21628 2335
rect -21674 2263 -21628 2301
rect -21674 2229 -21668 2263
rect -21634 2229 -21628 2263
rect -21674 2191 -21628 2229
rect -21674 2157 -21668 2191
rect -21634 2157 -21628 2191
rect -21674 2119 -21628 2157
rect -21674 2085 -21668 2119
rect -21634 2085 -21628 2119
rect -21674 2047 -21628 2085
rect -21674 2013 -21668 2047
rect -21634 2013 -21628 2047
rect -21674 1975 -21628 2013
rect -21674 1941 -21668 1975
rect -21634 1941 -21628 1975
rect -21674 1903 -21628 1941
rect -21674 1869 -21668 1903
rect -21634 1869 -21628 1903
rect -21674 1854 -21628 1869
rect -21578 2839 -21532 2854
rect -21578 2805 -21572 2839
rect -21538 2805 -21532 2839
rect -21578 2767 -21532 2805
rect -21578 2733 -21572 2767
rect -21538 2733 -21532 2767
rect -21578 2695 -21532 2733
rect -21578 2661 -21572 2695
rect -21538 2661 -21532 2695
rect -21578 2623 -21532 2661
rect -21578 2589 -21572 2623
rect -21538 2589 -21532 2623
rect -21578 2551 -21532 2589
rect -21578 2517 -21572 2551
rect -21538 2517 -21532 2551
rect -21578 2479 -21532 2517
rect -21578 2445 -21572 2479
rect -21538 2445 -21532 2479
rect -21578 2407 -21532 2445
rect -21578 2373 -21572 2407
rect -21538 2373 -21532 2407
rect -21578 2335 -21532 2373
rect -21578 2301 -21572 2335
rect -21538 2301 -21532 2335
rect -21578 2263 -21532 2301
rect -21578 2229 -21572 2263
rect -21538 2229 -21532 2263
rect -21578 2191 -21532 2229
rect -21578 2157 -21572 2191
rect -21538 2157 -21532 2191
rect -21578 2119 -21532 2157
rect -21578 2085 -21572 2119
rect -21538 2085 -21532 2119
rect -21578 2047 -21532 2085
rect -21578 2013 -21572 2047
rect -21538 2013 -21532 2047
rect -21578 1975 -21532 2013
rect -21578 1941 -21572 1975
rect -21538 1941 -21532 1975
rect -21578 1903 -21532 1941
rect -21578 1869 -21572 1903
rect -21538 1869 -21532 1903
rect -21578 1854 -21532 1869
rect -21350 2831 -21304 2846
rect -21350 2797 -21344 2831
rect -21310 2797 -21304 2831
rect -21350 2759 -21304 2797
rect -21350 2725 -21344 2759
rect -21310 2725 -21304 2759
rect -21350 2687 -21304 2725
rect -21350 2653 -21344 2687
rect -21310 2653 -21304 2687
rect -21350 2615 -21304 2653
rect -21350 2581 -21344 2615
rect -21310 2581 -21304 2615
rect -21350 2543 -21304 2581
rect -21350 2509 -21344 2543
rect -21310 2509 -21304 2543
rect -21350 2471 -21304 2509
rect -21350 2437 -21344 2471
rect -21310 2437 -21304 2471
rect -21350 2399 -21304 2437
rect -21350 2365 -21344 2399
rect -21310 2365 -21304 2399
rect -21350 2327 -21304 2365
rect -21350 2293 -21344 2327
rect -21310 2293 -21304 2327
rect -21350 2255 -21304 2293
rect -21350 2221 -21344 2255
rect -21310 2221 -21304 2255
rect -21350 2183 -21304 2221
rect -21350 2149 -21344 2183
rect -21310 2149 -21304 2183
rect -21350 2111 -21304 2149
rect -21350 2077 -21344 2111
rect -21310 2077 -21304 2111
rect -21350 2039 -21304 2077
rect -21350 2005 -21344 2039
rect -21310 2005 -21304 2039
rect -21350 1967 -21304 2005
rect -21350 1933 -21344 1967
rect -21310 1933 -21304 1967
rect -21350 1895 -21304 1933
rect -21350 1861 -21344 1895
rect -21310 1861 -21304 1895
rect -21350 1846 -21304 1861
rect -21254 2831 -21208 2846
rect -21254 2797 -21248 2831
rect -21214 2797 -21208 2831
rect -21254 2759 -21208 2797
rect -21254 2725 -21248 2759
rect -21214 2725 -21208 2759
rect -21254 2687 -21208 2725
rect -21254 2653 -21248 2687
rect -21214 2653 -21208 2687
rect -21254 2615 -21208 2653
rect -21254 2581 -21248 2615
rect -21214 2581 -21208 2615
rect -21254 2543 -21208 2581
rect -21254 2509 -21248 2543
rect -21214 2509 -21208 2543
rect -21254 2471 -21208 2509
rect -21254 2437 -21248 2471
rect -21214 2437 -21208 2471
rect -21254 2399 -21208 2437
rect -21254 2365 -21248 2399
rect -21214 2365 -21208 2399
rect -21254 2327 -21208 2365
rect -21254 2293 -21248 2327
rect -21214 2293 -21208 2327
rect -21254 2255 -21208 2293
rect -21254 2221 -21248 2255
rect -21214 2221 -21208 2255
rect -21254 2183 -21208 2221
rect -21254 2149 -21248 2183
rect -21214 2149 -21208 2183
rect -21254 2111 -21208 2149
rect -21254 2077 -21248 2111
rect -21214 2077 -21208 2111
rect -21254 2039 -21208 2077
rect -21254 2005 -21248 2039
rect -21214 2005 -21208 2039
rect -21254 1967 -21208 2005
rect -21254 1933 -21248 1967
rect -21214 1933 -21208 1967
rect -21254 1895 -21208 1933
rect -21254 1861 -21248 1895
rect -21214 1861 -21208 1895
rect -21254 1846 -21208 1861
rect -21158 2831 -21112 2846
rect -21158 2797 -21152 2831
rect -21118 2797 -21112 2831
rect -21158 2759 -21112 2797
rect -21158 2725 -21152 2759
rect -21118 2725 -21112 2759
rect -21158 2687 -21112 2725
rect -21158 2653 -21152 2687
rect -21118 2653 -21112 2687
rect -21158 2615 -21112 2653
rect -21158 2581 -21152 2615
rect -21118 2581 -21112 2615
rect -21158 2543 -21112 2581
rect -21158 2509 -21152 2543
rect -21118 2509 -21112 2543
rect -21158 2471 -21112 2509
rect -21158 2437 -21152 2471
rect -21118 2437 -21112 2471
rect -21158 2399 -21112 2437
rect -21158 2365 -21152 2399
rect -21118 2365 -21112 2399
rect -21158 2327 -21112 2365
rect -21158 2293 -21152 2327
rect -21118 2293 -21112 2327
rect -21158 2255 -21112 2293
rect -21158 2221 -21152 2255
rect -21118 2221 -21112 2255
rect -21158 2183 -21112 2221
rect -21158 2149 -21152 2183
rect -21118 2149 -21112 2183
rect -21158 2111 -21112 2149
rect -21158 2077 -21152 2111
rect -21118 2077 -21112 2111
rect -21158 2039 -21112 2077
rect -21158 2005 -21152 2039
rect -21118 2005 -21112 2039
rect -21158 1967 -21112 2005
rect -21158 1933 -21152 1967
rect -21118 1933 -21112 1967
rect -21158 1895 -21112 1933
rect -21158 1861 -21152 1895
rect -21118 1861 -21112 1895
rect -21158 1846 -21112 1861
rect -21062 2831 -21016 2846
rect -21062 2797 -21056 2831
rect -21022 2797 -21016 2831
rect -21062 2759 -21016 2797
rect -21062 2725 -21056 2759
rect -21022 2725 -21016 2759
rect -21062 2687 -21016 2725
rect -21062 2653 -21056 2687
rect -21022 2653 -21016 2687
rect -21062 2615 -21016 2653
rect -21062 2581 -21056 2615
rect -21022 2581 -21016 2615
rect -21062 2543 -21016 2581
rect -21062 2509 -21056 2543
rect -21022 2509 -21016 2543
rect -21062 2471 -21016 2509
rect -21062 2437 -21056 2471
rect -21022 2437 -21016 2471
rect -21062 2399 -21016 2437
rect -21062 2365 -21056 2399
rect -21022 2365 -21016 2399
rect -21062 2327 -21016 2365
rect -21062 2293 -21056 2327
rect -21022 2293 -21016 2327
rect -21062 2255 -21016 2293
rect -21062 2221 -21056 2255
rect -21022 2221 -21016 2255
rect -21062 2183 -21016 2221
rect -21062 2149 -21056 2183
rect -21022 2149 -21016 2183
rect -21062 2111 -21016 2149
rect -21062 2077 -21056 2111
rect -21022 2077 -21016 2111
rect -21062 2039 -21016 2077
rect -21062 2005 -21056 2039
rect -21022 2005 -21016 2039
rect -21062 1967 -21016 2005
rect -21062 1933 -21056 1967
rect -21022 1933 -21016 1967
rect -21062 1895 -21016 1933
rect -21062 1861 -21056 1895
rect -21022 1861 -21016 1895
rect -21062 1846 -21016 1861
rect -20966 2831 -20920 2846
rect -20966 2797 -20960 2831
rect -20926 2797 -20920 2831
rect -20966 2759 -20920 2797
rect -20966 2725 -20960 2759
rect -20926 2725 -20920 2759
rect -20966 2687 -20920 2725
rect -20966 2653 -20960 2687
rect -20926 2653 -20920 2687
rect -20966 2615 -20920 2653
rect -20966 2581 -20960 2615
rect -20926 2581 -20920 2615
rect -20966 2543 -20920 2581
rect -20966 2509 -20960 2543
rect -20926 2509 -20920 2543
rect -20966 2471 -20920 2509
rect -20966 2437 -20960 2471
rect -20926 2437 -20920 2471
rect -20966 2399 -20920 2437
rect -20966 2365 -20960 2399
rect -20926 2365 -20920 2399
rect -20966 2327 -20920 2365
rect -20966 2293 -20960 2327
rect -20926 2293 -20920 2327
rect -20966 2255 -20920 2293
rect -20966 2221 -20960 2255
rect -20926 2221 -20920 2255
rect -20966 2183 -20920 2221
rect -20966 2149 -20960 2183
rect -20926 2149 -20920 2183
rect -20966 2111 -20920 2149
rect -20966 2077 -20960 2111
rect -20926 2077 -20920 2111
rect -20966 2039 -20920 2077
rect -20966 2005 -20960 2039
rect -20926 2005 -20920 2039
rect -20966 1967 -20920 2005
rect -20966 1933 -20960 1967
rect -20926 1933 -20920 1967
rect -20966 1895 -20920 1933
rect -20966 1861 -20960 1895
rect -20926 1861 -20920 1895
rect -20966 1846 -20920 1861
rect -20870 2831 -20824 2846
rect -20870 2797 -20864 2831
rect -20830 2797 -20824 2831
rect -20870 2759 -20824 2797
rect -20870 2725 -20864 2759
rect -20830 2725 -20824 2759
rect -20870 2687 -20824 2725
rect -20870 2653 -20864 2687
rect -20830 2653 -20824 2687
rect -20870 2615 -20824 2653
rect -20870 2581 -20864 2615
rect -20830 2581 -20824 2615
rect -20870 2543 -20824 2581
rect -20870 2509 -20864 2543
rect -20830 2509 -20824 2543
rect -20870 2471 -20824 2509
rect -20870 2437 -20864 2471
rect -20830 2437 -20824 2471
rect -20870 2399 -20824 2437
rect -20870 2365 -20864 2399
rect -20830 2365 -20824 2399
rect -20870 2327 -20824 2365
rect -20870 2293 -20864 2327
rect -20830 2293 -20824 2327
rect -20870 2255 -20824 2293
rect -20870 2221 -20864 2255
rect -20830 2221 -20824 2255
rect -20870 2183 -20824 2221
rect -20870 2149 -20864 2183
rect -20830 2149 -20824 2183
rect -20870 2111 -20824 2149
rect -20870 2077 -20864 2111
rect -20830 2077 -20824 2111
rect -20870 2039 -20824 2077
rect -20870 2005 -20864 2039
rect -20830 2005 -20824 2039
rect -20870 1967 -20824 2005
rect -20870 1933 -20864 1967
rect -20830 1933 -20824 1967
rect -20870 1895 -20824 1933
rect -20870 1861 -20864 1895
rect -20830 1861 -20824 1895
rect -20870 1846 -20824 1861
rect -20774 2831 -20728 2846
rect -20774 2797 -20768 2831
rect -20734 2797 -20728 2831
rect -20774 2759 -20728 2797
rect -20774 2725 -20768 2759
rect -20734 2725 -20728 2759
rect -20774 2687 -20728 2725
rect -20774 2653 -20768 2687
rect -20734 2653 -20728 2687
rect -20774 2615 -20728 2653
rect -20774 2581 -20768 2615
rect -20734 2581 -20728 2615
rect -20774 2543 -20728 2581
rect -20774 2509 -20768 2543
rect -20734 2509 -20728 2543
rect -20774 2471 -20728 2509
rect -20774 2437 -20768 2471
rect -20734 2437 -20728 2471
rect -20774 2399 -20728 2437
rect -20774 2365 -20768 2399
rect -20734 2365 -20728 2399
rect -20774 2327 -20728 2365
rect -20774 2293 -20768 2327
rect -20734 2293 -20728 2327
rect -20774 2255 -20728 2293
rect -20774 2221 -20768 2255
rect -20734 2221 -20728 2255
rect -20774 2183 -20728 2221
rect -20774 2149 -20768 2183
rect -20734 2149 -20728 2183
rect -20774 2111 -20728 2149
rect -20774 2077 -20768 2111
rect -20734 2077 -20728 2111
rect -20774 2039 -20728 2077
rect -20774 2005 -20768 2039
rect -20734 2005 -20728 2039
rect -20774 1967 -20728 2005
rect -20774 1933 -20768 1967
rect -20734 1933 -20728 1967
rect -20774 1895 -20728 1933
rect -20774 1861 -20768 1895
rect -20734 1861 -20728 1895
rect -20774 1846 -20728 1861
rect -20678 2831 -20632 2846
rect -20678 2797 -20672 2831
rect -20638 2797 -20632 2831
rect -20678 2759 -20632 2797
rect -20678 2725 -20672 2759
rect -20638 2725 -20632 2759
rect -20678 2687 -20632 2725
rect -20678 2653 -20672 2687
rect -20638 2653 -20632 2687
rect -20678 2615 -20632 2653
rect -20678 2581 -20672 2615
rect -20638 2581 -20632 2615
rect -20678 2543 -20632 2581
rect -20678 2509 -20672 2543
rect -20638 2509 -20632 2543
rect -20678 2471 -20632 2509
rect -20678 2437 -20672 2471
rect -20638 2437 -20632 2471
rect -20678 2399 -20632 2437
rect -20678 2365 -20672 2399
rect -20638 2365 -20632 2399
rect -20678 2327 -20632 2365
rect -20678 2293 -20672 2327
rect -20638 2293 -20632 2327
rect -20678 2255 -20632 2293
rect -20678 2221 -20672 2255
rect -20638 2221 -20632 2255
rect -20678 2183 -20632 2221
rect -20678 2149 -20672 2183
rect -20638 2149 -20632 2183
rect -20678 2111 -20632 2149
rect -20678 2077 -20672 2111
rect -20638 2077 -20632 2111
rect -20678 2039 -20632 2077
rect -20678 2005 -20672 2039
rect -20638 2005 -20632 2039
rect -20678 1967 -20632 2005
rect -20678 1933 -20672 1967
rect -20638 1933 -20632 1967
rect -20678 1895 -20632 1933
rect -20678 1861 -20672 1895
rect -20638 1861 -20632 1895
rect -20678 1846 -20632 1861
rect -20582 2831 -20536 2846
rect -20582 2797 -20576 2831
rect -20542 2797 -20536 2831
rect -20582 2759 -20536 2797
rect -20582 2725 -20576 2759
rect -20542 2725 -20536 2759
rect -20582 2687 -20536 2725
rect -20582 2653 -20576 2687
rect -20542 2653 -20536 2687
rect -20582 2615 -20536 2653
rect -20582 2581 -20576 2615
rect -20542 2581 -20536 2615
rect -20582 2543 -20536 2581
rect -20582 2509 -20576 2543
rect -20542 2509 -20536 2543
rect -20582 2471 -20536 2509
rect -20582 2437 -20576 2471
rect -20542 2437 -20536 2471
rect -20582 2399 -20536 2437
rect -20582 2365 -20576 2399
rect -20542 2365 -20536 2399
rect -20582 2327 -20536 2365
rect -20582 2293 -20576 2327
rect -20542 2293 -20536 2327
rect -20582 2255 -20536 2293
rect -20582 2221 -20576 2255
rect -20542 2221 -20536 2255
rect -20582 2183 -20536 2221
rect -20582 2149 -20576 2183
rect -20542 2149 -20536 2183
rect -20582 2111 -20536 2149
rect -20582 2077 -20576 2111
rect -20542 2077 -20536 2111
rect -20582 2039 -20536 2077
rect -20582 2005 -20576 2039
rect -20542 2005 -20536 2039
rect -20582 1967 -20536 2005
rect -20582 1933 -20576 1967
rect -20542 1933 -20536 1967
rect -20582 1895 -20536 1933
rect -20582 1861 -20576 1895
rect -20542 1861 -20536 1895
rect -20582 1846 -20536 1861
rect -20486 2831 -20440 2846
rect -20486 2797 -20480 2831
rect -20446 2797 -20440 2831
rect -20486 2759 -20440 2797
rect -20486 2725 -20480 2759
rect -20446 2725 -20440 2759
rect -20486 2687 -20440 2725
rect -20486 2653 -20480 2687
rect -20446 2653 -20440 2687
rect -20486 2615 -20440 2653
rect -20486 2581 -20480 2615
rect -20446 2581 -20440 2615
rect -20486 2543 -20440 2581
rect -20486 2509 -20480 2543
rect -20446 2509 -20440 2543
rect -20486 2471 -20440 2509
rect -20486 2437 -20480 2471
rect -20446 2437 -20440 2471
rect -20486 2399 -20440 2437
rect -20486 2365 -20480 2399
rect -20446 2365 -20440 2399
rect -20486 2327 -20440 2365
rect -20486 2293 -20480 2327
rect -20446 2293 -20440 2327
rect -20486 2255 -20440 2293
rect -20486 2221 -20480 2255
rect -20446 2221 -20440 2255
rect -20486 2183 -20440 2221
rect -20486 2149 -20480 2183
rect -20446 2149 -20440 2183
rect -20486 2111 -20440 2149
rect -20486 2077 -20480 2111
rect -20446 2077 -20440 2111
rect -20486 2039 -20440 2077
rect -20486 2005 -20480 2039
rect -20446 2005 -20440 2039
rect -20486 1967 -20440 2005
rect -20486 1933 -20480 1967
rect -20446 1933 -20440 1967
rect -20486 1895 -20440 1933
rect -20486 1861 -20480 1895
rect -20446 1861 -20440 1895
rect -20486 1846 -20440 1861
rect -20390 2831 -20344 2846
rect -20390 2797 -20384 2831
rect -20350 2797 -20344 2831
rect -20390 2759 -20344 2797
rect -20390 2725 -20384 2759
rect -20350 2725 -20344 2759
rect -20390 2687 -20344 2725
rect -20390 2653 -20384 2687
rect -20350 2653 -20344 2687
rect -20390 2615 -20344 2653
rect -20390 2581 -20384 2615
rect -20350 2581 -20344 2615
rect -20390 2543 -20344 2581
rect -20390 2509 -20384 2543
rect -20350 2509 -20344 2543
rect -20390 2471 -20344 2509
rect -20390 2437 -20384 2471
rect -20350 2437 -20344 2471
rect -20390 2399 -20344 2437
rect -20390 2365 -20384 2399
rect -20350 2365 -20344 2399
rect -20390 2327 -20344 2365
rect -20390 2293 -20384 2327
rect -20350 2293 -20344 2327
rect -20390 2255 -20344 2293
rect -20390 2221 -20384 2255
rect -20350 2221 -20344 2255
rect -20390 2183 -20344 2221
rect -20390 2149 -20384 2183
rect -20350 2149 -20344 2183
rect -20390 2111 -20344 2149
rect -20390 2077 -20384 2111
rect -20350 2077 -20344 2111
rect -20390 2039 -20344 2077
rect -20390 2005 -20384 2039
rect -20350 2005 -20344 2039
rect -20390 1967 -20344 2005
rect -20390 1933 -20384 1967
rect -20350 1933 -20344 1967
rect -20390 1895 -20344 1933
rect -20390 1861 -20384 1895
rect -20350 1861 -20344 1895
rect -20390 1846 -20344 1861
rect -20294 2831 -20248 2846
rect -20294 2797 -20288 2831
rect -20254 2797 -20248 2831
rect -20294 2759 -20248 2797
rect -20294 2725 -20288 2759
rect -20254 2725 -20248 2759
rect -20294 2687 -20248 2725
rect -20294 2653 -20288 2687
rect -20254 2653 -20248 2687
rect -20294 2615 -20248 2653
rect -20294 2581 -20288 2615
rect -20254 2581 -20248 2615
rect -20294 2543 -20248 2581
rect -20294 2509 -20288 2543
rect -20254 2509 -20248 2543
rect -20294 2471 -20248 2509
rect -20294 2437 -20288 2471
rect -20254 2437 -20248 2471
rect -20294 2399 -20248 2437
rect -20294 2365 -20288 2399
rect -20254 2365 -20248 2399
rect -20294 2327 -20248 2365
rect -20294 2293 -20288 2327
rect -20254 2293 -20248 2327
rect -20294 2255 -20248 2293
rect -20294 2221 -20288 2255
rect -20254 2221 -20248 2255
rect -20294 2183 -20248 2221
rect -20294 2149 -20288 2183
rect -20254 2149 -20248 2183
rect -20294 2111 -20248 2149
rect -20294 2077 -20288 2111
rect -20254 2077 -20248 2111
rect -20294 2039 -20248 2077
rect -20294 2005 -20288 2039
rect -20254 2005 -20248 2039
rect -20294 1967 -20248 2005
rect -20294 1933 -20288 1967
rect -20254 1933 -20248 1967
rect -20294 1895 -20248 1933
rect -20294 1861 -20288 1895
rect -20254 1861 -20248 1895
rect -20294 1846 -20248 1861
rect -20198 2831 -20152 2846
rect -20198 2797 -20192 2831
rect -20158 2797 -20152 2831
rect -20198 2759 -20152 2797
rect -20198 2725 -20192 2759
rect -20158 2725 -20152 2759
rect -20198 2687 -20152 2725
rect -20198 2653 -20192 2687
rect -20158 2653 -20152 2687
rect -20198 2615 -20152 2653
rect -20198 2581 -20192 2615
rect -20158 2581 -20152 2615
rect -20198 2543 -20152 2581
rect -20198 2509 -20192 2543
rect -20158 2509 -20152 2543
rect -20198 2471 -20152 2509
rect -20198 2437 -20192 2471
rect -20158 2437 -20152 2471
rect -20198 2399 -20152 2437
rect -20198 2365 -20192 2399
rect -20158 2365 -20152 2399
rect -20198 2327 -20152 2365
rect -20198 2293 -20192 2327
rect -20158 2293 -20152 2327
rect -20198 2255 -20152 2293
rect -20198 2221 -20192 2255
rect -20158 2221 -20152 2255
rect -20198 2183 -20152 2221
rect -20198 2149 -20192 2183
rect -20158 2149 -20152 2183
rect -20198 2111 -20152 2149
rect -20198 2077 -20192 2111
rect -20158 2077 -20152 2111
rect -20198 2039 -20152 2077
rect -20198 2005 -20192 2039
rect -20158 2005 -20152 2039
rect -20198 1967 -20152 2005
rect -20198 1933 -20192 1967
rect -20158 1933 -20152 1967
rect -20198 1895 -20152 1933
rect -20198 1861 -20192 1895
rect -20158 1861 -20152 1895
rect -20198 1846 -20152 1861
rect -20102 2831 -20056 2846
rect -20102 2797 -20096 2831
rect -20062 2797 -20056 2831
rect -20102 2759 -20056 2797
rect -20102 2725 -20096 2759
rect -20062 2725 -20056 2759
rect -20102 2687 -20056 2725
rect -20102 2653 -20096 2687
rect -20062 2653 -20056 2687
rect -20102 2615 -20056 2653
rect -20102 2581 -20096 2615
rect -20062 2581 -20056 2615
rect -20102 2543 -20056 2581
rect -20102 2509 -20096 2543
rect -20062 2509 -20056 2543
rect -20102 2471 -20056 2509
rect -20102 2437 -20096 2471
rect -20062 2437 -20056 2471
rect -20102 2399 -20056 2437
rect -20102 2365 -20096 2399
rect -20062 2365 -20056 2399
rect -20102 2327 -20056 2365
rect -20102 2293 -20096 2327
rect -20062 2293 -20056 2327
rect -20102 2255 -20056 2293
rect -20102 2221 -20096 2255
rect -20062 2221 -20056 2255
rect -20102 2183 -20056 2221
rect -20102 2149 -20096 2183
rect -20062 2149 -20056 2183
rect -20102 2111 -20056 2149
rect -20102 2077 -20096 2111
rect -20062 2077 -20056 2111
rect -20102 2039 -20056 2077
rect -20102 2005 -20096 2039
rect -20062 2005 -20056 2039
rect -20102 1967 -20056 2005
rect -20102 1933 -20096 1967
rect -20062 1933 -20056 1967
rect -20102 1895 -20056 1933
rect -20102 1861 -20096 1895
rect -20062 1861 -20056 1895
rect -20102 1846 -20056 1861
rect -20006 2831 -19960 2846
rect -20006 2797 -20000 2831
rect -19966 2797 -19960 2831
rect -20006 2759 -19960 2797
rect -20006 2725 -20000 2759
rect -19966 2725 -19960 2759
rect -20006 2687 -19960 2725
rect -20006 2653 -20000 2687
rect -19966 2653 -19960 2687
rect -20006 2615 -19960 2653
rect -20006 2581 -20000 2615
rect -19966 2581 -19960 2615
rect -20006 2543 -19960 2581
rect -20006 2509 -20000 2543
rect -19966 2509 -19960 2543
rect -20006 2471 -19960 2509
rect -20006 2437 -20000 2471
rect -19966 2437 -19960 2471
rect -20006 2399 -19960 2437
rect -20006 2365 -20000 2399
rect -19966 2365 -19960 2399
rect -20006 2327 -19960 2365
rect -20006 2293 -20000 2327
rect -19966 2293 -19960 2327
rect -20006 2255 -19960 2293
rect -20006 2221 -20000 2255
rect -19966 2221 -19960 2255
rect -20006 2183 -19960 2221
rect -20006 2149 -20000 2183
rect -19966 2149 -19960 2183
rect -20006 2111 -19960 2149
rect -20006 2077 -20000 2111
rect -19966 2077 -19960 2111
rect -20006 2039 -19960 2077
rect -20006 2005 -20000 2039
rect -19966 2005 -19960 2039
rect -20006 1967 -19960 2005
rect -20006 1933 -20000 1967
rect -19966 1933 -19960 1967
rect -20006 1895 -19960 1933
rect -20006 1861 -20000 1895
rect -19966 1861 -19960 1895
rect -20006 1846 -19960 1861
rect -19910 2831 -19864 2846
rect -19910 2797 -19904 2831
rect -19870 2797 -19864 2831
rect -19910 2759 -19864 2797
rect -19910 2725 -19904 2759
rect -19870 2725 -19864 2759
rect -19910 2687 -19864 2725
rect -19910 2653 -19904 2687
rect -19870 2653 -19864 2687
rect -19910 2615 -19864 2653
rect -19910 2581 -19904 2615
rect -19870 2581 -19864 2615
rect -19910 2543 -19864 2581
rect -19910 2509 -19904 2543
rect -19870 2509 -19864 2543
rect -19910 2471 -19864 2509
rect -19910 2437 -19904 2471
rect -19870 2437 -19864 2471
rect -19910 2399 -19864 2437
rect -19910 2365 -19904 2399
rect -19870 2365 -19864 2399
rect -19910 2327 -19864 2365
rect -19910 2293 -19904 2327
rect -19870 2293 -19864 2327
rect -19910 2255 -19864 2293
rect -19910 2221 -19904 2255
rect -19870 2221 -19864 2255
rect -19910 2183 -19864 2221
rect -19910 2149 -19904 2183
rect -19870 2149 -19864 2183
rect -19910 2111 -19864 2149
rect -19910 2077 -19904 2111
rect -19870 2077 -19864 2111
rect -19910 2039 -19864 2077
rect -19910 2005 -19904 2039
rect -19870 2005 -19864 2039
rect -19910 1967 -19864 2005
rect -19910 1933 -19904 1967
rect -19870 1933 -19864 1967
rect -19910 1895 -19864 1933
rect -19910 1861 -19904 1895
rect -19870 1861 -19864 1895
rect -19910 1846 -19864 1861
rect -19672 2835 -19626 2850
rect -19672 2801 -19666 2835
rect -19632 2801 -19626 2835
rect -19672 2763 -19626 2801
rect -19672 2729 -19666 2763
rect -19632 2729 -19626 2763
rect -19672 2691 -19626 2729
rect -19672 2657 -19666 2691
rect -19632 2657 -19626 2691
rect -19672 2619 -19626 2657
rect -19672 2585 -19666 2619
rect -19632 2585 -19626 2619
rect -19672 2547 -19626 2585
rect -19672 2513 -19666 2547
rect -19632 2513 -19626 2547
rect -19672 2475 -19626 2513
rect -19672 2441 -19666 2475
rect -19632 2441 -19626 2475
rect -19672 2403 -19626 2441
rect -19672 2369 -19666 2403
rect -19632 2369 -19626 2403
rect -19672 2331 -19626 2369
rect -19672 2297 -19666 2331
rect -19632 2297 -19626 2331
rect -19672 2259 -19626 2297
rect -19672 2225 -19666 2259
rect -19632 2225 -19626 2259
rect -19672 2187 -19626 2225
rect -19672 2153 -19666 2187
rect -19632 2153 -19626 2187
rect -19672 2115 -19626 2153
rect -19672 2081 -19666 2115
rect -19632 2081 -19626 2115
rect -19672 2043 -19626 2081
rect -19672 2009 -19666 2043
rect -19632 2009 -19626 2043
rect -19672 1971 -19626 2009
rect -19672 1937 -19666 1971
rect -19632 1937 -19626 1971
rect -19672 1899 -19626 1937
rect -19672 1865 -19666 1899
rect -19632 1865 -19626 1899
rect -19672 1850 -19626 1865
rect -19576 2835 -19530 2850
rect -19576 2801 -19570 2835
rect -19536 2801 -19530 2835
rect -19576 2763 -19530 2801
rect -19576 2729 -19570 2763
rect -19536 2729 -19530 2763
rect -19576 2691 -19530 2729
rect -19576 2657 -19570 2691
rect -19536 2657 -19530 2691
rect -19576 2619 -19530 2657
rect -19576 2585 -19570 2619
rect -19536 2585 -19530 2619
rect -19576 2547 -19530 2585
rect -19576 2513 -19570 2547
rect -19536 2513 -19530 2547
rect -19576 2475 -19530 2513
rect -19576 2441 -19570 2475
rect -19536 2441 -19530 2475
rect -19576 2403 -19530 2441
rect -19576 2369 -19570 2403
rect -19536 2369 -19530 2403
rect -19576 2331 -19530 2369
rect -19576 2297 -19570 2331
rect -19536 2297 -19530 2331
rect -19576 2259 -19530 2297
rect -19576 2225 -19570 2259
rect -19536 2225 -19530 2259
rect -19576 2187 -19530 2225
rect -19576 2153 -19570 2187
rect -19536 2153 -19530 2187
rect -19576 2115 -19530 2153
rect -19576 2081 -19570 2115
rect -19536 2081 -19530 2115
rect -19576 2043 -19530 2081
rect -19576 2009 -19570 2043
rect -19536 2009 -19530 2043
rect -19576 1971 -19530 2009
rect -19576 1937 -19570 1971
rect -19536 1937 -19530 1971
rect -19576 1899 -19530 1937
rect -19576 1865 -19570 1899
rect -19536 1865 -19530 1899
rect -19576 1850 -19530 1865
rect -19480 2835 -19434 2850
rect -19480 2801 -19474 2835
rect -19440 2801 -19434 2835
rect -19480 2763 -19434 2801
rect -19480 2729 -19474 2763
rect -19440 2729 -19434 2763
rect -19480 2691 -19434 2729
rect -19480 2657 -19474 2691
rect -19440 2657 -19434 2691
rect -19480 2619 -19434 2657
rect -19480 2585 -19474 2619
rect -19440 2585 -19434 2619
rect -19480 2547 -19434 2585
rect -19480 2513 -19474 2547
rect -19440 2513 -19434 2547
rect -19480 2475 -19434 2513
rect -19480 2441 -19474 2475
rect -19440 2441 -19434 2475
rect -19480 2403 -19434 2441
rect -19480 2369 -19474 2403
rect -19440 2369 -19434 2403
rect -19480 2331 -19434 2369
rect -19480 2297 -19474 2331
rect -19440 2297 -19434 2331
rect -19480 2259 -19434 2297
rect -19480 2225 -19474 2259
rect -19440 2225 -19434 2259
rect -19480 2187 -19434 2225
rect -19480 2153 -19474 2187
rect -19440 2153 -19434 2187
rect -19480 2115 -19434 2153
rect -19480 2081 -19474 2115
rect -19440 2081 -19434 2115
rect -19480 2043 -19434 2081
rect -19480 2009 -19474 2043
rect -19440 2009 -19434 2043
rect -19480 1971 -19434 2009
rect -19480 1937 -19474 1971
rect -19440 1937 -19434 1971
rect -19480 1899 -19434 1937
rect -19480 1865 -19474 1899
rect -19440 1865 -19434 1899
rect -19480 1850 -19434 1865
rect -19384 2835 -19338 2850
rect -19384 2801 -19378 2835
rect -19344 2801 -19338 2835
rect -19384 2763 -19338 2801
rect -19384 2729 -19378 2763
rect -19344 2729 -19338 2763
rect -19384 2691 -19338 2729
rect -19384 2657 -19378 2691
rect -19344 2657 -19338 2691
rect -19384 2619 -19338 2657
rect -19384 2585 -19378 2619
rect -19344 2585 -19338 2619
rect -19384 2547 -19338 2585
rect -19384 2513 -19378 2547
rect -19344 2513 -19338 2547
rect -19384 2475 -19338 2513
rect -19384 2441 -19378 2475
rect -19344 2441 -19338 2475
rect -19384 2403 -19338 2441
rect -19384 2369 -19378 2403
rect -19344 2369 -19338 2403
rect -19384 2331 -19338 2369
rect -19384 2297 -19378 2331
rect -19344 2297 -19338 2331
rect -19384 2259 -19338 2297
rect -19384 2225 -19378 2259
rect -19344 2225 -19338 2259
rect -19384 2187 -19338 2225
rect -19384 2153 -19378 2187
rect -19344 2153 -19338 2187
rect -19384 2115 -19338 2153
rect -19384 2081 -19378 2115
rect -19344 2081 -19338 2115
rect -19384 2043 -19338 2081
rect -19384 2009 -19378 2043
rect -19344 2009 -19338 2043
rect -19384 1971 -19338 2009
rect -19384 1937 -19378 1971
rect -19344 1937 -19338 1971
rect -19384 1899 -19338 1937
rect -19384 1865 -19378 1899
rect -19344 1865 -19338 1899
rect -19384 1850 -19338 1865
rect -19288 2835 -19242 2850
rect -19288 2801 -19282 2835
rect -19248 2801 -19242 2835
rect -19288 2763 -19242 2801
rect -19288 2729 -19282 2763
rect -19248 2729 -19242 2763
rect -19288 2691 -19242 2729
rect -19288 2657 -19282 2691
rect -19248 2657 -19242 2691
rect -19288 2619 -19242 2657
rect -19288 2585 -19282 2619
rect -19248 2585 -19242 2619
rect -19288 2547 -19242 2585
rect -19288 2513 -19282 2547
rect -19248 2513 -19242 2547
rect -19288 2475 -19242 2513
rect -19288 2441 -19282 2475
rect -19248 2441 -19242 2475
rect -19288 2403 -19242 2441
rect -19288 2369 -19282 2403
rect -19248 2369 -19242 2403
rect -19288 2331 -19242 2369
rect -19288 2297 -19282 2331
rect -19248 2297 -19242 2331
rect -19288 2259 -19242 2297
rect -19288 2225 -19282 2259
rect -19248 2225 -19242 2259
rect -19288 2187 -19242 2225
rect -19288 2153 -19282 2187
rect -19248 2153 -19242 2187
rect -19288 2115 -19242 2153
rect -19288 2081 -19282 2115
rect -19248 2081 -19242 2115
rect -19288 2043 -19242 2081
rect -19288 2009 -19282 2043
rect -19248 2009 -19242 2043
rect -19288 1971 -19242 2009
rect -19288 1937 -19282 1971
rect -19248 1937 -19242 1971
rect -19288 1899 -19242 1937
rect -19288 1865 -19282 1899
rect -19248 1865 -19242 1899
rect -19288 1850 -19242 1865
rect -19192 2835 -19146 2850
rect -19192 2801 -19186 2835
rect -19152 2801 -19146 2835
rect -19192 2763 -19146 2801
rect -19192 2729 -19186 2763
rect -19152 2729 -19146 2763
rect -19192 2691 -19146 2729
rect -19192 2657 -19186 2691
rect -19152 2657 -19146 2691
rect -19192 2619 -19146 2657
rect -19192 2585 -19186 2619
rect -19152 2585 -19146 2619
rect -19192 2547 -19146 2585
rect -19192 2513 -19186 2547
rect -19152 2513 -19146 2547
rect -19192 2475 -19146 2513
rect -19192 2441 -19186 2475
rect -19152 2441 -19146 2475
rect -19192 2403 -19146 2441
rect -19192 2369 -19186 2403
rect -19152 2369 -19146 2403
rect -19192 2331 -19146 2369
rect -19192 2297 -19186 2331
rect -19152 2297 -19146 2331
rect -19192 2259 -19146 2297
rect -19192 2225 -19186 2259
rect -19152 2225 -19146 2259
rect -19192 2187 -19146 2225
rect -19192 2153 -19186 2187
rect -19152 2153 -19146 2187
rect -19192 2115 -19146 2153
rect -19192 2081 -19186 2115
rect -19152 2081 -19146 2115
rect -19192 2043 -19146 2081
rect -19192 2009 -19186 2043
rect -19152 2009 -19146 2043
rect -19192 1971 -19146 2009
rect -19192 1937 -19186 1971
rect -19152 1937 -19146 1971
rect -19192 1899 -19146 1937
rect -19192 1865 -19186 1899
rect -19152 1865 -19146 1899
rect -19192 1850 -19146 1865
rect -19096 2835 -19050 2850
rect -19096 2801 -19090 2835
rect -19056 2801 -19050 2835
rect -19096 2763 -19050 2801
rect -19096 2729 -19090 2763
rect -19056 2729 -19050 2763
rect -19096 2691 -19050 2729
rect -19096 2657 -19090 2691
rect -19056 2657 -19050 2691
rect -19096 2619 -19050 2657
rect -19096 2585 -19090 2619
rect -19056 2585 -19050 2619
rect -19096 2547 -19050 2585
rect -19096 2513 -19090 2547
rect -19056 2513 -19050 2547
rect -19096 2475 -19050 2513
rect -19096 2441 -19090 2475
rect -19056 2441 -19050 2475
rect -19096 2403 -19050 2441
rect -19096 2369 -19090 2403
rect -19056 2369 -19050 2403
rect -19096 2331 -19050 2369
rect -19096 2297 -19090 2331
rect -19056 2297 -19050 2331
rect -19096 2259 -19050 2297
rect -19096 2225 -19090 2259
rect -19056 2225 -19050 2259
rect -19096 2187 -19050 2225
rect -19096 2153 -19090 2187
rect -19056 2153 -19050 2187
rect -19096 2115 -19050 2153
rect -19096 2081 -19090 2115
rect -19056 2081 -19050 2115
rect -19096 2043 -19050 2081
rect -19096 2009 -19090 2043
rect -19056 2009 -19050 2043
rect -19096 1971 -19050 2009
rect -19096 1937 -19090 1971
rect -19056 1937 -19050 1971
rect -19096 1899 -19050 1937
rect -19096 1865 -19090 1899
rect -19056 1865 -19050 1899
rect -19096 1850 -19050 1865
rect -19000 2835 -18954 2850
rect -19000 2801 -18994 2835
rect -18960 2801 -18954 2835
rect -19000 2763 -18954 2801
rect -19000 2729 -18994 2763
rect -18960 2729 -18954 2763
rect -19000 2691 -18954 2729
rect -19000 2657 -18994 2691
rect -18960 2657 -18954 2691
rect -19000 2619 -18954 2657
rect -19000 2585 -18994 2619
rect -18960 2585 -18954 2619
rect -19000 2547 -18954 2585
rect -19000 2513 -18994 2547
rect -18960 2513 -18954 2547
rect -19000 2475 -18954 2513
rect -19000 2441 -18994 2475
rect -18960 2441 -18954 2475
rect -19000 2403 -18954 2441
rect -19000 2369 -18994 2403
rect -18960 2369 -18954 2403
rect -19000 2331 -18954 2369
rect -19000 2297 -18994 2331
rect -18960 2297 -18954 2331
rect -19000 2259 -18954 2297
rect -19000 2225 -18994 2259
rect -18960 2225 -18954 2259
rect -19000 2187 -18954 2225
rect -19000 2153 -18994 2187
rect -18960 2153 -18954 2187
rect -19000 2115 -18954 2153
rect -19000 2081 -18994 2115
rect -18960 2081 -18954 2115
rect -19000 2043 -18954 2081
rect -19000 2009 -18994 2043
rect -18960 2009 -18954 2043
rect -19000 1971 -18954 2009
rect -19000 1937 -18994 1971
rect -18960 1937 -18954 1971
rect -19000 1899 -18954 1937
rect -19000 1865 -18994 1899
rect -18960 1865 -18954 1899
rect -19000 1850 -18954 1865
rect -18904 2835 -18858 2850
rect -18904 2801 -18898 2835
rect -18864 2801 -18858 2835
rect -18904 2763 -18858 2801
rect -18904 2729 -18898 2763
rect -18864 2729 -18858 2763
rect -18904 2691 -18858 2729
rect -18904 2657 -18898 2691
rect -18864 2657 -18858 2691
rect -18904 2619 -18858 2657
rect -18904 2585 -18898 2619
rect -18864 2585 -18858 2619
rect -18904 2547 -18858 2585
rect -18904 2513 -18898 2547
rect -18864 2513 -18858 2547
rect -18904 2475 -18858 2513
rect -18904 2441 -18898 2475
rect -18864 2441 -18858 2475
rect -18904 2403 -18858 2441
rect -18904 2369 -18898 2403
rect -18864 2369 -18858 2403
rect -18904 2331 -18858 2369
rect -18904 2297 -18898 2331
rect -18864 2297 -18858 2331
rect -18904 2259 -18858 2297
rect -18904 2225 -18898 2259
rect -18864 2225 -18858 2259
rect -18904 2187 -18858 2225
rect -18904 2153 -18898 2187
rect -18864 2153 -18858 2187
rect -18904 2115 -18858 2153
rect -18904 2081 -18898 2115
rect -18864 2081 -18858 2115
rect -18904 2043 -18858 2081
rect -18904 2009 -18898 2043
rect -18864 2009 -18858 2043
rect -18904 1971 -18858 2009
rect -18904 1937 -18898 1971
rect -18864 1937 -18858 1971
rect -18904 1899 -18858 1937
rect -18904 1865 -18898 1899
rect -18864 1865 -18858 1899
rect -18904 1850 -18858 1865
rect -18808 2835 -18762 2850
rect -18808 2801 -18802 2835
rect -18768 2801 -18762 2835
rect -18808 2763 -18762 2801
rect -18808 2729 -18802 2763
rect -18768 2729 -18762 2763
rect -18808 2691 -18762 2729
rect -18808 2657 -18802 2691
rect -18768 2657 -18762 2691
rect -18808 2619 -18762 2657
rect -18808 2585 -18802 2619
rect -18768 2585 -18762 2619
rect -18808 2547 -18762 2585
rect -18808 2513 -18802 2547
rect -18768 2513 -18762 2547
rect -18808 2475 -18762 2513
rect -18808 2441 -18802 2475
rect -18768 2441 -18762 2475
rect -18808 2403 -18762 2441
rect -18808 2369 -18802 2403
rect -18768 2369 -18762 2403
rect -18808 2331 -18762 2369
rect -18808 2297 -18802 2331
rect -18768 2297 -18762 2331
rect -18808 2259 -18762 2297
rect -18808 2225 -18802 2259
rect -18768 2225 -18762 2259
rect -18808 2187 -18762 2225
rect -18808 2153 -18802 2187
rect -18768 2153 -18762 2187
rect -18808 2115 -18762 2153
rect -18808 2081 -18802 2115
rect -18768 2081 -18762 2115
rect -18808 2043 -18762 2081
rect -18808 2009 -18802 2043
rect -18768 2009 -18762 2043
rect -18808 1971 -18762 2009
rect -18808 1937 -18802 1971
rect -18768 1937 -18762 1971
rect -18808 1899 -18762 1937
rect -18808 1865 -18802 1899
rect -18768 1865 -18762 1899
rect -18808 1850 -18762 1865
rect -18712 2835 -18666 2850
rect -18712 2801 -18706 2835
rect -18672 2801 -18666 2835
rect -18712 2763 -18666 2801
rect -18712 2729 -18706 2763
rect -18672 2729 -18666 2763
rect -18712 2691 -18666 2729
rect -18712 2657 -18706 2691
rect -18672 2657 -18666 2691
rect -18712 2619 -18666 2657
rect -18712 2585 -18706 2619
rect -18672 2585 -18666 2619
rect -18712 2547 -18666 2585
rect -18712 2513 -18706 2547
rect -18672 2513 -18666 2547
rect -18712 2475 -18666 2513
rect -18712 2441 -18706 2475
rect -18672 2441 -18666 2475
rect -18712 2403 -18666 2441
rect -18712 2369 -18706 2403
rect -18672 2369 -18666 2403
rect -18712 2331 -18666 2369
rect -18712 2297 -18706 2331
rect -18672 2297 -18666 2331
rect -18712 2259 -18666 2297
rect -18712 2225 -18706 2259
rect -18672 2225 -18666 2259
rect -18712 2187 -18666 2225
rect -18712 2153 -18706 2187
rect -18672 2153 -18666 2187
rect -18712 2115 -18666 2153
rect -18712 2081 -18706 2115
rect -18672 2081 -18666 2115
rect -18712 2043 -18666 2081
rect -18712 2009 -18706 2043
rect -18672 2009 -18666 2043
rect -18712 1971 -18666 2009
rect -18712 1937 -18706 1971
rect -18672 1937 -18666 1971
rect -18712 1899 -18666 1937
rect -18712 1865 -18706 1899
rect -18672 1865 -18666 1899
rect -18712 1850 -18666 1865
rect -18500 2845 -18454 2860
rect -18500 2811 -18494 2845
rect -18460 2811 -18454 2845
rect -18500 2773 -18454 2811
rect -18500 2739 -18494 2773
rect -18460 2739 -18454 2773
rect -18500 2701 -18454 2739
rect -18500 2667 -18494 2701
rect -18460 2667 -18454 2701
rect -18500 2629 -18454 2667
rect -18500 2595 -18494 2629
rect -18460 2595 -18454 2629
rect -18500 2557 -18454 2595
rect -18500 2523 -18494 2557
rect -18460 2523 -18454 2557
rect -18500 2485 -18454 2523
rect -18500 2451 -18494 2485
rect -18460 2451 -18454 2485
rect -18500 2413 -18454 2451
rect -18500 2379 -18494 2413
rect -18460 2379 -18454 2413
rect -18500 2341 -18454 2379
rect -18500 2307 -18494 2341
rect -18460 2307 -18454 2341
rect -18500 2269 -18454 2307
rect -18500 2235 -18494 2269
rect -18460 2235 -18454 2269
rect -18500 2197 -18454 2235
rect -18500 2163 -18494 2197
rect -18460 2163 -18454 2197
rect -18500 2125 -18454 2163
rect -18500 2091 -18494 2125
rect -18460 2091 -18454 2125
rect -18500 2053 -18454 2091
rect -18500 2019 -18494 2053
rect -18460 2019 -18454 2053
rect -18500 1981 -18454 2019
rect -18500 1947 -18494 1981
rect -18460 1947 -18454 1981
rect -18500 1909 -18454 1947
rect -18500 1875 -18494 1909
rect -18460 1875 -18454 1909
rect -18500 1860 -18454 1875
rect -18404 2845 -18358 2860
rect -18404 2811 -18398 2845
rect -18364 2811 -18358 2845
rect -18404 2773 -18358 2811
rect -18404 2739 -18398 2773
rect -18364 2739 -18358 2773
rect -18404 2701 -18358 2739
rect -18404 2667 -18398 2701
rect -18364 2667 -18358 2701
rect -18404 2629 -18358 2667
rect -18404 2595 -18398 2629
rect -18364 2595 -18358 2629
rect -18404 2557 -18358 2595
rect -18404 2523 -18398 2557
rect -18364 2523 -18358 2557
rect -18404 2485 -18358 2523
rect -18404 2451 -18398 2485
rect -18364 2451 -18358 2485
rect -18404 2413 -18358 2451
rect -18404 2379 -18398 2413
rect -18364 2379 -18358 2413
rect -18404 2341 -18358 2379
rect -18404 2307 -18398 2341
rect -18364 2307 -18358 2341
rect -18404 2269 -18358 2307
rect -18404 2235 -18398 2269
rect -18364 2235 -18358 2269
rect -18404 2197 -18358 2235
rect -18404 2163 -18398 2197
rect -18364 2163 -18358 2197
rect -18404 2125 -18358 2163
rect -18404 2091 -18398 2125
rect -18364 2091 -18358 2125
rect -18404 2053 -18358 2091
rect -18404 2019 -18398 2053
rect -18364 2019 -18358 2053
rect -18404 1981 -18358 2019
rect -18404 1947 -18398 1981
rect -18364 1947 -18358 1981
rect -18404 1909 -18358 1947
rect -18404 1875 -18398 1909
rect -18364 1875 -18358 1909
rect -18404 1860 -18358 1875
rect -18308 2845 -18262 2860
rect -18308 2811 -18302 2845
rect -18268 2811 -18262 2845
rect -18308 2773 -18262 2811
rect -18308 2739 -18302 2773
rect -18268 2739 -18262 2773
rect -18308 2701 -18262 2739
rect -18308 2667 -18302 2701
rect -18268 2667 -18262 2701
rect -18308 2629 -18262 2667
rect -18308 2595 -18302 2629
rect -18268 2595 -18262 2629
rect -18308 2557 -18262 2595
rect -18308 2523 -18302 2557
rect -18268 2523 -18262 2557
rect -18308 2485 -18262 2523
rect -18308 2451 -18302 2485
rect -18268 2451 -18262 2485
rect -18308 2413 -18262 2451
rect -18308 2379 -18302 2413
rect -18268 2379 -18262 2413
rect -18308 2341 -18262 2379
rect -18308 2307 -18302 2341
rect -18268 2307 -18262 2341
rect -18308 2269 -18262 2307
rect -18308 2235 -18302 2269
rect -18268 2235 -18262 2269
rect -18308 2197 -18262 2235
rect -18308 2163 -18302 2197
rect -18268 2163 -18262 2197
rect -18308 2125 -18262 2163
rect -18308 2091 -18302 2125
rect -18268 2091 -18262 2125
rect -18308 2053 -18262 2091
rect -18308 2019 -18302 2053
rect -18268 2019 -18262 2053
rect -18308 1981 -18262 2019
rect -18308 1947 -18302 1981
rect -18268 1947 -18262 1981
rect -18308 1909 -18262 1947
rect -18308 1875 -18302 1909
rect -18268 1875 -18262 1909
rect -18308 1860 -18262 1875
rect -18212 2845 -18166 2860
rect -18212 2811 -18206 2845
rect -18172 2811 -18166 2845
rect -18212 2773 -18166 2811
rect -18212 2739 -18206 2773
rect -18172 2739 -18166 2773
rect -18212 2701 -18166 2739
rect -18212 2667 -18206 2701
rect -18172 2667 -18166 2701
rect -18212 2629 -18166 2667
rect -18212 2595 -18206 2629
rect -18172 2595 -18166 2629
rect -18212 2557 -18166 2595
rect -18212 2523 -18206 2557
rect -18172 2523 -18166 2557
rect -18212 2485 -18166 2523
rect -18212 2451 -18206 2485
rect -18172 2451 -18166 2485
rect -18212 2413 -18166 2451
rect -18212 2379 -18206 2413
rect -18172 2379 -18166 2413
rect -18212 2341 -18166 2379
rect -18212 2307 -18206 2341
rect -18172 2307 -18166 2341
rect -18212 2269 -18166 2307
rect -18212 2235 -18206 2269
rect -18172 2235 -18166 2269
rect -18212 2197 -18166 2235
rect -18212 2163 -18206 2197
rect -18172 2163 -18166 2197
rect -18212 2125 -18166 2163
rect -18212 2091 -18206 2125
rect -18172 2091 -18166 2125
rect -18212 2053 -18166 2091
rect -18212 2019 -18206 2053
rect -18172 2019 -18166 2053
rect -18212 1981 -18166 2019
rect -18212 1947 -18206 1981
rect -18172 1947 -18166 1981
rect -18212 1909 -18166 1947
rect -18212 1875 -18206 1909
rect -18172 1875 -18166 1909
rect -18212 1860 -18166 1875
rect -18116 2845 -18070 2860
rect -18116 2811 -18110 2845
rect -18076 2811 -18070 2845
rect -18116 2773 -18070 2811
rect -18116 2739 -18110 2773
rect -18076 2739 -18070 2773
rect -18116 2701 -18070 2739
rect -18116 2667 -18110 2701
rect -18076 2667 -18070 2701
rect -18116 2629 -18070 2667
rect -18116 2595 -18110 2629
rect -18076 2595 -18070 2629
rect -18116 2557 -18070 2595
rect -18116 2523 -18110 2557
rect -18076 2523 -18070 2557
rect -18116 2485 -18070 2523
rect -18116 2451 -18110 2485
rect -18076 2451 -18070 2485
rect -18116 2413 -18070 2451
rect -18116 2379 -18110 2413
rect -18076 2379 -18070 2413
rect -18116 2341 -18070 2379
rect -18116 2307 -18110 2341
rect -18076 2307 -18070 2341
rect -18116 2269 -18070 2307
rect -18116 2235 -18110 2269
rect -18076 2235 -18070 2269
rect -18116 2197 -18070 2235
rect -18116 2163 -18110 2197
rect -18076 2163 -18070 2197
rect -18116 2125 -18070 2163
rect -18116 2091 -18110 2125
rect -18076 2091 -18070 2125
rect -18116 2053 -18070 2091
rect -18116 2019 -18110 2053
rect -18076 2019 -18070 2053
rect -18116 1981 -18070 2019
rect -18116 1947 -18110 1981
rect -18076 1947 -18070 1981
rect -18116 1909 -18070 1947
rect -18116 1875 -18110 1909
rect -18076 1875 -18070 1909
rect -18116 1860 -18070 1875
rect -18020 2845 -17974 2860
rect -18020 2811 -18014 2845
rect -17980 2811 -17974 2845
rect -18020 2773 -17974 2811
rect -18020 2739 -18014 2773
rect -17980 2739 -17974 2773
rect -18020 2701 -17974 2739
rect -18020 2667 -18014 2701
rect -17980 2667 -17974 2701
rect -18020 2629 -17974 2667
rect -18020 2595 -18014 2629
rect -17980 2595 -17974 2629
rect -18020 2557 -17974 2595
rect -18020 2523 -18014 2557
rect -17980 2523 -17974 2557
rect -18020 2485 -17974 2523
rect -18020 2451 -18014 2485
rect -17980 2451 -17974 2485
rect -18020 2413 -17974 2451
rect -18020 2379 -18014 2413
rect -17980 2379 -17974 2413
rect -18020 2341 -17974 2379
rect -18020 2307 -18014 2341
rect -17980 2307 -17974 2341
rect -18020 2269 -17974 2307
rect -18020 2235 -18014 2269
rect -17980 2235 -17974 2269
rect -18020 2197 -17974 2235
rect -18020 2163 -18014 2197
rect -17980 2163 -17974 2197
rect -18020 2125 -17974 2163
rect -18020 2091 -18014 2125
rect -17980 2091 -17974 2125
rect -18020 2053 -17974 2091
rect -18020 2019 -18014 2053
rect -17980 2019 -17974 2053
rect -18020 1981 -17974 2019
rect -18020 1947 -18014 1981
rect -17980 1947 -17974 1981
rect -18020 1909 -17974 1947
rect -18020 1875 -18014 1909
rect -17980 1875 -17974 1909
rect -18020 1860 -17974 1875
rect -23126 1665 -22748 1668
rect -19126 1666 -18748 1668
rect -23126 1485 -23091 1665
rect -22783 1485 -22748 1665
rect -23126 1482 -22748 1485
rect -21126 1664 -20748 1666
rect -21126 1484 -21091 1664
rect -20783 1484 -20748 1664
rect -19126 1486 -19091 1666
rect -18783 1486 -18748 1666
rect -19126 1484 -18748 1486
rect -21126 1482 -20748 1484
rect -17380 -5888 -17074 3090
rect -14924 3086 -13854 3110
rect -13252 3157 -12200 3188
rect -13252 3123 -12288 3157
rect -12254 3123 -12200 3157
rect -13252 3092 -12200 3123
rect -12042 3178 -11962 3265
rect -11358 3281 -11260 3308
rect -11358 3247 -11328 3281
rect -11294 3247 -11260 3281
rect -11358 3184 -11260 3247
rect -8458 3285 -8346 3330
rect -8458 3251 -8418 3285
rect -8384 3251 -8346 3285
rect -12042 3159 -11410 3178
rect -12042 3125 -11472 3159
rect -11438 3125 -11410 3159
rect -12042 3108 -11410 3125
rect -11358 3158 -10914 3184
rect -8458 3168 -8346 3251
rect -6786 3291 -6686 3322
rect -6786 3257 -6754 3291
rect -6720 3257 -6686 3291
rect -6786 3186 -6686 3257
rect -5576 3297 -5496 3328
rect -5576 3263 -5550 3297
rect -5516 3263 -5496 3297
rect -14924 3028 -14812 3086
rect -14924 2994 -14886 3028
rect -14852 2994 -14812 3028
rect -14924 2954 -14812 2994
rect -13252 3030 -13152 3092
rect -13252 2996 -13218 3030
rect -13184 2996 -13152 3030
rect -12042 3074 -11962 3108
rect -12042 3040 -12020 3074
rect -11986 3040 -11962 3074
rect -12042 3018 -11962 3040
rect -11358 3106 -11002 3158
rect -10950 3106 -10914 3158
rect -11358 3080 -10914 3106
rect -10698 3140 -9588 3160
rect -10698 3106 -9678 3140
rect -9644 3106 -9588 3140
rect -10698 3088 -9588 3106
rect -8458 3142 -7388 3168
rect -8458 3108 -7475 3142
rect -7441 3108 -7388 3142
rect -10698 3086 -10368 3088
rect -11358 3044 -11260 3080
rect -13252 2970 -13152 2996
rect -11358 3010 -11328 3044
rect -11294 3010 -11260 3044
rect -11358 2984 -11260 3010
rect -16668 2851 -16622 2866
rect -16668 2817 -16662 2851
rect -16628 2817 -16622 2851
rect -16668 2779 -16622 2817
rect -16668 2745 -16662 2779
rect -16628 2745 -16622 2779
rect -16668 2707 -16622 2745
rect -16668 2673 -16662 2707
rect -16628 2673 -16622 2707
rect -16668 2635 -16622 2673
rect -16668 2601 -16662 2635
rect -16628 2601 -16622 2635
rect -16668 2563 -16622 2601
rect -16668 2529 -16662 2563
rect -16628 2529 -16622 2563
rect -16668 2491 -16622 2529
rect -16668 2457 -16662 2491
rect -16628 2457 -16622 2491
rect -16668 2419 -16622 2457
rect -16668 2385 -16662 2419
rect -16628 2385 -16622 2419
rect -16668 2347 -16622 2385
rect -16668 2313 -16662 2347
rect -16628 2313 -16622 2347
rect -16668 2275 -16622 2313
rect -16668 2241 -16662 2275
rect -16628 2241 -16622 2275
rect -16668 2203 -16622 2241
rect -16668 2169 -16662 2203
rect -16628 2169 -16622 2203
rect -16668 2131 -16622 2169
rect -16668 2097 -16662 2131
rect -16628 2097 -16622 2131
rect -16668 2059 -16622 2097
rect -16668 2025 -16662 2059
rect -16628 2025 -16622 2059
rect -16668 1987 -16622 2025
rect -16668 1953 -16662 1987
rect -16628 1953 -16622 1987
rect -16668 1915 -16622 1953
rect -16668 1881 -16662 1915
rect -16628 1881 -16622 1915
rect -16668 1866 -16622 1881
rect -16572 2851 -16526 2866
rect -16572 2817 -16566 2851
rect -16532 2817 -16526 2851
rect -16572 2779 -16526 2817
rect -16572 2745 -16566 2779
rect -16532 2745 -16526 2779
rect -16572 2707 -16526 2745
rect -16572 2673 -16566 2707
rect -16532 2673 -16526 2707
rect -16572 2635 -16526 2673
rect -16572 2601 -16566 2635
rect -16532 2601 -16526 2635
rect -16572 2563 -16526 2601
rect -16572 2529 -16566 2563
rect -16532 2529 -16526 2563
rect -16572 2491 -16526 2529
rect -16572 2457 -16566 2491
rect -16532 2457 -16526 2491
rect -16572 2419 -16526 2457
rect -16572 2385 -16566 2419
rect -16532 2385 -16526 2419
rect -16572 2347 -16526 2385
rect -16572 2313 -16566 2347
rect -16532 2313 -16526 2347
rect -16572 2275 -16526 2313
rect -16572 2241 -16566 2275
rect -16532 2241 -16526 2275
rect -16572 2203 -16526 2241
rect -16572 2169 -16566 2203
rect -16532 2169 -16526 2203
rect -16572 2131 -16526 2169
rect -16572 2097 -16566 2131
rect -16532 2097 -16526 2131
rect -16572 2059 -16526 2097
rect -16572 2025 -16566 2059
rect -16532 2025 -16526 2059
rect -16572 1987 -16526 2025
rect -16572 1953 -16566 1987
rect -16532 1953 -16526 1987
rect -16572 1915 -16526 1953
rect -16572 1881 -16566 1915
rect -16532 1881 -16526 1915
rect -16572 1866 -16526 1881
rect -16476 2851 -16430 2866
rect -16476 2817 -16470 2851
rect -16436 2817 -16430 2851
rect -16476 2779 -16430 2817
rect -16476 2745 -16470 2779
rect -16436 2745 -16430 2779
rect -16476 2707 -16430 2745
rect -16476 2673 -16470 2707
rect -16436 2673 -16430 2707
rect -16476 2635 -16430 2673
rect -16476 2601 -16470 2635
rect -16436 2601 -16430 2635
rect -16476 2563 -16430 2601
rect -16476 2529 -16470 2563
rect -16436 2529 -16430 2563
rect -16476 2491 -16430 2529
rect -16476 2457 -16470 2491
rect -16436 2457 -16430 2491
rect -16476 2419 -16430 2457
rect -16476 2385 -16470 2419
rect -16436 2385 -16430 2419
rect -16476 2347 -16430 2385
rect -16476 2313 -16470 2347
rect -16436 2313 -16430 2347
rect -16476 2275 -16430 2313
rect -16476 2241 -16470 2275
rect -16436 2241 -16430 2275
rect -16476 2203 -16430 2241
rect -16476 2169 -16470 2203
rect -16436 2169 -16430 2203
rect -16476 2131 -16430 2169
rect -16476 2097 -16470 2131
rect -16436 2097 -16430 2131
rect -16476 2059 -16430 2097
rect -16476 2025 -16470 2059
rect -16436 2025 -16430 2059
rect -16476 1987 -16430 2025
rect -16476 1953 -16470 1987
rect -16436 1953 -16430 1987
rect -16476 1915 -16430 1953
rect -16476 1881 -16470 1915
rect -16436 1881 -16430 1915
rect -16476 1866 -16430 1881
rect -16380 2851 -16334 2866
rect -16380 2817 -16374 2851
rect -16340 2817 -16334 2851
rect -16380 2779 -16334 2817
rect -16380 2745 -16374 2779
rect -16340 2745 -16334 2779
rect -16380 2707 -16334 2745
rect -16380 2673 -16374 2707
rect -16340 2673 -16334 2707
rect -16380 2635 -16334 2673
rect -16380 2601 -16374 2635
rect -16340 2601 -16334 2635
rect -16380 2563 -16334 2601
rect -16380 2529 -16374 2563
rect -16340 2529 -16334 2563
rect -16380 2491 -16334 2529
rect -16380 2457 -16374 2491
rect -16340 2457 -16334 2491
rect -16380 2419 -16334 2457
rect -16380 2385 -16374 2419
rect -16340 2385 -16334 2419
rect -16380 2347 -16334 2385
rect -16380 2313 -16374 2347
rect -16340 2313 -16334 2347
rect -16380 2275 -16334 2313
rect -16380 2241 -16374 2275
rect -16340 2241 -16334 2275
rect -16380 2203 -16334 2241
rect -16380 2169 -16374 2203
rect -16340 2169 -16334 2203
rect -16380 2131 -16334 2169
rect -16380 2097 -16374 2131
rect -16340 2097 -16334 2131
rect -16380 2059 -16334 2097
rect -16380 2025 -16374 2059
rect -16340 2025 -16334 2059
rect -16380 1987 -16334 2025
rect -16380 1953 -16374 1987
rect -16340 1953 -16334 1987
rect -16380 1915 -16334 1953
rect -16380 1881 -16374 1915
rect -16340 1881 -16334 1915
rect -16380 1866 -16334 1881
rect -16284 2851 -16238 2866
rect -16284 2817 -16278 2851
rect -16244 2817 -16238 2851
rect -16284 2779 -16238 2817
rect -16284 2745 -16278 2779
rect -16244 2745 -16238 2779
rect -16284 2707 -16238 2745
rect -16284 2673 -16278 2707
rect -16244 2673 -16238 2707
rect -16284 2635 -16238 2673
rect -16284 2601 -16278 2635
rect -16244 2601 -16238 2635
rect -16284 2563 -16238 2601
rect -16284 2529 -16278 2563
rect -16244 2529 -16238 2563
rect -16284 2491 -16238 2529
rect -16284 2457 -16278 2491
rect -16244 2457 -16238 2491
rect -16284 2419 -16238 2457
rect -16284 2385 -16278 2419
rect -16244 2385 -16238 2419
rect -16284 2347 -16238 2385
rect -16284 2313 -16278 2347
rect -16244 2313 -16238 2347
rect -16284 2275 -16238 2313
rect -16284 2241 -16278 2275
rect -16244 2241 -16238 2275
rect -16284 2203 -16238 2241
rect -16284 2169 -16278 2203
rect -16244 2169 -16238 2203
rect -16284 2131 -16238 2169
rect -16284 2097 -16278 2131
rect -16244 2097 -16238 2131
rect -16284 2059 -16238 2097
rect -16284 2025 -16278 2059
rect -16244 2025 -16238 2059
rect -16284 1987 -16238 2025
rect -16284 1953 -16278 1987
rect -16244 1953 -16238 1987
rect -16284 1915 -16238 1953
rect -16284 1881 -16278 1915
rect -16244 1881 -16238 1915
rect -16284 1866 -16238 1881
rect -16188 2851 -16142 2866
rect -16188 2817 -16182 2851
rect -16148 2817 -16142 2851
rect -16188 2779 -16142 2817
rect -16188 2745 -16182 2779
rect -16148 2745 -16142 2779
rect -16188 2707 -16142 2745
rect -16188 2673 -16182 2707
rect -16148 2673 -16142 2707
rect -16188 2635 -16142 2673
rect -16188 2601 -16182 2635
rect -16148 2601 -16142 2635
rect -16188 2563 -16142 2601
rect -16188 2529 -16182 2563
rect -16148 2529 -16142 2563
rect -16188 2491 -16142 2529
rect -16188 2457 -16182 2491
rect -16148 2457 -16142 2491
rect -16188 2419 -16142 2457
rect -16188 2385 -16182 2419
rect -16148 2385 -16142 2419
rect -16188 2347 -16142 2385
rect -16188 2313 -16182 2347
rect -16148 2313 -16142 2347
rect -16188 2275 -16142 2313
rect -16188 2241 -16182 2275
rect -16148 2241 -16142 2275
rect -16188 2203 -16142 2241
rect -16188 2169 -16182 2203
rect -16148 2169 -16142 2203
rect -16188 2131 -16142 2169
rect -16188 2097 -16182 2131
rect -16148 2097 -16142 2131
rect -16188 2059 -16142 2097
rect -16188 2025 -16182 2059
rect -16148 2025 -16142 2059
rect -16188 1987 -16142 2025
rect -16188 1953 -16182 1987
rect -16148 1953 -16142 1987
rect -16188 1915 -16142 1953
rect -16188 1881 -16182 1915
rect -16148 1881 -16142 1915
rect -16188 1866 -16142 1881
rect -16092 2851 -16046 2866
rect -16092 2817 -16086 2851
rect -16052 2817 -16046 2851
rect -16092 2779 -16046 2817
rect -16092 2745 -16086 2779
rect -16052 2745 -16046 2779
rect -16092 2707 -16046 2745
rect -16092 2673 -16086 2707
rect -16052 2673 -16046 2707
rect -16092 2635 -16046 2673
rect -16092 2601 -16086 2635
rect -16052 2601 -16046 2635
rect -16092 2563 -16046 2601
rect -16092 2529 -16086 2563
rect -16052 2529 -16046 2563
rect -16092 2491 -16046 2529
rect -16092 2457 -16086 2491
rect -16052 2457 -16046 2491
rect -16092 2419 -16046 2457
rect -16092 2385 -16086 2419
rect -16052 2385 -16046 2419
rect -16092 2347 -16046 2385
rect -16092 2313 -16086 2347
rect -16052 2313 -16046 2347
rect -16092 2275 -16046 2313
rect -16092 2241 -16086 2275
rect -16052 2241 -16046 2275
rect -16092 2203 -16046 2241
rect -16092 2169 -16086 2203
rect -16052 2169 -16046 2203
rect -16092 2131 -16046 2169
rect -16092 2097 -16086 2131
rect -16052 2097 -16046 2131
rect -16092 2059 -16046 2097
rect -16092 2025 -16086 2059
rect -16052 2025 -16046 2059
rect -16092 1987 -16046 2025
rect -16092 1953 -16086 1987
rect -16052 1953 -16046 1987
rect -16092 1915 -16046 1953
rect -16092 1881 -16086 1915
rect -16052 1881 -16046 1915
rect -16092 1866 -16046 1881
rect -15996 2851 -15950 2866
rect -15996 2817 -15990 2851
rect -15956 2817 -15950 2851
rect -15996 2779 -15950 2817
rect -15996 2745 -15990 2779
rect -15956 2745 -15950 2779
rect -15996 2707 -15950 2745
rect -15996 2673 -15990 2707
rect -15956 2673 -15950 2707
rect -15996 2635 -15950 2673
rect -15996 2601 -15990 2635
rect -15956 2601 -15950 2635
rect -15996 2563 -15950 2601
rect -15996 2529 -15990 2563
rect -15956 2529 -15950 2563
rect -15996 2491 -15950 2529
rect -15996 2457 -15990 2491
rect -15956 2457 -15950 2491
rect -15996 2419 -15950 2457
rect -15996 2385 -15990 2419
rect -15956 2385 -15950 2419
rect -15996 2347 -15950 2385
rect -15996 2313 -15990 2347
rect -15956 2313 -15950 2347
rect -15996 2275 -15950 2313
rect -15996 2241 -15990 2275
rect -15956 2241 -15950 2275
rect -15996 2203 -15950 2241
rect -15996 2169 -15990 2203
rect -15956 2169 -15950 2203
rect -15996 2131 -15950 2169
rect -15996 2097 -15990 2131
rect -15956 2097 -15950 2131
rect -15996 2059 -15950 2097
rect -15996 2025 -15990 2059
rect -15956 2025 -15950 2059
rect -15996 1987 -15950 2025
rect -15996 1953 -15990 1987
rect -15956 1953 -15950 1987
rect -15996 1915 -15950 1953
rect -15996 1881 -15990 1915
rect -15956 1881 -15950 1915
rect -15996 1866 -15950 1881
rect -15900 2851 -15854 2866
rect -15900 2817 -15894 2851
rect -15860 2817 -15854 2851
rect -15900 2779 -15854 2817
rect -15900 2745 -15894 2779
rect -15860 2745 -15854 2779
rect -15900 2707 -15854 2745
rect -15900 2673 -15894 2707
rect -15860 2673 -15854 2707
rect -15900 2635 -15854 2673
rect -15900 2601 -15894 2635
rect -15860 2601 -15854 2635
rect -15900 2563 -15854 2601
rect -15900 2529 -15894 2563
rect -15860 2529 -15854 2563
rect -15900 2491 -15854 2529
rect -15900 2457 -15894 2491
rect -15860 2457 -15854 2491
rect -15900 2419 -15854 2457
rect -15900 2385 -15894 2419
rect -15860 2385 -15854 2419
rect -15900 2347 -15854 2385
rect -15900 2313 -15894 2347
rect -15860 2313 -15854 2347
rect -15900 2275 -15854 2313
rect -15900 2241 -15894 2275
rect -15860 2241 -15854 2275
rect -15900 2203 -15854 2241
rect -15900 2169 -15894 2203
rect -15860 2169 -15854 2203
rect -15900 2131 -15854 2169
rect -15900 2097 -15894 2131
rect -15860 2097 -15854 2131
rect -15900 2059 -15854 2097
rect -15900 2025 -15894 2059
rect -15860 2025 -15854 2059
rect -15900 1987 -15854 2025
rect -15900 1953 -15894 1987
rect -15860 1953 -15854 1987
rect -15900 1915 -15854 1953
rect -15900 1881 -15894 1915
rect -15860 1881 -15854 1915
rect -15900 1866 -15854 1881
rect -15804 2851 -15758 2866
rect -15804 2817 -15798 2851
rect -15764 2817 -15758 2851
rect -15804 2779 -15758 2817
rect -15804 2745 -15798 2779
rect -15764 2745 -15758 2779
rect -15804 2707 -15758 2745
rect -15804 2673 -15798 2707
rect -15764 2673 -15758 2707
rect -15804 2635 -15758 2673
rect -15804 2601 -15798 2635
rect -15764 2601 -15758 2635
rect -15804 2563 -15758 2601
rect -15804 2529 -15798 2563
rect -15764 2529 -15758 2563
rect -15804 2491 -15758 2529
rect -15804 2457 -15798 2491
rect -15764 2457 -15758 2491
rect -15804 2419 -15758 2457
rect -15804 2385 -15798 2419
rect -15764 2385 -15758 2419
rect -15804 2347 -15758 2385
rect -15804 2313 -15798 2347
rect -15764 2313 -15758 2347
rect -15804 2275 -15758 2313
rect -15804 2241 -15798 2275
rect -15764 2241 -15758 2275
rect -15804 2203 -15758 2241
rect -15804 2169 -15798 2203
rect -15764 2169 -15758 2203
rect -15804 2131 -15758 2169
rect -15804 2097 -15798 2131
rect -15764 2097 -15758 2131
rect -15804 2059 -15758 2097
rect -15804 2025 -15798 2059
rect -15764 2025 -15758 2059
rect -15804 1987 -15758 2025
rect -15804 1953 -15798 1987
rect -15764 1953 -15758 1987
rect -15804 1915 -15758 1953
rect -15804 1881 -15798 1915
rect -15764 1881 -15758 1915
rect -15804 1866 -15758 1881
rect -15708 2851 -15662 2866
rect -15708 2817 -15702 2851
rect -15668 2817 -15662 2851
rect -15708 2779 -15662 2817
rect -15708 2745 -15702 2779
rect -15668 2745 -15662 2779
rect -15708 2707 -15662 2745
rect -15708 2673 -15702 2707
rect -15668 2673 -15662 2707
rect -15708 2635 -15662 2673
rect -15708 2601 -15702 2635
rect -15668 2601 -15662 2635
rect -15708 2563 -15662 2601
rect -15708 2529 -15702 2563
rect -15668 2529 -15662 2563
rect -15708 2491 -15662 2529
rect -15708 2457 -15702 2491
rect -15668 2457 -15662 2491
rect -15708 2419 -15662 2457
rect -15708 2385 -15702 2419
rect -15668 2385 -15662 2419
rect -15708 2347 -15662 2385
rect -15708 2313 -15702 2347
rect -15668 2313 -15662 2347
rect -15708 2275 -15662 2313
rect -15708 2241 -15702 2275
rect -15668 2241 -15662 2275
rect -15708 2203 -15662 2241
rect -15708 2169 -15702 2203
rect -15668 2169 -15662 2203
rect -15708 2131 -15662 2169
rect -15708 2097 -15702 2131
rect -15668 2097 -15662 2131
rect -15708 2059 -15662 2097
rect -15708 2025 -15702 2059
rect -15668 2025 -15662 2059
rect -15708 1987 -15662 2025
rect -15708 1953 -15702 1987
rect -15668 1953 -15662 1987
rect -15708 1915 -15662 1953
rect -15708 1881 -15702 1915
rect -15668 1881 -15662 1915
rect -15708 1866 -15662 1881
rect -15612 2851 -15566 2866
rect -15612 2817 -15606 2851
rect -15572 2817 -15566 2851
rect -15612 2779 -15566 2817
rect -15612 2745 -15606 2779
rect -15572 2745 -15566 2779
rect -15612 2707 -15566 2745
rect -15612 2673 -15606 2707
rect -15572 2673 -15566 2707
rect -15612 2635 -15566 2673
rect -15612 2601 -15606 2635
rect -15572 2601 -15566 2635
rect -15612 2563 -15566 2601
rect -15612 2529 -15606 2563
rect -15572 2529 -15566 2563
rect -15612 2491 -15566 2529
rect -15612 2457 -15606 2491
rect -15572 2457 -15566 2491
rect -15612 2419 -15566 2457
rect -15612 2385 -15606 2419
rect -15572 2385 -15566 2419
rect -15612 2347 -15566 2385
rect -15612 2313 -15606 2347
rect -15572 2313 -15566 2347
rect -15612 2275 -15566 2313
rect -15612 2241 -15606 2275
rect -15572 2241 -15566 2275
rect -15612 2203 -15566 2241
rect -15612 2169 -15606 2203
rect -15572 2169 -15566 2203
rect -15612 2131 -15566 2169
rect -15612 2097 -15606 2131
rect -15572 2097 -15566 2131
rect -15612 2059 -15566 2097
rect -15612 2025 -15606 2059
rect -15572 2025 -15566 2059
rect -15612 1987 -15566 2025
rect -15612 1953 -15606 1987
rect -15572 1953 -15566 1987
rect -15612 1915 -15566 1953
rect -15612 1881 -15606 1915
rect -15572 1881 -15566 1915
rect -15612 1866 -15566 1881
rect -15516 2851 -15470 2866
rect -15516 2817 -15510 2851
rect -15476 2817 -15470 2851
rect -15516 2779 -15470 2817
rect -15516 2745 -15510 2779
rect -15476 2745 -15470 2779
rect -15516 2707 -15470 2745
rect -15516 2673 -15510 2707
rect -15476 2673 -15470 2707
rect -15516 2635 -15470 2673
rect -15516 2601 -15510 2635
rect -15476 2601 -15470 2635
rect -15516 2563 -15470 2601
rect -15516 2529 -15510 2563
rect -15476 2529 -15470 2563
rect -15516 2491 -15470 2529
rect -15516 2457 -15510 2491
rect -15476 2457 -15470 2491
rect -15516 2419 -15470 2457
rect -15516 2385 -15510 2419
rect -15476 2385 -15470 2419
rect -15516 2347 -15470 2385
rect -15516 2313 -15510 2347
rect -15476 2313 -15470 2347
rect -15516 2275 -15470 2313
rect -15516 2241 -15510 2275
rect -15476 2241 -15470 2275
rect -15516 2203 -15470 2241
rect -15516 2169 -15510 2203
rect -15476 2169 -15470 2203
rect -15516 2131 -15470 2169
rect -15516 2097 -15510 2131
rect -15476 2097 -15470 2131
rect -15516 2059 -15470 2097
rect -15516 2025 -15510 2059
rect -15476 2025 -15470 2059
rect -15516 1987 -15470 2025
rect -15516 1953 -15510 1987
rect -15476 1953 -15470 1987
rect -15516 1915 -15470 1953
rect -15516 1881 -15510 1915
rect -15476 1881 -15470 1915
rect -15516 1866 -15470 1881
rect -15420 2851 -15374 2866
rect -15420 2817 -15414 2851
rect -15380 2817 -15374 2851
rect -15420 2779 -15374 2817
rect -15420 2745 -15414 2779
rect -15380 2745 -15374 2779
rect -15420 2707 -15374 2745
rect -15420 2673 -15414 2707
rect -15380 2673 -15374 2707
rect -15420 2635 -15374 2673
rect -15420 2601 -15414 2635
rect -15380 2601 -15374 2635
rect -15420 2563 -15374 2601
rect -15420 2529 -15414 2563
rect -15380 2529 -15374 2563
rect -15420 2491 -15374 2529
rect -15420 2457 -15414 2491
rect -15380 2457 -15374 2491
rect -15420 2419 -15374 2457
rect -15420 2385 -15414 2419
rect -15380 2385 -15374 2419
rect -15420 2347 -15374 2385
rect -15420 2313 -15414 2347
rect -15380 2313 -15374 2347
rect -15420 2275 -15374 2313
rect -15420 2241 -15414 2275
rect -15380 2241 -15374 2275
rect -15420 2203 -15374 2241
rect -15420 2169 -15414 2203
rect -15380 2169 -15374 2203
rect -15420 2131 -15374 2169
rect -15420 2097 -15414 2131
rect -15380 2097 -15374 2131
rect -15420 2059 -15374 2097
rect -15420 2025 -15414 2059
rect -15380 2025 -15374 2059
rect -15420 1987 -15374 2025
rect -15420 1953 -15414 1987
rect -15380 1953 -15374 1987
rect -15420 1915 -15374 1953
rect -15420 1881 -15414 1915
rect -15380 1881 -15374 1915
rect -15420 1866 -15374 1881
rect -15324 2851 -15278 2866
rect -15324 2817 -15318 2851
rect -15284 2817 -15278 2851
rect -15324 2779 -15278 2817
rect -15324 2745 -15318 2779
rect -15284 2745 -15278 2779
rect -15324 2707 -15278 2745
rect -15324 2673 -15318 2707
rect -15284 2673 -15278 2707
rect -15324 2635 -15278 2673
rect -15324 2601 -15318 2635
rect -15284 2601 -15278 2635
rect -15324 2563 -15278 2601
rect -15324 2529 -15318 2563
rect -15284 2529 -15278 2563
rect -15324 2491 -15278 2529
rect -15324 2457 -15318 2491
rect -15284 2457 -15278 2491
rect -15324 2419 -15278 2457
rect -15324 2385 -15318 2419
rect -15284 2385 -15278 2419
rect -15324 2347 -15278 2385
rect -15324 2313 -15318 2347
rect -15284 2313 -15278 2347
rect -15324 2275 -15278 2313
rect -15324 2241 -15318 2275
rect -15284 2241 -15278 2275
rect -15324 2203 -15278 2241
rect -15324 2169 -15318 2203
rect -15284 2169 -15278 2203
rect -15324 2131 -15278 2169
rect -15324 2097 -15318 2131
rect -15284 2097 -15278 2131
rect -15324 2059 -15278 2097
rect -15324 2025 -15318 2059
rect -15284 2025 -15278 2059
rect -15324 1987 -15278 2025
rect -15324 1953 -15318 1987
rect -15284 1953 -15278 1987
rect -15324 1915 -15278 1953
rect -15324 1881 -15318 1915
rect -15284 1881 -15278 1915
rect -15324 1866 -15278 1881
rect -15228 2851 -15182 2866
rect -15228 2817 -15222 2851
rect -15188 2817 -15182 2851
rect -15228 2779 -15182 2817
rect -15228 2745 -15222 2779
rect -15188 2745 -15182 2779
rect -15228 2707 -15182 2745
rect -15228 2673 -15222 2707
rect -15188 2673 -15182 2707
rect -15228 2635 -15182 2673
rect -15228 2601 -15222 2635
rect -15188 2601 -15182 2635
rect -15228 2563 -15182 2601
rect -15228 2529 -15222 2563
rect -15188 2529 -15182 2563
rect -15228 2491 -15182 2529
rect -15228 2457 -15222 2491
rect -15188 2457 -15182 2491
rect -15228 2419 -15182 2457
rect -15228 2385 -15222 2419
rect -15188 2385 -15182 2419
rect -15228 2347 -15182 2385
rect -15228 2313 -15222 2347
rect -15188 2313 -15182 2347
rect -15228 2275 -15182 2313
rect -15228 2241 -15222 2275
rect -15188 2241 -15182 2275
rect -15228 2203 -15182 2241
rect -15228 2169 -15222 2203
rect -15188 2169 -15182 2203
rect -15228 2131 -15182 2169
rect -15228 2097 -15222 2131
rect -15188 2097 -15182 2131
rect -15228 2059 -15182 2097
rect -15228 2025 -15222 2059
rect -15188 2025 -15182 2059
rect -15228 1987 -15182 2025
rect -15228 1953 -15222 1987
rect -15188 1953 -15182 1987
rect -15228 1915 -15182 1953
rect -15228 1881 -15222 1915
rect -15188 1881 -15182 1915
rect -15228 1866 -15182 1881
rect -15132 2851 -15086 2866
rect -15132 2817 -15126 2851
rect -15092 2817 -15086 2851
rect -15132 2779 -15086 2817
rect -15132 2745 -15126 2779
rect -15092 2745 -15086 2779
rect -15132 2707 -15086 2745
rect -15132 2673 -15126 2707
rect -15092 2673 -15086 2707
rect -15132 2635 -15086 2673
rect -15132 2601 -15126 2635
rect -15092 2601 -15086 2635
rect -15132 2563 -15086 2601
rect -15132 2529 -15126 2563
rect -15092 2529 -15086 2563
rect -15132 2491 -15086 2529
rect -15132 2457 -15126 2491
rect -15092 2457 -15086 2491
rect -15132 2419 -15086 2457
rect -15132 2385 -15126 2419
rect -15092 2385 -15086 2419
rect -15132 2347 -15086 2385
rect -15132 2313 -15126 2347
rect -15092 2313 -15086 2347
rect -15132 2275 -15086 2313
rect -15132 2241 -15126 2275
rect -15092 2241 -15086 2275
rect -15132 2203 -15086 2241
rect -15132 2169 -15126 2203
rect -15092 2169 -15086 2203
rect -15132 2131 -15086 2169
rect -15132 2097 -15126 2131
rect -15092 2097 -15086 2131
rect -15132 2059 -15086 2097
rect -15132 2025 -15126 2059
rect -15092 2025 -15086 2059
rect -15132 1987 -15086 2025
rect -15132 1953 -15126 1987
rect -15092 1953 -15086 1987
rect -15132 1915 -15086 1953
rect -15132 1881 -15126 1915
rect -15092 1881 -15086 1915
rect -15132 1866 -15086 1881
rect -15036 2851 -14990 2866
rect -15036 2817 -15030 2851
rect -14996 2817 -14990 2851
rect -15036 2779 -14990 2817
rect -15036 2745 -15030 2779
rect -14996 2745 -14990 2779
rect -15036 2707 -14990 2745
rect -15036 2673 -15030 2707
rect -14996 2673 -14990 2707
rect -15036 2635 -14990 2673
rect -15036 2601 -15030 2635
rect -14996 2601 -14990 2635
rect -15036 2563 -14990 2601
rect -15036 2529 -15030 2563
rect -14996 2529 -14990 2563
rect -15036 2491 -14990 2529
rect -15036 2457 -15030 2491
rect -14996 2457 -14990 2491
rect -15036 2419 -14990 2457
rect -15036 2385 -15030 2419
rect -14996 2385 -14990 2419
rect -15036 2347 -14990 2385
rect -15036 2313 -15030 2347
rect -14996 2313 -14990 2347
rect -15036 2275 -14990 2313
rect -15036 2241 -15030 2275
rect -14996 2241 -14990 2275
rect -15036 2203 -14990 2241
rect -15036 2169 -15030 2203
rect -14996 2169 -14990 2203
rect -15036 2131 -14990 2169
rect -15036 2097 -15030 2131
rect -14996 2097 -14990 2131
rect -15036 2059 -14990 2097
rect -15036 2025 -15030 2059
rect -14996 2025 -14990 2059
rect -15036 1987 -14990 2025
rect -15036 1953 -15030 1987
rect -14996 1953 -14990 1987
rect -15036 1915 -14990 1953
rect -15036 1881 -15030 1915
rect -14996 1881 -14990 1915
rect -15036 1866 -14990 1881
rect -14940 2851 -14894 2866
rect -14940 2817 -14934 2851
rect -14900 2817 -14894 2851
rect -14940 2779 -14894 2817
rect -14940 2745 -14934 2779
rect -14900 2745 -14894 2779
rect -14940 2707 -14894 2745
rect -14940 2673 -14934 2707
rect -14900 2673 -14894 2707
rect -14940 2635 -14894 2673
rect -14940 2601 -14934 2635
rect -14900 2601 -14894 2635
rect -14940 2563 -14894 2601
rect -14940 2529 -14934 2563
rect -14900 2529 -14894 2563
rect -14940 2491 -14894 2529
rect -14940 2457 -14934 2491
rect -14900 2457 -14894 2491
rect -14940 2419 -14894 2457
rect -14940 2385 -14934 2419
rect -14900 2385 -14894 2419
rect -14940 2347 -14894 2385
rect -14940 2313 -14934 2347
rect -14900 2313 -14894 2347
rect -14940 2275 -14894 2313
rect -14940 2241 -14934 2275
rect -14900 2241 -14894 2275
rect -14940 2203 -14894 2241
rect -14940 2169 -14934 2203
rect -14900 2169 -14894 2203
rect -14940 2131 -14894 2169
rect -14940 2097 -14934 2131
rect -14900 2097 -14894 2131
rect -14940 2059 -14894 2097
rect -14940 2025 -14934 2059
rect -14900 2025 -14894 2059
rect -14940 1987 -14894 2025
rect -14940 1953 -14934 1987
rect -14900 1953 -14894 1987
rect -14940 1915 -14894 1953
rect -14940 1881 -14934 1915
rect -14900 1881 -14894 1915
rect -14940 1866 -14894 1881
rect -14844 2851 -14798 2866
rect -14844 2817 -14838 2851
rect -14804 2817 -14798 2851
rect -14844 2779 -14798 2817
rect -14844 2745 -14838 2779
rect -14804 2745 -14798 2779
rect -14844 2707 -14798 2745
rect -14844 2673 -14838 2707
rect -14804 2673 -14798 2707
rect -14844 2635 -14798 2673
rect -14844 2601 -14838 2635
rect -14804 2601 -14798 2635
rect -14844 2563 -14798 2601
rect -14844 2529 -14838 2563
rect -14804 2529 -14798 2563
rect -14844 2491 -14798 2529
rect -14844 2457 -14838 2491
rect -14804 2457 -14798 2491
rect -14844 2419 -14798 2457
rect -14844 2385 -14838 2419
rect -14804 2385 -14798 2419
rect -14844 2347 -14798 2385
rect -14844 2313 -14838 2347
rect -14804 2313 -14798 2347
rect -14844 2275 -14798 2313
rect -14844 2241 -14838 2275
rect -14804 2241 -14798 2275
rect -14844 2203 -14798 2241
rect -14844 2169 -14838 2203
rect -14804 2169 -14798 2203
rect -14844 2131 -14798 2169
rect -14844 2097 -14838 2131
rect -14804 2097 -14798 2131
rect -14844 2059 -14798 2097
rect -14844 2025 -14838 2059
rect -14804 2025 -14798 2059
rect -14844 1987 -14798 2025
rect -14844 1953 -14838 1987
rect -14804 1953 -14798 1987
rect -14844 1915 -14798 1953
rect -14844 1881 -14838 1915
rect -14804 1881 -14798 1915
rect -14844 1866 -14798 1881
rect -14748 2851 -14702 2866
rect -14748 2817 -14742 2851
rect -14708 2817 -14702 2851
rect -14748 2779 -14702 2817
rect -14748 2745 -14742 2779
rect -14708 2745 -14702 2779
rect -14748 2707 -14702 2745
rect -14748 2673 -14742 2707
rect -14708 2673 -14702 2707
rect -14748 2635 -14702 2673
rect -14748 2601 -14742 2635
rect -14708 2601 -14702 2635
rect -14748 2563 -14702 2601
rect -14748 2529 -14742 2563
rect -14708 2529 -14702 2563
rect -14748 2491 -14702 2529
rect -14748 2457 -14742 2491
rect -14708 2457 -14702 2491
rect -14748 2419 -14702 2457
rect -14748 2385 -14742 2419
rect -14708 2385 -14702 2419
rect -14748 2347 -14702 2385
rect -14748 2313 -14742 2347
rect -14708 2313 -14702 2347
rect -14748 2275 -14702 2313
rect -14748 2241 -14742 2275
rect -14708 2241 -14702 2275
rect -14748 2203 -14702 2241
rect -14748 2169 -14742 2203
rect -14708 2169 -14702 2203
rect -14748 2131 -14702 2169
rect -14748 2097 -14742 2131
rect -14708 2097 -14702 2131
rect -14748 2059 -14702 2097
rect -14748 2025 -14742 2059
rect -14708 2025 -14702 2059
rect -14748 1987 -14702 2025
rect -14748 1953 -14742 1987
rect -14708 1953 -14702 1987
rect -14748 1915 -14702 1953
rect -14748 1881 -14742 1915
rect -14708 1881 -14702 1915
rect -14748 1866 -14702 1881
rect -14520 2843 -14474 2858
rect -14520 2809 -14514 2843
rect -14480 2809 -14474 2843
rect -14520 2771 -14474 2809
rect -14520 2737 -14514 2771
rect -14480 2737 -14474 2771
rect -14520 2699 -14474 2737
rect -14520 2665 -14514 2699
rect -14480 2665 -14474 2699
rect -14520 2627 -14474 2665
rect -14520 2593 -14514 2627
rect -14480 2593 -14474 2627
rect -14520 2555 -14474 2593
rect -14520 2521 -14514 2555
rect -14480 2521 -14474 2555
rect -14520 2483 -14474 2521
rect -14520 2449 -14514 2483
rect -14480 2449 -14474 2483
rect -14520 2411 -14474 2449
rect -14520 2377 -14514 2411
rect -14480 2377 -14474 2411
rect -14520 2339 -14474 2377
rect -14520 2305 -14514 2339
rect -14480 2305 -14474 2339
rect -14520 2267 -14474 2305
rect -14520 2233 -14514 2267
rect -14480 2233 -14474 2267
rect -14520 2195 -14474 2233
rect -14520 2161 -14514 2195
rect -14480 2161 -14474 2195
rect -14520 2123 -14474 2161
rect -14520 2089 -14514 2123
rect -14480 2089 -14474 2123
rect -14520 2051 -14474 2089
rect -14520 2017 -14514 2051
rect -14480 2017 -14474 2051
rect -14520 1979 -14474 2017
rect -14520 1945 -14514 1979
rect -14480 1945 -14474 1979
rect -14520 1907 -14474 1945
rect -14520 1873 -14514 1907
rect -14480 1873 -14474 1907
rect -14520 1858 -14474 1873
rect -14424 2843 -14378 2858
rect -14424 2809 -14418 2843
rect -14384 2809 -14378 2843
rect -14424 2771 -14378 2809
rect -14424 2737 -14418 2771
rect -14384 2737 -14378 2771
rect -14424 2699 -14378 2737
rect -14424 2665 -14418 2699
rect -14384 2665 -14378 2699
rect -14424 2627 -14378 2665
rect -14424 2593 -14418 2627
rect -14384 2593 -14378 2627
rect -14424 2555 -14378 2593
rect -14424 2521 -14418 2555
rect -14384 2521 -14378 2555
rect -14424 2483 -14378 2521
rect -14424 2449 -14418 2483
rect -14384 2449 -14378 2483
rect -14424 2411 -14378 2449
rect -14424 2377 -14418 2411
rect -14384 2377 -14378 2411
rect -14424 2339 -14378 2377
rect -14424 2305 -14418 2339
rect -14384 2305 -14378 2339
rect -14424 2267 -14378 2305
rect -14424 2233 -14418 2267
rect -14384 2233 -14378 2267
rect -14424 2195 -14378 2233
rect -14424 2161 -14418 2195
rect -14384 2161 -14378 2195
rect -14424 2123 -14378 2161
rect -14424 2089 -14418 2123
rect -14384 2089 -14378 2123
rect -14424 2051 -14378 2089
rect -14424 2017 -14418 2051
rect -14384 2017 -14378 2051
rect -14424 1979 -14378 2017
rect -14424 1945 -14418 1979
rect -14384 1945 -14378 1979
rect -14424 1907 -14378 1945
rect -14424 1873 -14418 1907
rect -14384 1873 -14378 1907
rect -14424 1858 -14378 1873
rect -14328 2843 -14282 2858
rect -14328 2809 -14322 2843
rect -14288 2809 -14282 2843
rect -14328 2771 -14282 2809
rect -14328 2737 -14322 2771
rect -14288 2737 -14282 2771
rect -14328 2699 -14282 2737
rect -14328 2665 -14322 2699
rect -14288 2665 -14282 2699
rect -14328 2627 -14282 2665
rect -14328 2593 -14322 2627
rect -14288 2593 -14282 2627
rect -14328 2555 -14282 2593
rect -14328 2521 -14322 2555
rect -14288 2521 -14282 2555
rect -14328 2483 -14282 2521
rect -14328 2449 -14322 2483
rect -14288 2449 -14282 2483
rect -14328 2411 -14282 2449
rect -14328 2377 -14322 2411
rect -14288 2377 -14282 2411
rect -14328 2339 -14282 2377
rect -14328 2305 -14322 2339
rect -14288 2305 -14282 2339
rect -14328 2267 -14282 2305
rect -14328 2233 -14322 2267
rect -14288 2233 -14282 2267
rect -14328 2195 -14282 2233
rect -14328 2161 -14322 2195
rect -14288 2161 -14282 2195
rect -14328 2123 -14282 2161
rect -14328 2089 -14322 2123
rect -14288 2089 -14282 2123
rect -14328 2051 -14282 2089
rect -14328 2017 -14322 2051
rect -14288 2017 -14282 2051
rect -14328 1979 -14282 2017
rect -14328 1945 -14322 1979
rect -14288 1945 -14282 1979
rect -14328 1907 -14282 1945
rect -14328 1873 -14322 1907
rect -14288 1873 -14282 1907
rect -14328 1858 -14282 1873
rect -14232 2843 -14186 2858
rect -14232 2809 -14226 2843
rect -14192 2809 -14186 2843
rect -14232 2771 -14186 2809
rect -14232 2737 -14226 2771
rect -14192 2737 -14186 2771
rect -14232 2699 -14186 2737
rect -14232 2665 -14226 2699
rect -14192 2665 -14186 2699
rect -14232 2627 -14186 2665
rect -14232 2593 -14226 2627
rect -14192 2593 -14186 2627
rect -14232 2555 -14186 2593
rect -14232 2521 -14226 2555
rect -14192 2521 -14186 2555
rect -14232 2483 -14186 2521
rect -14232 2449 -14226 2483
rect -14192 2449 -14186 2483
rect -14232 2411 -14186 2449
rect -14232 2377 -14226 2411
rect -14192 2377 -14186 2411
rect -14232 2339 -14186 2377
rect -14232 2305 -14226 2339
rect -14192 2305 -14186 2339
rect -14232 2267 -14186 2305
rect -14232 2233 -14226 2267
rect -14192 2233 -14186 2267
rect -14232 2195 -14186 2233
rect -14232 2161 -14226 2195
rect -14192 2161 -14186 2195
rect -14232 2123 -14186 2161
rect -14232 2089 -14226 2123
rect -14192 2089 -14186 2123
rect -14232 2051 -14186 2089
rect -14232 2017 -14226 2051
rect -14192 2017 -14186 2051
rect -14232 1979 -14186 2017
rect -14232 1945 -14226 1979
rect -14192 1945 -14186 1979
rect -14232 1907 -14186 1945
rect -14232 1873 -14226 1907
rect -14192 1873 -14186 1907
rect -14232 1858 -14186 1873
rect -14136 2843 -14090 2858
rect -14136 2809 -14130 2843
rect -14096 2809 -14090 2843
rect -14136 2771 -14090 2809
rect -14136 2737 -14130 2771
rect -14096 2737 -14090 2771
rect -14136 2699 -14090 2737
rect -14136 2665 -14130 2699
rect -14096 2665 -14090 2699
rect -14136 2627 -14090 2665
rect -14136 2593 -14130 2627
rect -14096 2593 -14090 2627
rect -14136 2555 -14090 2593
rect -14136 2521 -14130 2555
rect -14096 2521 -14090 2555
rect -14136 2483 -14090 2521
rect -14136 2449 -14130 2483
rect -14096 2449 -14090 2483
rect -14136 2411 -14090 2449
rect -14136 2377 -14130 2411
rect -14096 2377 -14090 2411
rect -14136 2339 -14090 2377
rect -14136 2305 -14130 2339
rect -14096 2305 -14090 2339
rect -14136 2267 -14090 2305
rect -14136 2233 -14130 2267
rect -14096 2233 -14090 2267
rect -14136 2195 -14090 2233
rect -14136 2161 -14130 2195
rect -14096 2161 -14090 2195
rect -14136 2123 -14090 2161
rect -14136 2089 -14130 2123
rect -14096 2089 -14090 2123
rect -14136 2051 -14090 2089
rect -14136 2017 -14130 2051
rect -14096 2017 -14090 2051
rect -14136 1979 -14090 2017
rect -14136 1945 -14130 1979
rect -14096 1945 -14090 1979
rect -14136 1907 -14090 1945
rect -14136 1873 -14130 1907
rect -14096 1873 -14090 1907
rect -14136 1858 -14090 1873
rect -14040 2843 -13994 2858
rect -14040 2809 -14034 2843
rect -14000 2809 -13994 2843
rect -14040 2771 -13994 2809
rect -14040 2737 -14034 2771
rect -14000 2737 -13994 2771
rect -14040 2699 -13994 2737
rect -14040 2665 -14034 2699
rect -14000 2665 -13994 2699
rect -14040 2627 -13994 2665
rect -14040 2593 -14034 2627
rect -14000 2593 -13994 2627
rect -14040 2555 -13994 2593
rect -14040 2521 -14034 2555
rect -14000 2521 -13994 2555
rect -14040 2483 -13994 2521
rect -14040 2449 -14034 2483
rect -14000 2449 -13994 2483
rect -14040 2411 -13994 2449
rect -14040 2377 -14034 2411
rect -14000 2377 -13994 2411
rect -14040 2339 -13994 2377
rect -14040 2305 -14034 2339
rect -14000 2305 -13994 2339
rect -14040 2267 -13994 2305
rect -14040 2233 -14034 2267
rect -14000 2233 -13994 2267
rect -14040 2195 -13994 2233
rect -14040 2161 -14034 2195
rect -14000 2161 -13994 2195
rect -14040 2123 -13994 2161
rect -14040 2089 -14034 2123
rect -14000 2089 -13994 2123
rect -14040 2051 -13994 2089
rect -14040 2017 -14034 2051
rect -14000 2017 -13994 2051
rect -14040 1979 -13994 2017
rect -14040 1945 -14034 1979
rect -14000 1945 -13994 1979
rect -14040 1907 -13994 1945
rect -14040 1873 -14034 1907
rect -14000 1873 -13994 1907
rect -14040 1858 -13994 1873
rect -13944 2843 -13898 2858
rect -13944 2809 -13938 2843
rect -13904 2809 -13898 2843
rect -13944 2771 -13898 2809
rect -13944 2737 -13938 2771
rect -13904 2737 -13898 2771
rect -13944 2699 -13898 2737
rect -13944 2665 -13938 2699
rect -13904 2665 -13898 2699
rect -13944 2627 -13898 2665
rect -13944 2593 -13938 2627
rect -13904 2593 -13898 2627
rect -13944 2555 -13898 2593
rect -13944 2521 -13938 2555
rect -13904 2521 -13898 2555
rect -13944 2483 -13898 2521
rect -13944 2449 -13938 2483
rect -13904 2449 -13898 2483
rect -13944 2411 -13898 2449
rect -13944 2377 -13938 2411
rect -13904 2377 -13898 2411
rect -13944 2339 -13898 2377
rect -13944 2305 -13938 2339
rect -13904 2305 -13898 2339
rect -13944 2267 -13898 2305
rect -13944 2233 -13938 2267
rect -13904 2233 -13898 2267
rect -13944 2195 -13898 2233
rect -13944 2161 -13938 2195
rect -13904 2161 -13898 2195
rect -13944 2123 -13898 2161
rect -13944 2089 -13938 2123
rect -13904 2089 -13898 2123
rect -13944 2051 -13898 2089
rect -13944 2017 -13938 2051
rect -13904 2017 -13898 2051
rect -13944 1979 -13898 2017
rect -13944 1945 -13938 1979
rect -13904 1945 -13898 1979
rect -13944 1907 -13898 1945
rect -13944 1873 -13938 1907
rect -13904 1873 -13898 1907
rect -13944 1858 -13898 1873
rect -13848 2843 -13802 2858
rect -13848 2809 -13842 2843
rect -13808 2809 -13802 2843
rect -13848 2771 -13802 2809
rect -13848 2737 -13842 2771
rect -13808 2737 -13802 2771
rect -13848 2699 -13802 2737
rect -13848 2665 -13842 2699
rect -13808 2665 -13802 2699
rect -13848 2627 -13802 2665
rect -13848 2593 -13842 2627
rect -13808 2593 -13802 2627
rect -13848 2555 -13802 2593
rect -13848 2521 -13842 2555
rect -13808 2521 -13802 2555
rect -13848 2483 -13802 2521
rect -13848 2449 -13842 2483
rect -13808 2449 -13802 2483
rect -13848 2411 -13802 2449
rect -13848 2377 -13842 2411
rect -13808 2377 -13802 2411
rect -13848 2339 -13802 2377
rect -13848 2305 -13842 2339
rect -13808 2305 -13802 2339
rect -13848 2267 -13802 2305
rect -13848 2233 -13842 2267
rect -13808 2233 -13802 2267
rect -13848 2195 -13802 2233
rect -13848 2161 -13842 2195
rect -13808 2161 -13802 2195
rect -13848 2123 -13802 2161
rect -13848 2089 -13842 2123
rect -13808 2089 -13802 2123
rect -13848 2051 -13802 2089
rect -13848 2017 -13842 2051
rect -13808 2017 -13802 2051
rect -13848 1979 -13802 2017
rect -13848 1945 -13842 1979
rect -13808 1945 -13802 1979
rect -13848 1907 -13802 1945
rect -13848 1873 -13842 1907
rect -13808 1873 -13802 1907
rect -13848 1858 -13802 1873
rect -13752 2843 -13706 2858
rect -13752 2809 -13746 2843
rect -13712 2809 -13706 2843
rect -13752 2771 -13706 2809
rect -13752 2737 -13746 2771
rect -13712 2737 -13706 2771
rect -13752 2699 -13706 2737
rect -13752 2665 -13746 2699
rect -13712 2665 -13706 2699
rect -13752 2627 -13706 2665
rect -13752 2593 -13746 2627
rect -13712 2593 -13706 2627
rect -13752 2555 -13706 2593
rect -13752 2521 -13746 2555
rect -13712 2521 -13706 2555
rect -13752 2483 -13706 2521
rect -13752 2449 -13746 2483
rect -13712 2449 -13706 2483
rect -13752 2411 -13706 2449
rect -13752 2377 -13746 2411
rect -13712 2377 -13706 2411
rect -13752 2339 -13706 2377
rect -13752 2305 -13746 2339
rect -13712 2305 -13706 2339
rect -13752 2267 -13706 2305
rect -13752 2233 -13746 2267
rect -13712 2233 -13706 2267
rect -13752 2195 -13706 2233
rect -13752 2161 -13746 2195
rect -13712 2161 -13706 2195
rect -13752 2123 -13706 2161
rect -13752 2089 -13746 2123
rect -13712 2089 -13706 2123
rect -13752 2051 -13706 2089
rect -13752 2017 -13746 2051
rect -13712 2017 -13706 2051
rect -13752 1979 -13706 2017
rect -13752 1945 -13746 1979
rect -13712 1945 -13706 1979
rect -13752 1907 -13706 1945
rect -13752 1873 -13746 1907
rect -13712 1873 -13706 1907
rect -13752 1858 -13706 1873
rect -13656 2843 -13610 2858
rect -13656 2809 -13650 2843
rect -13616 2809 -13610 2843
rect -13656 2771 -13610 2809
rect -13656 2737 -13650 2771
rect -13616 2737 -13610 2771
rect -13656 2699 -13610 2737
rect -13656 2665 -13650 2699
rect -13616 2665 -13610 2699
rect -13656 2627 -13610 2665
rect -13656 2593 -13650 2627
rect -13616 2593 -13610 2627
rect -13656 2555 -13610 2593
rect -13656 2521 -13650 2555
rect -13616 2521 -13610 2555
rect -13656 2483 -13610 2521
rect -13656 2449 -13650 2483
rect -13616 2449 -13610 2483
rect -13656 2411 -13610 2449
rect -13656 2377 -13650 2411
rect -13616 2377 -13610 2411
rect -13656 2339 -13610 2377
rect -13656 2305 -13650 2339
rect -13616 2305 -13610 2339
rect -13656 2267 -13610 2305
rect -13656 2233 -13650 2267
rect -13616 2233 -13610 2267
rect -13656 2195 -13610 2233
rect -13656 2161 -13650 2195
rect -13616 2161 -13610 2195
rect -13656 2123 -13610 2161
rect -13656 2089 -13650 2123
rect -13616 2089 -13610 2123
rect -13656 2051 -13610 2089
rect -13656 2017 -13650 2051
rect -13616 2017 -13610 2051
rect -13656 1979 -13610 2017
rect -13656 1945 -13650 1979
rect -13616 1945 -13610 1979
rect -13656 1907 -13610 1945
rect -13656 1873 -13650 1907
rect -13616 1873 -13610 1907
rect -13656 1858 -13610 1873
rect -13560 2843 -13514 2858
rect -13560 2809 -13554 2843
rect -13520 2809 -13514 2843
rect -13560 2771 -13514 2809
rect -13560 2737 -13554 2771
rect -13520 2737 -13514 2771
rect -13560 2699 -13514 2737
rect -13560 2665 -13554 2699
rect -13520 2665 -13514 2699
rect -13560 2627 -13514 2665
rect -13560 2593 -13554 2627
rect -13520 2593 -13514 2627
rect -13560 2555 -13514 2593
rect -13560 2521 -13554 2555
rect -13520 2521 -13514 2555
rect -13560 2483 -13514 2521
rect -13560 2449 -13554 2483
rect -13520 2449 -13514 2483
rect -13560 2411 -13514 2449
rect -13560 2377 -13554 2411
rect -13520 2377 -13514 2411
rect -13560 2339 -13514 2377
rect -13560 2305 -13554 2339
rect -13520 2305 -13514 2339
rect -13560 2267 -13514 2305
rect -13560 2233 -13554 2267
rect -13520 2233 -13514 2267
rect -13560 2195 -13514 2233
rect -13560 2161 -13554 2195
rect -13520 2161 -13514 2195
rect -13560 2123 -13514 2161
rect -13560 2089 -13554 2123
rect -13520 2089 -13514 2123
rect -13560 2051 -13514 2089
rect -13560 2017 -13554 2051
rect -13520 2017 -13514 2051
rect -13560 1979 -13514 2017
rect -13560 1945 -13554 1979
rect -13520 1945 -13514 1979
rect -13560 1907 -13514 1945
rect -13560 1873 -13554 1907
rect -13520 1873 -13514 1907
rect -13560 1858 -13514 1873
rect -13464 2843 -13418 2858
rect -13464 2809 -13458 2843
rect -13424 2809 -13418 2843
rect -13464 2771 -13418 2809
rect -13464 2737 -13458 2771
rect -13424 2737 -13418 2771
rect -13464 2699 -13418 2737
rect -13464 2665 -13458 2699
rect -13424 2665 -13418 2699
rect -13464 2627 -13418 2665
rect -13464 2593 -13458 2627
rect -13424 2593 -13418 2627
rect -13464 2555 -13418 2593
rect -13464 2521 -13458 2555
rect -13424 2521 -13418 2555
rect -13464 2483 -13418 2521
rect -13464 2449 -13458 2483
rect -13424 2449 -13418 2483
rect -13464 2411 -13418 2449
rect -13464 2377 -13458 2411
rect -13424 2377 -13418 2411
rect -13464 2339 -13418 2377
rect -13464 2305 -13458 2339
rect -13424 2305 -13418 2339
rect -13464 2267 -13418 2305
rect -13464 2233 -13458 2267
rect -13424 2233 -13418 2267
rect -13464 2195 -13418 2233
rect -13464 2161 -13458 2195
rect -13424 2161 -13418 2195
rect -13464 2123 -13418 2161
rect -13464 2089 -13458 2123
rect -13424 2089 -13418 2123
rect -13464 2051 -13418 2089
rect -13464 2017 -13458 2051
rect -13424 2017 -13418 2051
rect -13464 1979 -13418 2017
rect -13464 1945 -13458 1979
rect -13424 1945 -13418 1979
rect -13464 1907 -13418 1945
rect -13464 1873 -13458 1907
rect -13424 1873 -13418 1907
rect -13464 1858 -13418 1873
rect -13368 2843 -13322 2858
rect -13368 2809 -13362 2843
rect -13328 2809 -13322 2843
rect -13368 2771 -13322 2809
rect -13368 2737 -13362 2771
rect -13328 2737 -13322 2771
rect -13368 2699 -13322 2737
rect -13368 2665 -13362 2699
rect -13328 2665 -13322 2699
rect -13368 2627 -13322 2665
rect -13368 2593 -13362 2627
rect -13328 2593 -13322 2627
rect -13368 2555 -13322 2593
rect -13368 2521 -13362 2555
rect -13328 2521 -13322 2555
rect -13368 2483 -13322 2521
rect -13368 2449 -13362 2483
rect -13328 2449 -13322 2483
rect -13368 2411 -13322 2449
rect -13368 2377 -13362 2411
rect -13328 2377 -13322 2411
rect -13368 2339 -13322 2377
rect -13368 2305 -13362 2339
rect -13328 2305 -13322 2339
rect -13368 2267 -13322 2305
rect -13368 2233 -13362 2267
rect -13328 2233 -13322 2267
rect -13368 2195 -13322 2233
rect -13368 2161 -13362 2195
rect -13328 2161 -13322 2195
rect -13368 2123 -13322 2161
rect -13368 2089 -13362 2123
rect -13328 2089 -13322 2123
rect -13368 2051 -13322 2089
rect -13368 2017 -13362 2051
rect -13328 2017 -13322 2051
rect -13368 1979 -13322 2017
rect -13368 1945 -13362 1979
rect -13328 1945 -13322 1979
rect -13368 1907 -13322 1945
rect -13368 1873 -13362 1907
rect -13328 1873 -13322 1907
rect -13368 1858 -13322 1873
rect -13272 2843 -13226 2858
rect -13272 2809 -13266 2843
rect -13232 2809 -13226 2843
rect -13272 2771 -13226 2809
rect -13272 2737 -13266 2771
rect -13232 2737 -13226 2771
rect -13272 2699 -13226 2737
rect -13272 2665 -13266 2699
rect -13232 2665 -13226 2699
rect -13272 2627 -13226 2665
rect -13272 2593 -13266 2627
rect -13232 2593 -13226 2627
rect -13272 2555 -13226 2593
rect -13272 2521 -13266 2555
rect -13232 2521 -13226 2555
rect -13272 2483 -13226 2521
rect -13272 2449 -13266 2483
rect -13232 2449 -13226 2483
rect -13272 2411 -13226 2449
rect -13272 2377 -13266 2411
rect -13232 2377 -13226 2411
rect -13272 2339 -13226 2377
rect -13272 2305 -13266 2339
rect -13232 2305 -13226 2339
rect -13272 2267 -13226 2305
rect -13272 2233 -13266 2267
rect -13232 2233 -13226 2267
rect -13272 2195 -13226 2233
rect -13272 2161 -13266 2195
rect -13232 2161 -13226 2195
rect -13272 2123 -13226 2161
rect -13272 2089 -13266 2123
rect -13232 2089 -13226 2123
rect -13272 2051 -13226 2089
rect -13272 2017 -13266 2051
rect -13232 2017 -13226 2051
rect -13272 1979 -13226 2017
rect -13272 1945 -13266 1979
rect -13232 1945 -13226 1979
rect -13272 1907 -13226 1945
rect -13272 1873 -13266 1907
rect -13232 1873 -13226 1907
rect -13272 1858 -13226 1873
rect -13176 2843 -13130 2858
rect -13176 2809 -13170 2843
rect -13136 2809 -13130 2843
rect -13176 2771 -13130 2809
rect -13176 2737 -13170 2771
rect -13136 2737 -13130 2771
rect -13176 2699 -13130 2737
rect -13176 2665 -13170 2699
rect -13136 2665 -13130 2699
rect -13176 2627 -13130 2665
rect -13176 2593 -13170 2627
rect -13136 2593 -13130 2627
rect -13176 2555 -13130 2593
rect -13176 2521 -13170 2555
rect -13136 2521 -13130 2555
rect -13176 2483 -13130 2521
rect -13176 2449 -13170 2483
rect -13136 2449 -13130 2483
rect -13176 2411 -13130 2449
rect -13176 2377 -13170 2411
rect -13136 2377 -13130 2411
rect -13176 2339 -13130 2377
rect -13176 2305 -13170 2339
rect -13136 2305 -13130 2339
rect -13176 2267 -13130 2305
rect -13176 2233 -13170 2267
rect -13136 2233 -13130 2267
rect -13176 2195 -13130 2233
rect -13176 2161 -13170 2195
rect -13136 2161 -13130 2195
rect -13176 2123 -13130 2161
rect -13176 2089 -13170 2123
rect -13136 2089 -13130 2123
rect -13176 2051 -13130 2089
rect -13176 2017 -13170 2051
rect -13136 2017 -13130 2051
rect -13176 1979 -13130 2017
rect -13176 1945 -13170 1979
rect -13136 1945 -13130 1979
rect -13176 1907 -13130 1945
rect -13176 1873 -13170 1907
rect -13136 1873 -13130 1907
rect -13176 1858 -13130 1873
rect -13080 2843 -13034 2858
rect -13080 2809 -13074 2843
rect -13040 2809 -13034 2843
rect -13080 2771 -13034 2809
rect -13080 2737 -13074 2771
rect -13040 2737 -13034 2771
rect -13080 2699 -13034 2737
rect -13080 2665 -13074 2699
rect -13040 2665 -13034 2699
rect -13080 2627 -13034 2665
rect -13080 2593 -13074 2627
rect -13040 2593 -13034 2627
rect -13080 2555 -13034 2593
rect -13080 2521 -13074 2555
rect -13040 2521 -13034 2555
rect -13080 2483 -13034 2521
rect -13080 2449 -13074 2483
rect -13040 2449 -13034 2483
rect -13080 2411 -13034 2449
rect -13080 2377 -13074 2411
rect -13040 2377 -13034 2411
rect -13080 2339 -13034 2377
rect -13080 2305 -13074 2339
rect -13040 2305 -13034 2339
rect -13080 2267 -13034 2305
rect -13080 2233 -13074 2267
rect -13040 2233 -13034 2267
rect -13080 2195 -13034 2233
rect -13080 2161 -13074 2195
rect -13040 2161 -13034 2195
rect -13080 2123 -13034 2161
rect -13080 2089 -13074 2123
rect -13040 2089 -13034 2123
rect -13080 2051 -13034 2089
rect -13080 2017 -13074 2051
rect -13040 2017 -13034 2051
rect -13080 1979 -13034 2017
rect -13080 1945 -13074 1979
rect -13040 1945 -13034 1979
rect -13080 1907 -13034 1945
rect -13080 1873 -13074 1907
rect -13040 1873 -13034 1907
rect -13080 1858 -13034 1873
rect -12842 2847 -12796 2862
rect -12842 2813 -12836 2847
rect -12802 2813 -12796 2847
rect -12842 2775 -12796 2813
rect -12842 2741 -12836 2775
rect -12802 2741 -12796 2775
rect -12842 2703 -12796 2741
rect -12842 2669 -12836 2703
rect -12802 2669 -12796 2703
rect -12842 2631 -12796 2669
rect -12842 2597 -12836 2631
rect -12802 2597 -12796 2631
rect -12842 2559 -12796 2597
rect -12842 2525 -12836 2559
rect -12802 2525 -12796 2559
rect -12842 2487 -12796 2525
rect -12842 2453 -12836 2487
rect -12802 2453 -12796 2487
rect -12842 2415 -12796 2453
rect -12842 2381 -12836 2415
rect -12802 2381 -12796 2415
rect -12842 2343 -12796 2381
rect -12842 2309 -12836 2343
rect -12802 2309 -12796 2343
rect -12842 2271 -12796 2309
rect -12842 2237 -12836 2271
rect -12802 2237 -12796 2271
rect -12842 2199 -12796 2237
rect -12842 2165 -12836 2199
rect -12802 2165 -12796 2199
rect -12842 2127 -12796 2165
rect -12842 2093 -12836 2127
rect -12802 2093 -12796 2127
rect -12842 2055 -12796 2093
rect -12842 2021 -12836 2055
rect -12802 2021 -12796 2055
rect -12842 1983 -12796 2021
rect -12842 1949 -12836 1983
rect -12802 1949 -12796 1983
rect -12842 1911 -12796 1949
rect -12842 1877 -12836 1911
rect -12802 1877 -12796 1911
rect -12842 1862 -12796 1877
rect -12746 2847 -12700 2862
rect -12746 2813 -12740 2847
rect -12706 2813 -12700 2847
rect -12746 2775 -12700 2813
rect -12746 2741 -12740 2775
rect -12706 2741 -12700 2775
rect -12746 2703 -12700 2741
rect -12746 2669 -12740 2703
rect -12706 2669 -12700 2703
rect -12746 2631 -12700 2669
rect -12746 2597 -12740 2631
rect -12706 2597 -12700 2631
rect -12746 2559 -12700 2597
rect -12746 2525 -12740 2559
rect -12706 2525 -12700 2559
rect -12746 2487 -12700 2525
rect -12746 2453 -12740 2487
rect -12706 2453 -12700 2487
rect -12746 2415 -12700 2453
rect -12746 2381 -12740 2415
rect -12706 2381 -12700 2415
rect -12746 2343 -12700 2381
rect -12746 2309 -12740 2343
rect -12706 2309 -12700 2343
rect -12746 2271 -12700 2309
rect -12746 2237 -12740 2271
rect -12706 2237 -12700 2271
rect -12746 2199 -12700 2237
rect -12746 2165 -12740 2199
rect -12706 2165 -12700 2199
rect -12746 2127 -12700 2165
rect -12746 2093 -12740 2127
rect -12706 2093 -12700 2127
rect -12746 2055 -12700 2093
rect -12746 2021 -12740 2055
rect -12706 2021 -12700 2055
rect -12746 1983 -12700 2021
rect -12746 1949 -12740 1983
rect -12706 1949 -12700 1983
rect -12746 1911 -12700 1949
rect -12746 1877 -12740 1911
rect -12706 1877 -12700 1911
rect -12746 1862 -12700 1877
rect -12650 2847 -12604 2862
rect -12650 2813 -12644 2847
rect -12610 2813 -12604 2847
rect -12650 2775 -12604 2813
rect -12650 2741 -12644 2775
rect -12610 2741 -12604 2775
rect -12650 2703 -12604 2741
rect -12650 2669 -12644 2703
rect -12610 2669 -12604 2703
rect -12650 2631 -12604 2669
rect -12650 2597 -12644 2631
rect -12610 2597 -12604 2631
rect -12650 2559 -12604 2597
rect -12650 2525 -12644 2559
rect -12610 2525 -12604 2559
rect -12650 2487 -12604 2525
rect -12650 2453 -12644 2487
rect -12610 2453 -12604 2487
rect -12650 2415 -12604 2453
rect -12650 2381 -12644 2415
rect -12610 2381 -12604 2415
rect -12650 2343 -12604 2381
rect -12650 2309 -12644 2343
rect -12610 2309 -12604 2343
rect -12650 2271 -12604 2309
rect -12650 2237 -12644 2271
rect -12610 2237 -12604 2271
rect -12650 2199 -12604 2237
rect -12650 2165 -12644 2199
rect -12610 2165 -12604 2199
rect -12650 2127 -12604 2165
rect -12650 2093 -12644 2127
rect -12610 2093 -12604 2127
rect -12650 2055 -12604 2093
rect -12650 2021 -12644 2055
rect -12610 2021 -12604 2055
rect -12650 1983 -12604 2021
rect -12650 1949 -12644 1983
rect -12610 1949 -12604 1983
rect -12650 1911 -12604 1949
rect -12650 1877 -12644 1911
rect -12610 1877 -12604 1911
rect -12650 1862 -12604 1877
rect -12554 2847 -12508 2862
rect -12554 2813 -12548 2847
rect -12514 2813 -12508 2847
rect -12554 2775 -12508 2813
rect -12554 2741 -12548 2775
rect -12514 2741 -12508 2775
rect -12554 2703 -12508 2741
rect -12554 2669 -12548 2703
rect -12514 2669 -12508 2703
rect -12554 2631 -12508 2669
rect -12554 2597 -12548 2631
rect -12514 2597 -12508 2631
rect -12554 2559 -12508 2597
rect -12554 2525 -12548 2559
rect -12514 2525 -12508 2559
rect -12554 2487 -12508 2525
rect -12554 2453 -12548 2487
rect -12514 2453 -12508 2487
rect -12554 2415 -12508 2453
rect -12554 2381 -12548 2415
rect -12514 2381 -12508 2415
rect -12554 2343 -12508 2381
rect -12554 2309 -12548 2343
rect -12514 2309 -12508 2343
rect -12554 2271 -12508 2309
rect -12554 2237 -12548 2271
rect -12514 2237 -12508 2271
rect -12554 2199 -12508 2237
rect -12554 2165 -12548 2199
rect -12514 2165 -12508 2199
rect -12554 2127 -12508 2165
rect -12554 2093 -12548 2127
rect -12514 2093 -12508 2127
rect -12554 2055 -12508 2093
rect -12554 2021 -12548 2055
rect -12514 2021 -12508 2055
rect -12554 1983 -12508 2021
rect -12554 1949 -12548 1983
rect -12514 1949 -12508 1983
rect -12554 1911 -12508 1949
rect -12554 1877 -12548 1911
rect -12514 1877 -12508 1911
rect -12554 1862 -12508 1877
rect -12458 2847 -12412 2862
rect -12458 2813 -12452 2847
rect -12418 2813 -12412 2847
rect -12458 2775 -12412 2813
rect -12458 2741 -12452 2775
rect -12418 2741 -12412 2775
rect -12458 2703 -12412 2741
rect -12458 2669 -12452 2703
rect -12418 2669 -12412 2703
rect -12458 2631 -12412 2669
rect -12458 2597 -12452 2631
rect -12418 2597 -12412 2631
rect -12458 2559 -12412 2597
rect -12458 2525 -12452 2559
rect -12418 2525 -12412 2559
rect -12458 2487 -12412 2525
rect -12458 2453 -12452 2487
rect -12418 2453 -12412 2487
rect -12458 2415 -12412 2453
rect -12458 2381 -12452 2415
rect -12418 2381 -12412 2415
rect -12458 2343 -12412 2381
rect -12458 2309 -12452 2343
rect -12418 2309 -12412 2343
rect -12458 2271 -12412 2309
rect -12458 2237 -12452 2271
rect -12418 2237 -12412 2271
rect -12458 2199 -12412 2237
rect -12458 2165 -12452 2199
rect -12418 2165 -12412 2199
rect -12458 2127 -12412 2165
rect -12458 2093 -12452 2127
rect -12418 2093 -12412 2127
rect -12458 2055 -12412 2093
rect -12458 2021 -12452 2055
rect -12418 2021 -12412 2055
rect -12458 1983 -12412 2021
rect -12458 1949 -12452 1983
rect -12418 1949 -12412 1983
rect -12458 1911 -12412 1949
rect -12458 1877 -12452 1911
rect -12418 1877 -12412 1911
rect -12458 1862 -12412 1877
rect -12362 2847 -12316 2862
rect -12362 2813 -12356 2847
rect -12322 2813 -12316 2847
rect -12362 2775 -12316 2813
rect -12362 2741 -12356 2775
rect -12322 2741 -12316 2775
rect -12362 2703 -12316 2741
rect -12362 2669 -12356 2703
rect -12322 2669 -12316 2703
rect -12362 2631 -12316 2669
rect -12362 2597 -12356 2631
rect -12322 2597 -12316 2631
rect -12362 2559 -12316 2597
rect -12362 2525 -12356 2559
rect -12322 2525 -12316 2559
rect -12362 2487 -12316 2525
rect -12362 2453 -12356 2487
rect -12322 2453 -12316 2487
rect -12362 2415 -12316 2453
rect -12362 2381 -12356 2415
rect -12322 2381 -12316 2415
rect -12362 2343 -12316 2381
rect -12362 2309 -12356 2343
rect -12322 2309 -12316 2343
rect -12362 2271 -12316 2309
rect -12362 2237 -12356 2271
rect -12322 2237 -12316 2271
rect -12362 2199 -12316 2237
rect -12362 2165 -12356 2199
rect -12322 2165 -12316 2199
rect -12362 2127 -12316 2165
rect -12362 2093 -12356 2127
rect -12322 2093 -12316 2127
rect -12362 2055 -12316 2093
rect -12362 2021 -12356 2055
rect -12322 2021 -12316 2055
rect -12362 1983 -12316 2021
rect -12362 1949 -12356 1983
rect -12322 1949 -12316 1983
rect -12362 1911 -12316 1949
rect -12362 1877 -12356 1911
rect -12322 1877 -12316 1911
rect -12362 1862 -12316 1877
rect -12266 2847 -12220 2862
rect -12266 2813 -12260 2847
rect -12226 2813 -12220 2847
rect -12266 2775 -12220 2813
rect -12266 2741 -12260 2775
rect -12226 2741 -12220 2775
rect -12266 2703 -12220 2741
rect -12266 2669 -12260 2703
rect -12226 2669 -12220 2703
rect -12266 2631 -12220 2669
rect -12266 2597 -12260 2631
rect -12226 2597 -12220 2631
rect -12266 2559 -12220 2597
rect -12266 2525 -12260 2559
rect -12226 2525 -12220 2559
rect -12266 2487 -12220 2525
rect -12266 2453 -12260 2487
rect -12226 2453 -12220 2487
rect -12266 2415 -12220 2453
rect -12266 2381 -12260 2415
rect -12226 2381 -12220 2415
rect -12266 2343 -12220 2381
rect -12266 2309 -12260 2343
rect -12226 2309 -12220 2343
rect -12266 2271 -12220 2309
rect -12266 2237 -12260 2271
rect -12226 2237 -12220 2271
rect -12266 2199 -12220 2237
rect -12266 2165 -12260 2199
rect -12226 2165 -12220 2199
rect -12266 2127 -12220 2165
rect -12266 2093 -12260 2127
rect -12226 2093 -12220 2127
rect -12266 2055 -12220 2093
rect -12266 2021 -12260 2055
rect -12226 2021 -12220 2055
rect -12266 1983 -12220 2021
rect -12266 1949 -12260 1983
rect -12226 1949 -12220 1983
rect -12266 1911 -12220 1949
rect -12266 1877 -12260 1911
rect -12226 1877 -12220 1911
rect -12266 1862 -12220 1877
rect -12170 2847 -12124 2862
rect -12170 2813 -12164 2847
rect -12130 2813 -12124 2847
rect -12170 2775 -12124 2813
rect -12170 2741 -12164 2775
rect -12130 2741 -12124 2775
rect -12170 2703 -12124 2741
rect -12170 2669 -12164 2703
rect -12130 2669 -12124 2703
rect -12170 2631 -12124 2669
rect -12170 2597 -12164 2631
rect -12130 2597 -12124 2631
rect -12170 2559 -12124 2597
rect -12170 2525 -12164 2559
rect -12130 2525 -12124 2559
rect -12170 2487 -12124 2525
rect -12170 2453 -12164 2487
rect -12130 2453 -12124 2487
rect -12170 2415 -12124 2453
rect -12170 2381 -12164 2415
rect -12130 2381 -12124 2415
rect -12170 2343 -12124 2381
rect -12170 2309 -12164 2343
rect -12130 2309 -12124 2343
rect -12170 2271 -12124 2309
rect -12170 2237 -12164 2271
rect -12130 2237 -12124 2271
rect -12170 2199 -12124 2237
rect -12170 2165 -12164 2199
rect -12130 2165 -12124 2199
rect -12170 2127 -12124 2165
rect -12170 2093 -12164 2127
rect -12130 2093 -12124 2127
rect -12170 2055 -12124 2093
rect -12170 2021 -12164 2055
rect -12130 2021 -12124 2055
rect -12170 1983 -12124 2021
rect -12170 1949 -12164 1983
rect -12130 1949 -12124 1983
rect -12170 1911 -12124 1949
rect -12170 1877 -12164 1911
rect -12130 1877 -12124 1911
rect -12170 1862 -12124 1877
rect -12074 2847 -12028 2862
rect -12074 2813 -12068 2847
rect -12034 2813 -12028 2847
rect -12074 2775 -12028 2813
rect -12074 2741 -12068 2775
rect -12034 2741 -12028 2775
rect -12074 2703 -12028 2741
rect -12074 2669 -12068 2703
rect -12034 2669 -12028 2703
rect -12074 2631 -12028 2669
rect -12074 2597 -12068 2631
rect -12034 2597 -12028 2631
rect -12074 2559 -12028 2597
rect -12074 2525 -12068 2559
rect -12034 2525 -12028 2559
rect -12074 2487 -12028 2525
rect -12074 2453 -12068 2487
rect -12034 2453 -12028 2487
rect -12074 2415 -12028 2453
rect -12074 2381 -12068 2415
rect -12034 2381 -12028 2415
rect -12074 2343 -12028 2381
rect -12074 2309 -12068 2343
rect -12034 2309 -12028 2343
rect -12074 2271 -12028 2309
rect -12074 2237 -12068 2271
rect -12034 2237 -12028 2271
rect -12074 2199 -12028 2237
rect -12074 2165 -12068 2199
rect -12034 2165 -12028 2199
rect -12074 2127 -12028 2165
rect -12074 2093 -12068 2127
rect -12034 2093 -12028 2127
rect -12074 2055 -12028 2093
rect -12074 2021 -12068 2055
rect -12034 2021 -12028 2055
rect -12074 1983 -12028 2021
rect -12074 1949 -12068 1983
rect -12034 1949 -12028 1983
rect -12074 1911 -12028 1949
rect -12074 1877 -12068 1911
rect -12034 1877 -12028 1911
rect -12074 1862 -12028 1877
rect -11978 2847 -11932 2862
rect -11978 2813 -11972 2847
rect -11938 2813 -11932 2847
rect -11978 2775 -11932 2813
rect -11978 2741 -11972 2775
rect -11938 2741 -11932 2775
rect -11978 2703 -11932 2741
rect -11978 2669 -11972 2703
rect -11938 2669 -11932 2703
rect -11978 2631 -11932 2669
rect -11978 2597 -11972 2631
rect -11938 2597 -11932 2631
rect -11978 2559 -11932 2597
rect -11978 2525 -11972 2559
rect -11938 2525 -11932 2559
rect -11978 2487 -11932 2525
rect -11978 2453 -11972 2487
rect -11938 2453 -11932 2487
rect -11978 2415 -11932 2453
rect -11978 2381 -11972 2415
rect -11938 2381 -11932 2415
rect -11978 2343 -11932 2381
rect -11978 2309 -11972 2343
rect -11938 2309 -11932 2343
rect -11978 2271 -11932 2309
rect -11978 2237 -11972 2271
rect -11938 2237 -11932 2271
rect -11978 2199 -11932 2237
rect -11978 2165 -11972 2199
rect -11938 2165 -11932 2199
rect -11978 2127 -11932 2165
rect -11978 2093 -11972 2127
rect -11938 2093 -11932 2127
rect -11978 2055 -11932 2093
rect -11978 2021 -11972 2055
rect -11938 2021 -11932 2055
rect -11978 1983 -11932 2021
rect -11978 1949 -11972 1983
rect -11938 1949 -11932 1983
rect -11978 1911 -11932 1949
rect -11978 1877 -11972 1911
rect -11938 1877 -11932 1911
rect -11978 1862 -11932 1877
rect -11882 2847 -11836 2862
rect -11882 2813 -11876 2847
rect -11842 2813 -11836 2847
rect -11882 2775 -11836 2813
rect -11882 2741 -11876 2775
rect -11842 2741 -11836 2775
rect -11882 2703 -11836 2741
rect -11882 2669 -11876 2703
rect -11842 2669 -11836 2703
rect -11882 2631 -11836 2669
rect -11882 2597 -11876 2631
rect -11842 2597 -11836 2631
rect -11882 2559 -11836 2597
rect -11882 2525 -11876 2559
rect -11842 2525 -11836 2559
rect -11882 2487 -11836 2525
rect -11882 2453 -11876 2487
rect -11842 2453 -11836 2487
rect -11882 2415 -11836 2453
rect -11882 2381 -11876 2415
rect -11842 2381 -11836 2415
rect -11882 2343 -11836 2381
rect -11882 2309 -11876 2343
rect -11842 2309 -11836 2343
rect -11882 2271 -11836 2309
rect -11882 2237 -11876 2271
rect -11842 2237 -11836 2271
rect -11882 2199 -11836 2237
rect -11882 2165 -11876 2199
rect -11842 2165 -11836 2199
rect -11882 2127 -11836 2165
rect -11882 2093 -11876 2127
rect -11842 2093 -11836 2127
rect -11882 2055 -11836 2093
rect -11882 2021 -11876 2055
rect -11842 2021 -11836 2055
rect -11882 1983 -11836 2021
rect -11882 1949 -11876 1983
rect -11842 1949 -11836 1983
rect -11882 1911 -11836 1949
rect -11882 1877 -11876 1911
rect -11842 1877 -11836 1911
rect -11882 1862 -11836 1877
rect -11670 2857 -11624 2872
rect -11670 2823 -11664 2857
rect -11630 2823 -11624 2857
rect -11670 2785 -11624 2823
rect -11670 2751 -11664 2785
rect -11630 2751 -11624 2785
rect -11670 2713 -11624 2751
rect -11670 2679 -11664 2713
rect -11630 2679 -11624 2713
rect -11670 2641 -11624 2679
rect -11670 2607 -11664 2641
rect -11630 2607 -11624 2641
rect -11670 2569 -11624 2607
rect -11670 2535 -11664 2569
rect -11630 2535 -11624 2569
rect -11670 2497 -11624 2535
rect -11670 2463 -11664 2497
rect -11630 2463 -11624 2497
rect -11670 2425 -11624 2463
rect -11670 2391 -11664 2425
rect -11630 2391 -11624 2425
rect -11670 2353 -11624 2391
rect -11670 2319 -11664 2353
rect -11630 2319 -11624 2353
rect -11670 2281 -11624 2319
rect -11670 2247 -11664 2281
rect -11630 2247 -11624 2281
rect -11670 2209 -11624 2247
rect -11670 2175 -11664 2209
rect -11630 2175 -11624 2209
rect -11670 2137 -11624 2175
rect -11670 2103 -11664 2137
rect -11630 2103 -11624 2137
rect -11670 2065 -11624 2103
rect -11670 2031 -11664 2065
rect -11630 2031 -11624 2065
rect -11670 1993 -11624 2031
rect -11670 1959 -11664 1993
rect -11630 1959 -11624 1993
rect -11670 1921 -11624 1959
rect -11670 1887 -11664 1921
rect -11630 1887 -11624 1921
rect -11670 1872 -11624 1887
rect -11574 2857 -11528 2872
rect -11574 2823 -11568 2857
rect -11534 2823 -11528 2857
rect -11574 2785 -11528 2823
rect -11574 2751 -11568 2785
rect -11534 2751 -11528 2785
rect -11574 2713 -11528 2751
rect -11574 2679 -11568 2713
rect -11534 2679 -11528 2713
rect -11574 2641 -11528 2679
rect -11574 2607 -11568 2641
rect -11534 2607 -11528 2641
rect -11574 2569 -11528 2607
rect -11574 2535 -11568 2569
rect -11534 2535 -11528 2569
rect -11574 2497 -11528 2535
rect -11574 2463 -11568 2497
rect -11534 2463 -11528 2497
rect -11574 2425 -11528 2463
rect -11574 2391 -11568 2425
rect -11534 2391 -11528 2425
rect -11574 2353 -11528 2391
rect -11574 2319 -11568 2353
rect -11534 2319 -11528 2353
rect -11574 2281 -11528 2319
rect -11574 2247 -11568 2281
rect -11534 2247 -11528 2281
rect -11574 2209 -11528 2247
rect -11574 2175 -11568 2209
rect -11534 2175 -11528 2209
rect -11574 2137 -11528 2175
rect -11574 2103 -11568 2137
rect -11534 2103 -11528 2137
rect -11574 2065 -11528 2103
rect -11574 2031 -11568 2065
rect -11534 2031 -11528 2065
rect -11574 1993 -11528 2031
rect -11574 1959 -11568 1993
rect -11534 1959 -11528 1993
rect -11574 1921 -11528 1959
rect -11574 1887 -11568 1921
rect -11534 1887 -11528 1921
rect -11574 1872 -11528 1887
rect -11478 2857 -11432 2872
rect -11478 2823 -11472 2857
rect -11438 2823 -11432 2857
rect -11478 2785 -11432 2823
rect -11478 2751 -11472 2785
rect -11438 2751 -11432 2785
rect -11478 2713 -11432 2751
rect -11478 2679 -11472 2713
rect -11438 2679 -11432 2713
rect -11478 2641 -11432 2679
rect -11478 2607 -11472 2641
rect -11438 2607 -11432 2641
rect -11478 2569 -11432 2607
rect -11478 2535 -11472 2569
rect -11438 2535 -11432 2569
rect -11478 2497 -11432 2535
rect -11478 2463 -11472 2497
rect -11438 2463 -11432 2497
rect -11478 2425 -11432 2463
rect -11478 2391 -11472 2425
rect -11438 2391 -11432 2425
rect -11478 2353 -11432 2391
rect -11478 2319 -11472 2353
rect -11438 2319 -11432 2353
rect -11478 2281 -11432 2319
rect -11478 2247 -11472 2281
rect -11438 2247 -11432 2281
rect -11478 2209 -11432 2247
rect -11478 2175 -11472 2209
rect -11438 2175 -11432 2209
rect -11478 2137 -11432 2175
rect -11478 2103 -11472 2137
rect -11438 2103 -11432 2137
rect -11478 2065 -11432 2103
rect -11478 2031 -11472 2065
rect -11438 2031 -11432 2065
rect -11478 1993 -11432 2031
rect -11478 1959 -11472 1993
rect -11438 1959 -11432 1993
rect -11478 1921 -11432 1959
rect -11478 1887 -11472 1921
rect -11438 1887 -11432 1921
rect -11478 1872 -11432 1887
rect -11382 2857 -11336 2872
rect -11382 2823 -11376 2857
rect -11342 2823 -11336 2857
rect -11382 2785 -11336 2823
rect -11382 2751 -11376 2785
rect -11342 2751 -11336 2785
rect -11382 2713 -11336 2751
rect -11382 2679 -11376 2713
rect -11342 2679 -11336 2713
rect -11382 2641 -11336 2679
rect -11382 2607 -11376 2641
rect -11342 2607 -11336 2641
rect -11382 2569 -11336 2607
rect -11382 2535 -11376 2569
rect -11342 2535 -11336 2569
rect -11382 2497 -11336 2535
rect -11382 2463 -11376 2497
rect -11342 2463 -11336 2497
rect -11382 2425 -11336 2463
rect -11382 2391 -11376 2425
rect -11342 2391 -11336 2425
rect -11382 2353 -11336 2391
rect -11382 2319 -11376 2353
rect -11342 2319 -11336 2353
rect -11382 2281 -11336 2319
rect -11382 2247 -11376 2281
rect -11342 2247 -11336 2281
rect -11382 2209 -11336 2247
rect -11382 2175 -11376 2209
rect -11342 2175 -11336 2209
rect -11382 2137 -11336 2175
rect -11382 2103 -11376 2137
rect -11342 2103 -11336 2137
rect -11382 2065 -11336 2103
rect -11382 2031 -11376 2065
rect -11342 2031 -11336 2065
rect -11382 1993 -11336 2031
rect -11382 1959 -11376 1993
rect -11342 1959 -11336 1993
rect -11382 1921 -11336 1959
rect -11382 1887 -11376 1921
rect -11342 1887 -11336 1921
rect -11382 1872 -11336 1887
rect -11286 2857 -11240 2872
rect -11286 2823 -11280 2857
rect -11246 2823 -11240 2857
rect -11286 2785 -11240 2823
rect -11286 2751 -11280 2785
rect -11246 2751 -11240 2785
rect -11286 2713 -11240 2751
rect -11286 2679 -11280 2713
rect -11246 2679 -11240 2713
rect -11286 2641 -11240 2679
rect -11286 2607 -11280 2641
rect -11246 2607 -11240 2641
rect -11286 2569 -11240 2607
rect -11286 2535 -11280 2569
rect -11246 2535 -11240 2569
rect -11286 2497 -11240 2535
rect -11286 2463 -11280 2497
rect -11246 2463 -11240 2497
rect -11286 2425 -11240 2463
rect -11286 2391 -11280 2425
rect -11246 2391 -11240 2425
rect -11286 2353 -11240 2391
rect -11286 2319 -11280 2353
rect -11246 2319 -11240 2353
rect -11286 2281 -11240 2319
rect -11286 2247 -11280 2281
rect -11246 2247 -11240 2281
rect -11286 2209 -11240 2247
rect -11286 2175 -11280 2209
rect -11246 2175 -11240 2209
rect -11286 2137 -11240 2175
rect -11286 2103 -11280 2137
rect -11246 2103 -11240 2137
rect -11286 2065 -11240 2103
rect -11286 2031 -11280 2065
rect -11246 2031 -11240 2065
rect -11286 1993 -11240 2031
rect -11286 1959 -11280 1993
rect -11246 1959 -11240 1993
rect -11286 1921 -11240 1959
rect -11286 1887 -11280 1921
rect -11246 1887 -11240 1921
rect -11286 1872 -11240 1887
rect -11190 2857 -11144 2872
rect -11190 2823 -11184 2857
rect -11150 2823 -11144 2857
rect -11190 2785 -11144 2823
rect -11190 2751 -11184 2785
rect -11150 2751 -11144 2785
rect -11190 2713 -11144 2751
rect -11190 2679 -11184 2713
rect -11150 2679 -11144 2713
rect -11190 2641 -11144 2679
rect -11190 2607 -11184 2641
rect -11150 2607 -11144 2641
rect -11190 2569 -11144 2607
rect -11190 2535 -11184 2569
rect -11150 2535 -11144 2569
rect -11190 2497 -11144 2535
rect -11190 2463 -11184 2497
rect -11150 2463 -11144 2497
rect -11190 2425 -11144 2463
rect -11190 2391 -11184 2425
rect -11150 2391 -11144 2425
rect -11190 2353 -11144 2391
rect -11190 2319 -11184 2353
rect -11150 2319 -11144 2353
rect -11190 2281 -11144 2319
rect -11190 2247 -11184 2281
rect -11150 2247 -11144 2281
rect -11190 2209 -11144 2247
rect -11190 2175 -11184 2209
rect -11150 2175 -11144 2209
rect -11190 2137 -11144 2175
rect -11190 2103 -11184 2137
rect -11150 2103 -11144 2137
rect -11190 2065 -11144 2103
rect -11190 2031 -11184 2065
rect -11150 2031 -11144 2065
rect -11190 1993 -11144 2031
rect -11190 1959 -11184 1993
rect -11150 1959 -11144 1993
rect -11190 1921 -11144 1959
rect -11190 1887 -11184 1921
rect -11150 1887 -11144 1921
rect -11190 1872 -11144 1887
rect -16644 1677 -16266 1680
rect -16644 1497 -16609 1677
rect -16301 1497 -16266 1677
rect -16644 1494 -16266 1497
rect -14442 1678 -14068 1680
rect -14442 1498 -14409 1678
rect -14101 1498 -14068 1678
rect -14442 1496 -14068 1498
rect -12042 1677 -11664 1680
rect -12042 1497 -12007 1677
rect -11699 1497 -11664 1677
rect -12042 1494 -11664 1497
rect -10698 -5914 -10398 3086
rect -8458 3084 -7388 3108
rect -6786 3155 -5734 3186
rect -6786 3121 -5822 3155
rect -5788 3121 -5734 3155
rect -6786 3090 -5734 3121
rect -5576 3176 -5496 3263
rect -4892 3279 -4794 3306
rect -4892 3245 -4862 3279
rect -4828 3245 -4794 3279
rect -4892 3182 -4794 3245
rect -5576 3157 -4944 3176
rect -5576 3123 -5006 3157
rect -4972 3123 -4944 3157
rect -5576 3106 -4944 3123
rect -4892 3151 -4448 3182
rect -8458 3026 -8346 3084
rect -8458 2992 -8420 3026
rect -8386 2992 -8346 3026
rect -8458 2952 -8346 2992
rect -6786 3028 -6686 3090
rect -6786 2994 -6752 3028
rect -6718 2994 -6686 3028
rect -5576 3072 -5496 3106
rect -5576 3038 -5554 3072
rect -5520 3038 -5496 3072
rect -5576 3016 -5496 3038
rect -4892 3099 -4538 3151
rect -4486 3099 -4448 3151
rect -4892 3078 -4448 3099
rect -4892 3042 -4794 3078
rect -4576 3068 -4448 3078
rect -6786 2968 -6686 2994
rect -4892 3008 -4862 3042
rect -4828 3008 -4794 3042
rect -4892 2982 -4794 3008
rect -10202 2849 -10156 2864
rect -10202 2815 -10196 2849
rect -10162 2815 -10156 2849
rect -10202 2777 -10156 2815
rect -10202 2743 -10196 2777
rect -10162 2743 -10156 2777
rect -10202 2705 -10156 2743
rect -10202 2671 -10196 2705
rect -10162 2671 -10156 2705
rect -10202 2633 -10156 2671
rect -10202 2599 -10196 2633
rect -10162 2599 -10156 2633
rect -10202 2561 -10156 2599
rect -10202 2527 -10196 2561
rect -10162 2527 -10156 2561
rect -10202 2489 -10156 2527
rect -10202 2455 -10196 2489
rect -10162 2455 -10156 2489
rect -10202 2417 -10156 2455
rect -10202 2383 -10196 2417
rect -10162 2383 -10156 2417
rect -10202 2345 -10156 2383
rect -10202 2311 -10196 2345
rect -10162 2311 -10156 2345
rect -10202 2273 -10156 2311
rect -10202 2239 -10196 2273
rect -10162 2239 -10156 2273
rect -10202 2201 -10156 2239
rect -10202 2167 -10196 2201
rect -10162 2167 -10156 2201
rect -10202 2129 -10156 2167
rect -10202 2095 -10196 2129
rect -10162 2095 -10156 2129
rect -10202 2057 -10156 2095
rect -10202 2023 -10196 2057
rect -10162 2023 -10156 2057
rect -10202 1985 -10156 2023
rect -10202 1951 -10196 1985
rect -10162 1951 -10156 1985
rect -10202 1913 -10156 1951
rect -10202 1879 -10196 1913
rect -10162 1879 -10156 1913
rect -10202 1864 -10156 1879
rect -10106 2849 -10060 2864
rect -10106 2815 -10100 2849
rect -10066 2815 -10060 2849
rect -10106 2777 -10060 2815
rect -10106 2743 -10100 2777
rect -10066 2743 -10060 2777
rect -10106 2705 -10060 2743
rect -10106 2671 -10100 2705
rect -10066 2671 -10060 2705
rect -10106 2633 -10060 2671
rect -10106 2599 -10100 2633
rect -10066 2599 -10060 2633
rect -10106 2561 -10060 2599
rect -10106 2527 -10100 2561
rect -10066 2527 -10060 2561
rect -10106 2489 -10060 2527
rect -10106 2455 -10100 2489
rect -10066 2455 -10060 2489
rect -10106 2417 -10060 2455
rect -10106 2383 -10100 2417
rect -10066 2383 -10060 2417
rect -10106 2345 -10060 2383
rect -10106 2311 -10100 2345
rect -10066 2311 -10060 2345
rect -10106 2273 -10060 2311
rect -10106 2239 -10100 2273
rect -10066 2239 -10060 2273
rect -10106 2201 -10060 2239
rect -10106 2167 -10100 2201
rect -10066 2167 -10060 2201
rect -10106 2129 -10060 2167
rect -10106 2095 -10100 2129
rect -10066 2095 -10060 2129
rect -10106 2057 -10060 2095
rect -10106 2023 -10100 2057
rect -10066 2023 -10060 2057
rect -10106 1985 -10060 2023
rect -10106 1951 -10100 1985
rect -10066 1951 -10060 1985
rect -10106 1913 -10060 1951
rect -10106 1879 -10100 1913
rect -10066 1879 -10060 1913
rect -10106 1864 -10060 1879
rect -10010 2849 -9964 2864
rect -10010 2815 -10004 2849
rect -9970 2815 -9964 2849
rect -10010 2777 -9964 2815
rect -10010 2743 -10004 2777
rect -9970 2743 -9964 2777
rect -10010 2705 -9964 2743
rect -10010 2671 -10004 2705
rect -9970 2671 -9964 2705
rect -10010 2633 -9964 2671
rect -10010 2599 -10004 2633
rect -9970 2599 -9964 2633
rect -10010 2561 -9964 2599
rect -10010 2527 -10004 2561
rect -9970 2527 -9964 2561
rect -10010 2489 -9964 2527
rect -10010 2455 -10004 2489
rect -9970 2455 -9964 2489
rect -10010 2417 -9964 2455
rect -10010 2383 -10004 2417
rect -9970 2383 -9964 2417
rect -10010 2345 -9964 2383
rect -10010 2311 -10004 2345
rect -9970 2311 -9964 2345
rect -10010 2273 -9964 2311
rect -10010 2239 -10004 2273
rect -9970 2239 -9964 2273
rect -10010 2201 -9964 2239
rect -10010 2167 -10004 2201
rect -9970 2167 -9964 2201
rect -10010 2129 -9964 2167
rect -10010 2095 -10004 2129
rect -9970 2095 -9964 2129
rect -10010 2057 -9964 2095
rect -10010 2023 -10004 2057
rect -9970 2023 -9964 2057
rect -10010 1985 -9964 2023
rect -10010 1951 -10004 1985
rect -9970 1951 -9964 1985
rect -10010 1913 -9964 1951
rect -10010 1879 -10004 1913
rect -9970 1879 -9964 1913
rect -10010 1864 -9964 1879
rect -9914 2849 -9868 2864
rect -9914 2815 -9908 2849
rect -9874 2815 -9868 2849
rect -9914 2777 -9868 2815
rect -9914 2743 -9908 2777
rect -9874 2743 -9868 2777
rect -9914 2705 -9868 2743
rect -9914 2671 -9908 2705
rect -9874 2671 -9868 2705
rect -9914 2633 -9868 2671
rect -9914 2599 -9908 2633
rect -9874 2599 -9868 2633
rect -9914 2561 -9868 2599
rect -9914 2527 -9908 2561
rect -9874 2527 -9868 2561
rect -9914 2489 -9868 2527
rect -9914 2455 -9908 2489
rect -9874 2455 -9868 2489
rect -9914 2417 -9868 2455
rect -9914 2383 -9908 2417
rect -9874 2383 -9868 2417
rect -9914 2345 -9868 2383
rect -9914 2311 -9908 2345
rect -9874 2311 -9868 2345
rect -9914 2273 -9868 2311
rect -9914 2239 -9908 2273
rect -9874 2239 -9868 2273
rect -9914 2201 -9868 2239
rect -9914 2167 -9908 2201
rect -9874 2167 -9868 2201
rect -9914 2129 -9868 2167
rect -9914 2095 -9908 2129
rect -9874 2095 -9868 2129
rect -9914 2057 -9868 2095
rect -9914 2023 -9908 2057
rect -9874 2023 -9868 2057
rect -9914 1985 -9868 2023
rect -9914 1951 -9908 1985
rect -9874 1951 -9868 1985
rect -9914 1913 -9868 1951
rect -9914 1879 -9908 1913
rect -9874 1879 -9868 1913
rect -9914 1864 -9868 1879
rect -9818 2849 -9772 2864
rect -9818 2815 -9812 2849
rect -9778 2815 -9772 2849
rect -9818 2777 -9772 2815
rect -9818 2743 -9812 2777
rect -9778 2743 -9772 2777
rect -9818 2705 -9772 2743
rect -9818 2671 -9812 2705
rect -9778 2671 -9772 2705
rect -9818 2633 -9772 2671
rect -9818 2599 -9812 2633
rect -9778 2599 -9772 2633
rect -9818 2561 -9772 2599
rect -9818 2527 -9812 2561
rect -9778 2527 -9772 2561
rect -9818 2489 -9772 2527
rect -9818 2455 -9812 2489
rect -9778 2455 -9772 2489
rect -9818 2417 -9772 2455
rect -9818 2383 -9812 2417
rect -9778 2383 -9772 2417
rect -9818 2345 -9772 2383
rect -9818 2311 -9812 2345
rect -9778 2311 -9772 2345
rect -9818 2273 -9772 2311
rect -9818 2239 -9812 2273
rect -9778 2239 -9772 2273
rect -9818 2201 -9772 2239
rect -9818 2167 -9812 2201
rect -9778 2167 -9772 2201
rect -9818 2129 -9772 2167
rect -9818 2095 -9812 2129
rect -9778 2095 -9772 2129
rect -9818 2057 -9772 2095
rect -9818 2023 -9812 2057
rect -9778 2023 -9772 2057
rect -9818 1985 -9772 2023
rect -9818 1951 -9812 1985
rect -9778 1951 -9772 1985
rect -9818 1913 -9772 1951
rect -9818 1879 -9812 1913
rect -9778 1879 -9772 1913
rect -9818 1864 -9772 1879
rect -9722 2849 -9676 2864
rect -9722 2815 -9716 2849
rect -9682 2815 -9676 2849
rect -9722 2777 -9676 2815
rect -9722 2743 -9716 2777
rect -9682 2743 -9676 2777
rect -9722 2705 -9676 2743
rect -9722 2671 -9716 2705
rect -9682 2671 -9676 2705
rect -9722 2633 -9676 2671
rect -9722 2599 -9716 2633
rect -9682 2599 -9676 2633
rect -9722 2561 -9676 2599
rect -9722 2527 -9716 2561
rect -9682 2527 -9676 2561
rect -9722 2489 -9676 2527
rect -9722 2455 -9716 2489
rect -9682 2455 -9676 2489
rect -9722 2417 -9676 2455
rect -9722 2383 -9716 2417
rect -9682 2383 -9676 2417
rect -9722 2345 -9676 2383
rect -9722 2311 -9716 2345
rect -9682 2311 -9676 2345
rect -9722 2273 -9676 2311
rect -9722 2239 -9716 2273
rect -9682 2239 -9676 2273
rect -9722 2201 -9676 2239
rect -9722 2167 -9716 2201
rect -9682 2167 -9676 2201
rect -9722 2129 -9676 2167
rect -9722 2095 -9716 2129
rect -9682 2095 -9676 2129
rect -9722 2057 -9676 2095
rect -9722 2023 -9716 2057
rect -9682 2023 -9676 2057
rect -9722 1985 -9676 2023
rect -9722 1951 -9716 1985
rect -9682 1951 -9676 1985
rect -9722 1913 -9676 1951
rect -9722 1879 -9716 1913
rect -9682 1879 -9676 1913
rect -9722 1864 -9676 1879
rect -9626 2849 -9580 2864
rect -9626 2815 -9620 2849
rect -9586 2815 -9580 2849
rect -9626 2777 -9580 2815
rect -9626 2743 -9620 2777
rect -9586 2743 -9580 2777
rect -9626 2705 -9580 2743
rect -9626 2671 -9620 2705
rect -9586 2671 -9580 2705
rect -9626 2633 -9580 2671
rect -9626 2599 -9620 2633
rect -9586 2599 -9580 2633
rect -9626 2561 -9580 2599
rect -9626 2527 -9620 2561
rect -9586 2527 -9580 2561
rect -9626 2489 -9580 2527
rect -9626 2455 -9620 2489
rect -9586 2455 -9580 2489
rect -9626 2417 -9580 2455
rect -9626 2383 -9620 2417
rect -9586 2383 -9580 2417
rect -9626 2345 -9580 2383
rect -9626 2311 -9620 2345
rect -9586 2311 -9580 2345
rect -9626 2273 -9580 2311
rect -9626 2239 -9620 2273
rect -9586 2239 -9580 2273
rect -9626 2201 -9580 2239
rect -9626 2167 -9620 2201
rect -9586 2167 -9580 2201
rect -9626 2129 -9580 2167
rect -9626 2095 -9620 2129
rect -9586 2095 -9580 2129
rect -9626 2057 -9580 2095
rect -9626 2023 -9620 2057
rect -9586 2023 -9580 2057
rect -9626 1985 -9580 2023
rect -9626 1951 -9620 1985
rect -9586 1951 -9580 1985
rect -9626 1913 -9580 1951
rect -9626 1879 -9620 1913
rect -9586 1879 -9580 1913
rect -9626 1864 -9580 1879
rect -9530 2849 -9484 2864
rect -9530 2815 -9524 2849
rect -9490 2815 -9484 2849
rect -9530 2777 -9484 2815
rect -9530 2743 -9524 2777
rect -9490 2743 -9484 2777
rect -9530 2705 -9484 2743
rect -9530 2671 -9524 2705
rect -9490 2671 -9484 2705
rect -9530 2633 -9484 2671
rect -9530 2599 -9524 2633
rect -9490 2599 -9484 2633
rect -9530 2561 -9484 2599
rect -9530 2527 -9524 2561
rect -9490 2527 -9484 2561
rect -9530 2489 -9484 2527
rect -9530 2455 -9524 2489
rect -9490 2455 -9484 2489
rect -9530 2417 -9484 2455
rect -9530 2383 -9524 2417
rect -9490 2383 -9484 2417
rect -9530 2345 -9484 2383
rect -9530 2311 -9524 2345
rect -9490 2311 -9484 2345
rect -9530 2273 -9484 2311
rect -9530 2239 -9524 2273
rect -9490 2239 -9484 2273
rect -9530 2201 -9484 2239
rect -9530 2167 -9524 2201
rect -9490 2167 -9484 2201
rect -9530 2129 -9484 2167
rect -9530 2095 -9524 2129
rect -9490 2095 -9484 2129
rect -9530 2057 -9484 2095
rect -9530 2023 -9524 2057
rect -9490 2023 -9484 2057
rect -9530 1985 -9484 2023
rect -9530 1951 -9524 1985
rect -9490 1951 -9484 1985
rect -9530 1913 -9484 1951
rect -9530 1879 -9524 1913
rect -9490 1879 -9484 1913
rect -9530 1864 -9484 1879
rect -9434 2849 -9388 2864
rect -9434 2815 -9428 2849
rect -9394 2815 -9388 2849
rect -9434 2777 -9388 2815
rect -9434 2743 -9428 2777
rect -9394 2743 -9388 2777
rect -9434 2705 -9388 2743
rect -9434 2671 -9428 2705
rect -9394 2671 -9388 2705
rect -9434 2633 -9388 2671
rect -9434 2599 -9428 2633
rect -9394 2599 -9388 2633
rect -9434 2561 -9388 2599
rect -9434 2527 -9428 2561
rect -9394 2527 -9388 2561
rect -9434 2489 -9388 2527
rect -9434 2455 -9428 2489
rect -9394 2455 -9388 2489
rect -9434 2417 -9388 2455
rect -9434 2383 -9428 2417
rect -9394 2383 -9388 2417
rect -9434 2345 -9388 2383
rect -9434 2311 -9428 2345
rect -9394 2311 -9388 2345
rect -9434 2273 -9388 2311
rect -9434 2239 -9428 2273
rect -9394 2239 -9388 2273
rect -9434 2201 -9388 2239
rect -9434 2167 -9428 2201
rect -9394 2167 -9388 2201
rect -9434 2129 -9388 2167
rect -9434 2095 -9428 2129
rect -9394 2095 -9388 2129
rect -9434 2057 -9388 2095
rect -9434 2023 -9428 2057
rect -9394 2023 -9388 2057
rect -9434 1985 -9388 2023
rect -9434 1951 -9428 1985
rect -9394 1951 -9388 1985
rect -9434 1913 -9388 1951
rect -9434 1879 -9428 1913
rect -9394 1879 -9388 1913
rect -9434 1864 -9388 1879
rect -9338 2849 -9292 2864
rect -9338 2815 -9332 2849
rect -9298 2815 -9292 2849
rect -9338 2777 -9292 2815
rect -9338 2743 -9332 2777
rect -9298 2743 -9292 2777
rect -9338 2705 -9292 2743
rect -9338 2671 -9332 2705
rect -9298 2671 -9292 2705
rect -9338 2633 -9292 2671
rect -9338 2599 -9332 2633
rect -9298 2599 -9292 2633
rect -9338 2561 -9292 2599
rect -9338 2527 -9332 2561
rect -9298 2527 -9292 2561
rect -9338 2489 -9292 2527
rect -9338 2455 -9332 2489
rect -9298 2455 -9292 2489
rect -9338 2417 -9292 2455
rect -9338 2383 -9332 2417
rect -9298 2383 -9292 2417
rect -9338 2345 -9292 2383
rect -9338 2311 -9332 2345
rect -9298 2311 -9292 2345
rect -9338 2273 -9292 2311
rect -9338 2239 -9332 2273
rect -9298 2239 -9292 2273
rect -9338 2201 -9292 2239
rect -9338 2167 -9332 2201
rect -9298 2167 -9292 2201
rect -9338 2129 -9292 2167
rect -9338 2095 -9332 2129
rect -9298 2095 -9292 2129
rect -9338 2057 -9292 2095
rect -9338 2023 -9332 2057
rect -9298 2023 -9292 2057
rect -9338 1985 -9292 2023
rect -9338 1951 -9332 1985
rect -9298 1951 -9292 1985
rect -9338 1913 -9292 1951
rect -9338 1879 -9332 1913
rect -9298 1879 -9292 1913
rect -9338 1864 -9292 1879
rect -9242 2849 -9196 2864
rect -9242 2815 -9236 2849
rect -9202 2815 -9196 2849
rect -9242 2777 -9196 2815
rect -9242 2743 -9236 2777
rect -9202 2743 -9196 2777
rect -9242 2705 -9196 2743
rect -9242 2671 -9236 2705
rect -9202 2671 -9196 2705
rect -9242 2633 -9196 2671
rect -9242 2599 -9236 2633
rect -9202 2599 -9196 2633
rect -9242 2561 -9196 2599
rect -9242 2527 -9236 2561
rect -9202 2527 -9196 2561
rect -9242 2489 -9196 2527
rect -9242 2455 -9236 2489
rect -9202 2455 -9196 2489
rect -9242 2417 -9196 2455
rect -9242 2383 -9236 2417
rect -9202 2383 -9196 2417
rect -9242 2345 -9196 2383
rect -9242 2311 -9236 2345
rect -9202 2311 -9196 2345
rect -9242 2273 -9196 2311
rect -9242 2239 -9236 2273
rect -9202 2239 -9196 2273
rect -9242 2201 -9196 2239
rect -9242 2167 -9236 2201
rect -9202 2167 -9196 2201
rect -9242 2129 -9196 2167
rect -9242 2095 -9236 2129
rect -9202 2095 -9196 2129
rect -9242 2057 -9196 2095
rect -9242 2023 -9236 2057
rect -9202 2023 -9196 2057
rect -9242 1985 -9196 2023
rect -9242 1951 -9236 1985
rect -9202 1951 -9196 1985
rect -9242 1913 -9196 1951
rect -9242 1879 -9236 1913
rect -9202 1879 -9196 1913
rect -9242 1864 -9196 1879
rect -9146 2849 -9100 2864
rect -9146 2815 -9140 2849
rect -9106 2815 -9100 2849
rect -9146 2777 -9100 2815
rect -9146 2743 -9140 2777
rect -9106 2743 -9100 2777
rect -9146 2705 -9100 2743
rect -9146 2671 -9140 2705
rect -9106 2671 -9100 2705
rect -9146 2633 -9100 2671
rect -9146 2599 -9140 2633
rect -9106 2599 -9100 2633
rect -9146 2561 -9100 2599
rect -9146 2527 -9140 2561
rect -9106 2527 -9100 2561
rect -9146 2489 -9100 2527
rect -9146 2455 -9140 2489
rect -9106 2455 -9100 2489
rect -9146 2417 -9100 2455
rect -9146 2383 -9140 2417
rect -9106 2383 -9100 2417
rect -9146 2345 -9100 2383
rect -9146 2311 -9140 2345
rect -9106 2311 -9100 2345
rect -9146 2273 -9100 2311
rect -9146 2239 -9140 2273
rect -9106 2239 -9100 2273
rect -9146 2201 -9100 2239
rect -9146 2167 -9140 2201
rect -9106 2167 -9100 2201
rect -9146 2129 -9100 2167
rect -9146 2095 -9140 2129
rect -9106 2095 -9100 2129
rect -9146 2057 -9100 2095
rect -9146 2023 -9140 2057
rect -9106 2023 -9100 2057
rect -9146 1985 -9100 2023
rect -9146 1951 -9140 1985
rect -9106 1951 -9100 1985
rect -9146 1913 -9100 1951
rect -9146 1879 -9140 1913
rect -9106 1879 -9100 1913
rect -9146 1864 -9100 1879
rect -9050 2849 -9004 2864
rect -9050 2815 -9044 2849
rect -9010 2815 -9004 2849
rect -9050 2777 -9004 2815
rect -9050 2743 -9044 2777
rect -9010 2743 -9004 2777
rect -9050 2705 -9004 2743
rect -9050 2671 -9044 2705
rect -9010 2671 -9004 2705
rect -9050 2633 -9004 2671
rect -9050 2599 -9044 2633
rect -9010 2599 -9004 2633
rect -9050 2561 -9004 2599
rect -9050 2527 -9044 2561
rect -9010 2527 -9004 2561
rect -9050 2489 -9004 2527
rect -9050 2455 -9044 2489
rect -9010 2455 -9004 2489
rect -9050 2417 -9004 2455
rect -9050 2383 -9044 2417
rect -9010 2383 -9004 2417
rect -9050 2345 -9004 2383
rect -9050 2311 -9044 2345
rect -9010 2311 -9004 2345
rect -9050 2273 -9004 2311
rect -9050 2239 -9044 2273
rect -9010 2239 -9004 2273
rect -9050 2201 -9004 2239
rect -9050 2167 -9044 2201
rect -9010 2167 -9004 2201
rect -9050 2129 -9004 2167
rect -9050 2095 -9044 2129
rect -9010 2095 -9004 2129
rect -9050 2057 -9004 2095
rect -9050 2023 -9044 2057
rect -9010 2023 -9004 2057
rect -9050 1985 -9004 2023
rect -9050 1951 -9044 1985
rect -9010 1951 -9004 1985
rect -9050 1913 -9004 1951
rect -9050 1879 -9044 1913
rect -9010 1879 -9004 1913
rect -9050 1864 -9004 1879
rect -8954 2849 -8908 2864
rect -8954 2815 -8948 2849
rect -8914 2815 -8908 2849
rect -8954 2777 -8908 2815
rect -8954 2743 -8948 2777
rect -8914 2743 -8908 2777
rect -8954 2705 -8908 2743
rect -8954 2671 -8948 2705
rect -8914 2671 -8908 2705
rect -8954 2633 -8908 2671
rect -8954 2599 -8948 2633
rect -8914 2599 -8908 2633
rect -8954 2561 -8908 2599
rect -8954 2527 -8948 2561
rect -8914 2527 -8908 2561
rect -8954 2489 -8908 2527
rect -8954 2455 -8948 2489
rect -8914 2455 -8908 2489
rect -8954 2417 -8908 2455
rect -8954 2383 -8948 2417
rect -8914 2383 -8908 2417
rect -8954 2345 -8908 2383
rect -8954 2311 -8948 2345
rect -8914 2311 -8908 2345
rect -8954 2273 -8908 2311
rect -8954 2239 -8948 2273
rect -8914 2239 -8908 2273
rect -8954 2201 -8908 2239
rect -8954 2167 -8948 2201
rect -8914 2167 -8908 2201
rect -8954 2129 -8908 2167
rect -8954 2095 -8948 2129
rect -8914 2095 -8908 2129
rect -8954 2057 -8908 2095
rect -8954 2023 -8948 2057
rect -8914 2023 -8908 2057
rect -8954 1985 -8908 2023
rect -8954 1951 -8948 1985
rect -8914 1951 -8908 1985
rect -8954 1913 -8908 1951
rect -8954 1879 -8948 1913
rect -8914 1879 -8908 1913
rect -8954 1864 -8908 1879
rect -8858 2849 -8812 2864
rect -8858 2815 -8852 2849
rect -8818 2815 -8812 2849
rect -8858 2777 -8812 2815
rect -8858 2743 -8852 2777
rect -8818 2743 -8812 2777
rect -8858 2705 -8812 2743
rect -8858 2671 -8852 2705
rect -8818 2671 -8812 2705
rect -8858 2633 -8812 2671
rect -8858 2599 -8852 2633
rect -8818 2599 -8812 2633
rect -8858 2561 -8812 2599
rect -8858 2527 -8852 2561
rect -8818 2527 -8812 2561
rect -8858 2489 -8812 2527
rect -8858 2455 -8852 2489
rect -8818 2455 -8812 2489
rect -8858 2417 -8812 2455
rect -8858 2383 -8852 2417
rect -8818 2383 -8812 2417
rect -8858 2345 -8812 2383
rect -8858 2311 -8852 2345
rect -8818 2311 -8812 2345
rect -8858 2273 -8812 2311
rect -8858 2239 -8852 2273
rect -8818 2239 -8812 2273
rect -8858 2201 -8812 2239
rect -8858 2167 -8852 2201
rect -8818 2167 -8812 2201
rect -8858 2129 -8812 2167
rect -8858 2095 -8852 2129
rect -8818 2095 -8812 2129
rect -8858 2057 -8812 2095
rect -8858 2023 -8852 2057
rect -8818 2023 -8812 2057
rect -8858 1985 -8812 2023
rect -8858 1951 -8852 1985
rect -8818 1951 -8812 1985
rect -8858 1913 -8812 1951
rect -8858 1879 -8852 1913
rect -8818 1879 -8812 1913
rect -8858 1864 -8812 1879
rect -8762 2849 -8716 2864
rect -8762 2815 -8756 2849
rect -8722 2815 -8716 2849
rect -8762 2777 -8716 2815
rect -8762 2743 -8756 2777
rect -8722 2743 -8716 2777
rect -8762 2705 -8716 2743
rect -8762 2671 -8756 2705
rect -8722 2671 -8716 2705
rect -8762 2633 -8716 2671
rect -8762 2599 -8756 2633
rect -8722 2599 -8716 2633
rect -8762 2561 -8716 2599
rect -8762 2527 -8756 2561
rect -8722 2527 -8716 2561
rect -8762 2489 -8716 2527
rect -8762 2455 -8756 2489
rect -8722 2455 -8716 2489
rect -8762 2417 -8716 2455
rect -8762 2383 -8756 2417
rect -8722 2383 -8716 2417
rect -8762 2345 -8716 2383
rect -8762 2311 -8756 2345
rect -8722 2311 -8716 2345
rect -8762 2273 -8716 2311
rect -8762 2239 -8756 2273
rect -8722 2239 -8716 2273
rect -8762 2201 -8716 2239
rect -8762 2167 -8756 2201
rect -8722 2167 -8716 2201
rect -8762 2129 -8716 2167
rect -8762 2095 -8756 2129
rect -8722 2095 -8716 2129
rect -8762 2057 -8716 2095
rect -8762 2023 -8756 2057
rect -8722 2023 -8716 2057
rect -8762 1985 -8716 2023
rect -8762 1951 -8756 1985
rect -8722 1951 -8716 1985
rect -8762 1913 -8716 1951
rect -8762 1879 -8756 1913
rect -8722 1879 -8716 1913
rect -8762 1864 -8716 1879
rect -8666 2849 -8620 2864
rect -8666 2815 -8660 2849
rect -8626 2815 -8620 2849
rect -8666 2777 -8620 2815
rect -8666 2743 -8660 2777
rect -8626 2743 -8620 2777
rect -8666 2705 -8620 2743
rect -8666 2671 -8660 2705
rect -8626 2671 -8620 2705
rect -8666 2633 -8620 2671
rect -8666 2599 -8660 2633
rect -8626 2599 -8620 2633
rect -8666 2561 -8620 2599
rect -8666 2527 -8660 2561
rect -8626 2527 -8620 2561
rect -8666 2489 -8620 2527
rect -8666 2455 -8660 2489
rect -8626 2455 -8620 2489
rect -8666 2417 -8620 2455
rect -8666 2383 -8660 2417
rect -8626 2383 -8620 2417
rect -8666 2345 -8620 2383
rect -8666 2311 -8660 2345
rect -8626 2311 -8620 2345
rect -8666 2273 -8620 2311
rect -8666 2239 -8660 2273
rect -8626 2239 -8620 2273
rect -8666 2201 -8620 2239
rect -8666 2167 -8660 2201
rect -8626 2167 -8620 2201
rect -8666 2129 -8620 2167
rect -8666 2095 -8660 2129
rect -8626 2095 -8620 2129
rect -8666 2057 -8620 2095
rect -8666 2023 -8660 2057
rect -8626 2023 -8620 2057
rect -8666 1985 -8620 2023
rect -8666 1951 -8660 1985
rect -8626 1951 -8620 1985
rect -8666 1913 -8620 1951
rect -8666 1879 -8660 1913
rect -8626 1879 -8620 1913
rect -8666 1864 -8620 1879
rect -8570 2849 -8524 2864
rect -8570 2815 -8564 2849
rect -8530 2815 -8524 2849
rect -8570 2777 -8524 2815
rect -8570 2743 -8564 2777
rect -8530 2743 -8524 2777
rect -8570 2705 -8524 2743
rect -8570 2671 -8564 2705
rect -8530 2671 -8524 2705
rect -8570 2633 -8524 2671
rect -8570 2599 -8564 2633
rect -8530 2599 -8524 2633
rect -8570 2561 -8524 2599
rect -8570 2527 -8564 2561
rect -8530 2527 -8524 2561
rect -8570 2489 -8524 2527
rect -8570 2455 -8564 2489
rect -8530 2455 -8524 2489
rect -8570 2417 -8524 2455
rect -8570 2383 -8564 2417
rect -8530 2383 -8524 2417
rect -8570 2345 -8524 2383
rect -8570 2311 -8564 2345
rect -8530 2311 -8524 2345
rect -8570 2273 -8524 2311
rect -8570 2239 -8564 2273
rect -8530 2239 -8524 2273
rect -8570 2201 -8524 2239
rect -8570 2167 -8564 2201
rect -8530 2167 -8524 2201
rect -8570 2129 -8524 2167
rect -8570 2095 -8564 2129
rect -8530 2095 -8524 2129
rect -8570 2057 -8524 2095
rect -8570 2023 -8564 2057
rect -8530 2023 -8524 2057
rect -8570 1985 -8524 2023
rect -8570 1951 -8564 1985
rect -8530 1951 -8524 1985
rect -8570 1913 -8524 1951
rect -8570 1879 -8564 1913
rect -8530 1879 -8524 1913
rect -8570 1864 -8524 1879
rect -8474 2849 -8428 2864
rect -8474 2815 -8468 2849
rect -8434 2815 -8428 2849
rect -8474 2777 -8428 2815
rect -8474 2743 -8468 2777
rect -8434 2743 -8428 2777
rect -8474 2705 -8428 2743
rect -8474 2671 -8468 2705
rect -8434 2671 -8428 2705
rect -8474 2633 -8428 2671
rect -8474 2599 -8468 2633
rect -8434 2599 -8428 2633
rect -8474 2561 -8428 2599
rect -8474 2527 -8468 2561
rect -8434 2527 -8428 2561
rect -8474 2489 -8428 2527
rect -8474 2455 -8468 2489
rect -8434 2455 -8428 2489
rect -8474 2417 -8428 2455
rect -8474 2383 -8468 2417
rect -8434 2383 -8428 2417
rect -8474 2345 -8428 2383
rect -8474 2311 -8468 2345
rect -8434 2311 -8428 2345
rect -8474 2273 -8428 2311
rect -8474 2239 -8468 2273
rect -8434 2239 -8428 2273
rect -8474 2201 -8428 2239
rect -8474 2167 -8468 2201
rect -8434 2167 -8428 2201
rect -8474 2129 -8428 2167
rect -8474 2095 -8468 2129
rect -8434 2095 -8428 2129
rect -8474 2057 -8428 2095
rect -8474 2023 -8468 2057
rect -8434 2023 -8428 2057
rect -8474 1985 -8428 2023
rect -8474 1951 -8468 1985
rect -8434 1951 -8428 1985
rect -8474 1913 -8428 1951
rect -8474 1879 -8468 1913
rect -8434 1879 -8428 1913
rect -8474 1864 -8428 1879
rect -8378 2849 -8332 2864
rect -8378 2815 -8372 2849
rect -8338 2815 -8332 2849
rect -8378 2777 -8332 2815
rect -8378 2743 -8372 2777
rect -8338 2743 -8332 2777
rect -8378 2705 -8332 2743
rect -8378 2671 -8372 2705
rect -8338 2671 -8332 2705
rect -8378 2633 -8332 2671
rect -8378 2599 -8372 2633
rect -8338 2599 -8332 2633
rect -8378 2561 -8332 2599
rect -8378 2527 -8372 2561
rect -8338 2527 -8332 2561
rect -8378 2489 -8332 2527
rect -8378 2455 -8372 2489
rect -8338 2455 -8332 2489
rect -8378 2417 -8332 2455
rect -8378 2383 -8372 2417
rect -8338 2383 -8332 2417
rect -8378 2345 -8332 2383
rect -8378 2311 -8372 2345
rect -8338 2311 -8332 2345
rect -8378 2273 -8332 2311
rect -8378 2239 -8372 2273
rect -8338 2239 -8332 2273
rect -8378 2201 -8332 2239
rect -8378 2167 -8372 2201
rect -8338 2167 -8332 2201
rect -8378 2129 -8332 2167
rect -8378 2095 -8372 2129
rect -8338 2095 -8332 2129
rect -8378 2057 -8332 2095
rect -8378 2023 -8372 2057
rect -8338 2023 -8332 2057
rect -8378 1985 -8332 2023
rect -8378 1951 -8372 1985
rect -8338 1951 -8332 1985
rect -8378 1913 -8332 1951
rect -8378 1879 -8372 1913
rect -8338 1879 -8332 1913
rect -8378 1864 -8332 1879
rect -8282 2849 -8236 2864
rect -8282 2815 -8276 2849
rect -8242 2815 -8236 2849
rect -8282 2777 -8236 2815
rect -8282 2743 -8276 2777
rect -8242 2743 -8236 2777
rect -8282 2705 -8236 2743
rect -8282 2671 -8276 2705
rect -8242 2671 -8236 2705
rect -8282 2633 -8236 2671
rect -8282 2599 -8276 2633
rect -8242 2599 -8236 2633
rect -8282 2561 -8236 2599
rect -8282 2527 -8276 2561
rect -8242 2527 -8236 2561
rect -8282 2489 -8236 2527
rect -8282 2455 -8276 2489
rect -8242 2455 -8236 2489
rect -8282 2417 -8236 2455
rect -8282 2383 -8276 2417
rect -8242 2383 -8236 2417
rect -8282 2345 -8236 2383
rect -8282 2311 -8276 2345
rect -8242 2311 -8236 2345
rect -8282 2273 -8236 2311
rect -8282 2239 -8276 2273
rect -8242 2239 -8236 2273
rect -8282 2201 -8236 2239
rect -8282 2167 -8276 2201
rect -8242 2167 -8236 2201
rect -8282 2129 -8236 2167
rect -8282 2095 -8276 2129
rect -8242 2095 -8236 2129
rect -8282 2057 -8236 2095
rect -8282 2023 -8276 2057
rect -8242 2023 -8236 2057
rect -8282 1985 -8236 2023
rect -8282 1951 -8276 1985
rect -8242 1951 -8236 1985
rect -8282 1913 -8236 1951
rect -8282 1879 -8276 1913
rect -8242 1879 -8236 1913
rect -8282 1864 -8236 1879
rect -8054 2841 -8008 2856
rect -8054 2807 -8048 2841
rect -8014 2807 -8008 2841
rect -8054 2769 -8008 2807
rect -8054 2735 -8048 2769
rect -8014 2735 -8008 2769
rect -8054 2697 -8008 2735
rect -8054 2663 -8048 2697
rect -8014 2663 -8008 2697
rect -8054 2625 -8008 2663
rect -8054 2591 -8048 2625
rect -8014 2591 -8008 2625
rect -8054 2553 -8008 2591
rect -8054 2519 -8048 2553
rect -8014 2519 -8008 2553
rect -8054 2481 -8008 2519
rect -8054 2447 -8048 2481
rect -8014 2447 -8008 2481
rect -8054 2409 -8008 2447
rect -8054 2375 -8048 2409
rect -8014 2375 -8008 2409
rect -8054 2337 -8008 2375
rect -8054 2303 -8048 2337
rect -8014 2303 -8008 2337
rect -8054 2265 -8008 2303
rect -8054 2231 -8048 2265
rect -8014 2231 -8008 2265
rect -8054 2193 -8008 2231
rect -8054 2159 -8048 2193
rect -8014 2159 -8008 2193
rect -8054 2121 -8008 2159
rect -8054 2087 -8048 2121
rect -8014 2087 -8008 2121
rect -8054 2049 -8008 2087
rect -8054 2015 -8048 2049
rect -8014 2015 -8008 2049
rect -8054 1977 -8008 2015
rect -8054 1943 -8048 1977
rect -8014 1943 -8008 1977
rect -8054 1905 -8008 1943
rect -8054 1871 -8048 1905
rect -8014 1871 -8008 1905
rect -8054 1856 -8008 1871
rect -7958 2841 -7912 2856
rect -7958 2807 -7952 2841
rect -7918 2807 -7912 2841
rect -7958 2769 -7912 2807
rect -7958 2735 -7952 2769
rect -7918 2735 -7912 2769
rect -7958 2697 -7912 2735
rect -7958 2663 -7952 2697
rect -7918 2663 -7912 2697
rect -7958 2625 -7912 2663
rect -7958 2591 -7952 2625
rect -7918 2591 -7912 2625
rect -7958 2553 -7912 2591
rect -7958 2519 -7952 2553
rect -7918 2519 -7912 2553
rect -7958 2481 -7912 2519
rect -7958 2447 -7952 2481
rect -7918 2447 -7912 2481
rect -7958 2409 -7912 2447
rect -7958 2375 -7952 2409
rect -7918 2375 -7912 2409
rect -7958 2337 -7912 2375
rect -7958 2303 -7952 2337
rect -7918 2303 -7912 2337
rect -7958 2265 -7912 2303
rect -7958 2231 -7952 2265
rect -7918 2231 -7912 2265
rect -7958 2193 -7912 2231
rect -7958 2159 -7952 2193
rect -7918 2159 -7912 2193
rect -7958 2121 -7912 2159
rect -7958 2087 -7952 2121
rect -7918 2087 -7912 2121
rect -7958 2049 -7912 2087
rect -7958 2015 -7952 2049
rect -7918 2015 -7912 2049
rect -7958 1977 -7912 2015
rect -7958 1943 -7952 1977
rect -7918 1943 -7912 1977
rect -7958 1905 -7912 1943
rect -7958 1871 -7952 1905
rect -7918 1871 -7912 1905
rect -7958 1856 -7912 1871
rect -7862 2841 -7816 2856
rect -7862 2807 -7856 2841
rect -7822 2807 -7816 2841
rect -7862 2769 -7816 2807
rect -7862 2735 -7856 2769
rect -7822 2735 -7816 2769
rect -7862 2697 -7816 2735
rect -7862 2663 -7856 2697
rect -7822 2663 -7816 2697
rect -7862 2625 -7816 2663
rect -7862 2591 -7856 2625
rect -7822 2591 -7816 2625
rect -7862 2553 -7816 2591
rect -7862 2519 -7856 2553
rect -7822 2519 -7816 2553
rect -7862 2481 -7816 2519
rect -7862 2447 -7856 2481
rect -7822 2447 -7816 2481
rect -7862 2409 -7816 2447
rect -7862 2375 -7856 2409
rect -7822 2375 -7816 2409
rect -7862 2337 -7816 2375
rect -7862 2303 -7856 2337
rect -7822 2303 -7816 2337
rect -7862 2265 -7816 2303
rect -7862 2231 -7856 2265
rect -7822 2231 -7816 2265
rect -7862 2193 -7816 2231
rect -7862 2159 -7856 2193
rect -7822 2159 -7816 2193
rect -7862 2121 -7816 2159
rect -7862 2087 -7856 2121
rect -7822 2087 -7816 2121
rect -7862 2049 -7816 2087
rect -7862 2015 -7856 2049
rect -7822 2015 -7816 2049
rect -7862 1977 -7816 2015
rect -7862 1943 -7856 1977
rect -7822 1943 -7816 1977
rect -7862 1905 -7816 1943
rect -7862 1871 -7856 1905
rect -7822 1871 -7816 1905
rect -7862 1856 -7816 1871
rect -7766 2841 -7720 2856
rect -7766 2807 -7760 2841
rect -7726 2807 -7720 2841
rect -7766 2769 -7720 2807
rect -7766 2735 -7760 2769
rect -7726 2735 -7720 2769
rect -7766 2697 -7720 2735
rect -7766 2663 -7760 2697
rect -7726 2663 -7720 2697
rect -7766 2625 -7720 2663
rect -7766 2591 -7760 2625
rect -7726 2591 -7720 2625
rect -7766 2553 -7720 2591
rect -7766 2519 -7760 2553
rect -7726 2519 -7720 2553
rect -7766 2481 -7720 2519
rect -7766 2447 -7760 2481
rect -7726 2447 -7720 2481
rect -7766 2409 -7720 2447
rect -7766 2375 -7760 2409
rect -7726 2375 -7720 2409
rect -7766 2337 -7720 2375
rect -7766 2303 -7760 2337
rect -7726 2303 -7720 2337
rect -7766 2265 -7720 2303
rect -7766 2231 -7760 2265
rect -7726 2231 -7720 2265
rect -7766 2193 -7720 2231
rect -7766 2159 -7760 2193
rect -7726 2159 -7720 2193
rect -7766 2121 -7720 2159
rect -7766 2087 -7760 2121
rect -7726 2087 -7720 2121
rect -7766 2049 -7720 2087
rect -7766 2015 -7760 2049
rect -7726 2015 -7720 2049
rect -7766 1977 -7720 2015
rect -7766 1943 -7760 1977
rect -7726 1943 -7720 1977
rect -7766 1905 -7720 1943
rect -7766 1871 -7760 1905
rect -7726 1871 -7720 1905
rect -7766 1856 -7720 1871
rect -7670 2841 -7624 2856
rect -7670 2807 -7664 2841
rect -7630 2807 -7624 2841
rect -7670 2769 -7624 2807
rect -7670 2735 -7664 2769
rect -7630 2735 -7624 2769
rect -7670 2697 -7624 2735
rect -7670 2663 -7664 2697
rect -7630 2663 -7624 2697
rect -7670 2625 -7624 2663
rect -7670 2591 -7664 2625
rect -7630 2591 -7624 2625
rect -7670 2553 -7624 2591
rect -7670 2519 -7664 2553
rect -7630 2519 -7624 2553
rect -7670 2481 -7624 2519
rect -7670 2447 -7664 2481
rect -7630 2447 -7624 2481
rect -7670 2409 -7624 2447
rect -7670 2375 -7664 2409
rect -7630 2375 -7624 2409
rect -7670 2337 -7624 2375
rect -7670 2303 -7664 2337
rect -7630 2303 -7624 2337
rect -7670 2265 -7624 2303
rect -7670 2231 -7664 2265
rect -7630 2231 -7624 2265
rect -7670 2193 -7624 2231
rect -7670 2159 -7664 2193
rect -7630 2159 -7624 2193
rect -7670 2121 -7624 2159
rect -7670 2087 -7664 2121
rect -7630 2087 -7624 2121
rect -7670 2049 -7624 2087
rect -7670 2015 -7664 2049
rect -7630 2015 -7624 2049
rect -7670 1977 -7624 2015
rect -7670 1943 -7664 1977
rect -7630 1943 -7624 1977
rect -7670 1905 -7624 1943
rect -7670 1871 -7664 1905
rect -7630 1871 -7624 1905
rect -7670 1856 -7624 1871
rect -7574 2841 -7528 2856
rect -7574 2807 -7568 2841
rect -7534 2807 -7528 2841
rect -7574 2769 -7528 2807
rect -7574 2735 -7568 2769
rect -7534 2735 -7528 2769
rect -7574 2697 -7528 2735
rect -7574 2663 -7568 2697
rect -7534 2663 -7528 2697
rect -7574 2625 -7528 2663
rect -7574 2591 -7568 2625
rect -7534 2591 -7528 2625
rect -7574 2553 -7528 2591
rect -7574 2519 -7568 2553
rect -7534 2519 -7528 2553
rect -7574 2481 -7528 2519
rect -7574 2447 -7568 2481
rect -7534 2447 -7528 2481
rect -7574 2409 -7528 2447
rect -7574 2375 -7568 2409
rect -7534 2375 -7528 2409
rect -7574 2337 -7528 2375
rect -7574 2303 -7568 2337
rect -7534 2303 -7528 2337
rect -7574 2265 -7528 2303
rect -7574 2231 -7568 2265
rect -7534 2231 -7528 2265
rect -7574 2193 -7528 2231
rect -7574 2159 -7568 2193
rect -7534 2159 -7528 2193
rect -7574 2121 -7528 2159
rect -7574 2087 -7568 2121
rect -7534 2087 -7528 2121
rect -7574 2049 -7528 2087
rect -7574 2015 -7568 2049
rect -7534 2015 -7528 2049
rect -7574 1977 -7528 2015
rect -7574 1943 -7568 1977
rect -7534 1943 -7528 1977
rect -7574 1905 -7528 1943
rect -7574 1871 -7568 1905
rect -7534 1871 -7528 1905
rect -7574 1856 -7528 1871
rect -7478 2841 -7432 2856
rect -7478 2807 -7472 2841
rect -7438 2807 -7432 2841
rect -7478 2769 -7432 2807
rect -7478 2735 -7472 2769
rect -7438 2735 -7432 2769
rect -7478 2697 -7432 2735
rect -7478 2663 -7472 2697
rect -7438 2663 -7432 2697
rect -7478 2625 -7432 2663
rect -7478 2591 -7472 2625
rect -7438 2591 -7432 2625
rect -7478 2553 -7432 2591
rect -7478 2519 -7472 2553
rect -7438 2519 -7432 2553
rect -7478 2481 -7432 2519
rect -7478 2447 -7472 2481
rect -7438 2447 -7432 2481
rect -7478 2409 -7432 2447
rect -7478 2375 -7472 2409
rect -7438 2375 -7432 2409
rect -7478 2337 -7432 2375
rect -7478 2303 -7472 2337
rect -7438 2303 -7432 2337
rect -7478 2265 -7432 2303
rect -7478 2231 -7472 2265
rect -7438 2231 -7432 2265
rect -7478 2193 -7432 2231
rect -7478 2159 -7472 2193
rect -7438 2159 -7432 2193
rect -7478 2121 -7432 2159
rect -7478 2087 -7472 2121
rect -7438 2087 -7432 2121
rect -7478 2049 -7432 2087
rect -7478 2015 -7472 2049
rect -7438 2015 -7432 2049
rect -7478 1977 -7432 2015
rect -7478 1943 -7472 1977
rect -7438 1943 -7432 1977
rect -7478 1905 -7432 1943
rect -7478 1871 -7472 1905
rect -7438 1871 -7432 1905
rect -7478 1856 -7432 1871
rect -7382 2841 -7336 2856
rect -7382 2807 -7376 2841
rect -7342 2807 -7336 2841
rect -7382 2769 -7336 2807
rect -7382 2735 -7376 2769
rect -7342 2735 -7336 2769
rect -7382 2697 -7336 2735
rect -7382 2663 -7376 2697
rect -7342 2663 -7336 2697
rect -7382 2625 -7336 2663
rect -7382 2591 -7376 2625
rect -7342 2591 -7336 2625
rect -7382 2553 -7336 2591
rect -7382 2519 -7376 2553
rect -7342 2519 -7336 2553
rect -7382 2481 -7336 2519
rect -7382 2447 -7376 2481
rect -7342 2447 -7336 2481
rect -7382 2409 -7336 2447
rect -7382 2375 -7376 2409
rect -7342 2375 -7336 2409
rect -7382 2337 -7336 2375
rect -7382 2303 -7376 2337
rect -7342 2303 -7336 2337
rect -7382 2265 -7336 2303
rect -7382 2231 -7376 2265
rect -7342 2231 -7336 2265
rect -7382 2193 -7336 2231
rect -7382 2159 -7376 2193
rect -7342 2159 -7336 2193
rect -7382 2121 -7336 2159
rect -7382 2087 -7376 2121
rect -7342 2087 -7336 2121
rect -7382 2049 -7336 2087
rect -7382 2015 -7376 2049
rect -7342 2015 -7336 2049
rect -7382 1977 -7336 2015
rect -7382 1943 -7376 1977
rect -7342 1943 -7336 1977
rect -7382 1905 -7336 1943
rect -7382 1871 -7376 1905
rect -7342 1871 -7336 1905
rect -7382 1856 -7336 1871
rect -7286 2841 -7240 2856
rect -7286 2807 -7280 2841
rect -7246 2807 -7240 2841
rect -7286 2769 -7240 2807
rect -7286 2735 -7280 2769
rect -7246 2735 -7240 2769
rect -7286 2697 -7240 2735
rect -7286 2663 -7280 2697
rect -7246 2663 -7240 2697
rect -7286 2625 -7240 2663
rect -7286 2591 -7280 2625
rect -7246 2591 -7240 2625
rect -7286 2553 -7240 2591
rect -7286 2519 -7280 2553
rect -7246 2519 -7240 2553
rect -7286 2481 -7240 2519
rect -7286 2447 -7280 2481
rect -7246 2447 -7240 2481
rect -7286 2409 -7240 2447
rect -7286 2375 -7280 2409
rect -7246 2375 -7240 2409
rect -7286 2337 -7240 2375
rect -7286 2303 -7280 2337
rect -7246 2303 -7240 2337
rect -7286 2265 -7240 2303
rect -7286 2231 -7280 2265
rect -7246 2231 -7240 2265
rect -7286 2193 -7240 2231
rect -7286 2159 -7280 2193
rect -7246 2159 -7240 2193
rect -7286 2121 -7240 2159
rect -7286 2087 -7280 2121
rect -7246 2087 -7240 2121
rect -7286 2049 -7240 2087
rect -7286 2015 -7280 2049
rect -7246 2015 -7240 2049
rect -7286 1977 -7240 2015
rect -7286 1943 -7280 1977
rect -7246 1943 -7240 1977
rect -7286 1905 -7240 1943
rect -7286 1871 -7280 1905
rect -7246 1871 -7240 1905
rect -7286 1856 -7240 1871
rect -7190 2841 -7144 2856
rect -7190 2807 -7184 2841
rect -7150 2807 -7144 2841
rect -7190 2769 -7144 2807
rect -7190 2735 -7184 2769
rect -7150 2735 -7144 2769
rect -7190 2697 -7144 2735
rect -7190 2663 -7184 2697
rect -7150 2663 -7144 2697
rect -7190 2625 -7144 2663
rect -7190 2591 -7184 2625
rect -7150 2591 -7144 2625
rect -7190 2553 -7144 2591
rect -7190 2519 -7184 2553
rect -7150 2519 -7144 2553
rect -7190 2481 -7144 2519
rect -7190 2447 -7184 2481
rect -7150 2447 -7144 2481
rect -7190 2409 -7144 2447
rect -7190 2375 -7184 2409
rect -7150 2375 -7144 2409
rect -7190 2337 -7144 2375
rect -7190 2303 -7184 2337
rect -7150 2303 -7144 2337
rect -7190 2265 -7144 2303
rect -7190 2231 -7184 2265
rect -7150 2231 -7144 2265
rect -7190 2193 -7144 2231
rect -7190 2159 -7184 2193
rect -7150 2159 -7144 2193
rect -7190 2121 -7144 2159
rect -7190 2087 -7184 2121
rect -7150 2087 -7144 2121
rect -7190 2049 -7144 2087
rect -7190 2015 -7184 2049
rect -7150 2015 -7144 2049
rect -7190 1977 -7144 2015
rect -7190 1943 -7184 1977
rect -7150 1943 -7144 1977
rect -7190 1905 -7144 1943
rect -7190 1871 -7184 1905
rect -7150 1871 -7144 1905
rect -7190 1856 -7144 1871
rect -7094 2841 -7048 2856
rect -7094 2807 -7088 2841
rect -7054 2807 -7048 2841
rect -7094 2769 -7048 2807
rect -7094 2735 -7088 2769
rect -7054 2735 -7048 2769
rect -7094 2697 -7048 2735
rect -7094 2663 -7088 2697
rect -7054 2663 -7048 2697
rect -7094 2625 -7048 2663
rect -7094 2591 -7088 2625
rect -7054 2591 -7048 2625
rect -7094 2553 -7048 2591
rect -7094 2519 -7088 2553
rect -7054 2519 -7048 2553
rect -7094 2481 -7048 2519
rect -7094 2447 -7088 2481
rect -7054 2447 -7048 2481
rect -7094 2409 -7048 2447
rect -7094 2375 -7088 2409
rect -7054 2375 -7048 2409
rect -7094 2337 -7048 2375
rect -7094 2303 -7088 2337
rect -7054 2303 -7048 2337
rect -7094 2265 -7048 2303
rect -7094 2231 -7088 2265
rect -7054 2231 -7048 2265
rect -7094 2193 -7048 2231
rect -7094 2159 -7088 2193
rect -7054 2159 -7048 2193
rect -7094 2121 -7048 2159
rect -7094 2087 -7088 2121
rect -7054 2087 -7048 2121
rect -7094 2049 -7048 2087
rect -7094 2015 -7088 2049
rect -7054 2015 -7048 2049
rect -7094 1977 -7048 2015
rect -7094 1943 -7088 1977
rect -7054 1943 -7048 1977
rect -7094 1905 -7048 1943
rect -7094 1871 -7088 1905
rect -7054 1871 -7048 1905
rect -7094 1856 -7048 1871
rect -6998 2841 -6952 2856
rect -6998 2807 -6992 2841
rect -6958 2807 -6952 2841
rect -6998 2769 -6952 2807
rect -6998 2735 -6992 2769
rect -6958 2735 -6952 2769
rect -6998 2697 -6952 2735
rect -6998 2663 -6992 2697
rect -6958 2663 -6952 2697
rect -6998 2625 -6952 2663
rect -6998 2591 -6992 2625
rect -6958 2591 -6952 2625
rect -6998 2553 -6952 2591
rect -6998 2519 -6992 2553
rect -6958 2519 -6952 2553
rect -6998 2481 -6952 2519
rect -6998 2447 -6992 2481
rect -6958 2447 -6952 2481
rect -6998 2409 -6952 2447
rect -6998 2375 -6992 2409
rect -6958 2375 -6952 2409
rect -6998 2337 -6952 2375
rect -6998 2303 -6992 2337
rect -6958 2303 -6952 2337
rect -6998 2265 -6952 2303
rect -6998 2231 -6992 2265
rect -6958 2231 -6952 2265
rect -6998 2193 -6952 2231
rect -6998 2159 -6992 2193
rect -6958 2159 -6952 2193
rect -6998 2121 -6952 2159
rect -6998 2087 -6992 2121
rect -6958 2087 -6952 2121
rect -6998 2049 -6952 2087
rect -6998 2015 -6992 2049
rect -6958 2015 -6952 2049
rect -6998 1977 -6952 2015
rect -6998 1943 -6992 1977
rect -6958 1943 -6952 1977
rect -6998 1905 -6952 1943
rect -6998 1871 -6992 1905
rect -6958 1871 -6952 1905
rect -6998 1856 -6952 1871
rect -6902 2841 -6856 2856
rect -6902 2807 -6896 2841
rect -6862 2807 -6856 2841
rect -6902 2769 -6856 2807
rect -6902 2735 -6896 2769
rect -6862 2735 -6856 2769
rect -6902 2697 -6856 2735
rect -6902 2663 -6896 2697
rect -6862 2663 -6856 2697
rect -6902 2625 -6856 2663
rect -6902 2591 -6896 2625
rect -6862 2591 -6856 2625
rect -6902 2553 -6856 2591
rect -6902 2519 -6896 2553
rect -6862 2519 -6856 2553
rect -6902 2481 -6856 2519
rect -6902 2447 -6896 2481
rect -6862 2447 -6856 2481
rect -6902 2409 -6856 2447
rect -6902 2375 -6896 2409
rect -6862 2375 -6856 2409
rect -6902 2337 -6856 2375
rect -6902 2303 -6896 2337
rect -6862 2303 -6856 2337
rect -6902 2265 -6856 2303
rect -6902 2231 -6896 2265
rect -6862 2231 -6856 2265
rect -6902 2193 -6856 2231
rect -6902 2159 -6896 2193
rect -6862 2159 -6856 2193
rect -6902 2121 -6856 2159
rect -6902 2087 -6896 2121
rect -6862 2087 -6856 2121
rect -6902 2049 -6856 2087
rect -6902 2015 -6896 2049
rect -6862 2015 -6856 2049
rect -6902 1977 -6856 2015
rect -6902 1943 -6896 1977
rect -6862 1943 -6856 1977
rect -6902 1905 -6856 1943
rect -6902 1871 -6896 1905
rect -6862 1871 -6856 1905
rect -6902 1856 -6856 1871
rect -6806 2841 -6760 2856
rect -6806 2807 -6800 2841
rect -6766 2807 -6760 2841
rect -6806 2769 -6760 2807
rect -6806 2735 -6800 2769
rect -6766 2735 -6760 2769
rect -6806 2697 -6760 2735
rect -6806 2663 -6800 2697
rect -6766 2663 -6760 2697
rect -6806 2625 -6760 2663
rect -6806 2591 -6800 2625
rect -6766 2591 -6760 2625
rect -6806 2553 -6760 2591
rect -6806 2519 -6800 2553
rect -6766 2519 -6760 2553
rect -6806 2481 -6760 2519
rect -6806 2447 -6800 2481
rect -6766 2447 -6760 2481
rect -6806 2409 -6760 2447
rect -6806 2375 -6800 2409
rect -6766 2375 -6760 2409
rect -6806 2337 -6760 2375
rect -6806 2303 -6800 2337
rect -6766 2303 -6760 2337
rect -6806 2265 -6760 2303
rect -6806 2231 -6800 2265
rect -6766 2231 -6760 2265
rect -6806 2193 -6760 2231
rect -6806 2159 -6800 2193
rect -6766 2159 -6760 2193
rect -6806 2121 -6760 2159
rect -6806 2087 -6800 2121
rect -6766 2087 -6760 2121
rect -6806 2049 -6760 2087
rect -6806 2015 -6800 2049
rect -6766 2015 -6760 2049
rect -6806 1977 -6760 2015
rect -6806 1943 -6800 1977
rect -6766 1943 -6760 1977
rect -6806 1905 -6760 1943
rect -6806 1871 -6800 1905
rect -6766 1871 -6760 1905
rect -6806 1856 -6760 1871
rect -6710 2841 -6664 2856
rect -6710 2807 -6704 2841
rect -6670 2807 -6664 2841
rect -6710 2769 -6664 2807
rect -6710 2735 -6704 2769
rect -6670 2735 -6664 2769
rect -6710 2697 -6664 2735
rect -6710 2663 -6704 2697
rect -6670 2663 -6664 2697
rect -6710 2625 -6664 2663
rect -6710 2591 -6704 2625
rect -6670 2591 -6664 2625
rect -6710 2553 -6664 2591
rect -6710 2519 -6704 2553
rect -6670 2519 -6664 2553
rect -6710 2481 -6664 2519
rect -6710 2447 -6704 2481
rect -6670 2447 -6664 2481
rect -6710 2409 -6664 2447
rect -6710 2375 -6704 2409
rect -6670 2375 -6664 2409
rect -6710 2337 -6664 2375
rect -6710 2303 -6704 2337
rect -6670 2303 -6664 2337
rect -6710 2265 -6664 2303
rect -6710 2231 -6704 2265
rect -6670 2231 -6664 2265
rect -6710 2193 -6664 2231
rect -6710 2159 -6704 2193
rect -6670 2159 -6664 2193
rect -6710 2121 -6664 2159
rect -6710 2087 -6704 2121
rect -6670 2087 -6664 2121
rect -6710 2049 -6664 2087
rect -6710 2015 -6704 2049
rect -6670 2015 -6664 2049
rect -6710 1977 -6664 2015
rect -6710 1943 -6704 1977
rect -6670 1943 -6664 1977
rect -6710 1905 -6664 1943
rect -6710 1871 -6704 1905
rect -6670 1871 -6664 1905
rect -6710 1856 -6664 1871
rect -6614 2841 -6568 2856
rect -6614 2807 -6608 2841
rect -6574 2807 -6568 2841
rect -6614 2769 -6568 2807
rect -6614 2735 -6608 2769
rect -6574 2735 -6568 2769
rect -6614 2697 -6568 2735
rect -6614 2663 -6608 2697
rect -6574 2663 -6568 2697
rect -6614 2625 -6568 2663
rect -6614 2591 -6608 2625
rect -6574 2591 -6568 2625
rect -6614 2553 -6568 2591
rect -6614 2519 -6608 2553
rect -6574 2519 -6568 2553
rect -6614 2481 -6568 2519
rect -6614 2447 -6608 2481
rect -6574 2447 -6568 2481
rect -6614 2409 -6568 2447
rect -6614 2375 -6608 2409
rect -6574 2375 -6568 2409
rect -6614 2337 -6568 2375
rect -6614 2303 -6608 2337
rect -6574 2303 -6568 2337
rect -6614 2265 -6568 2303
rect -6614 2231 -6608 2265
rect -6574 2231 -6568 2265
rect -6614 2193 -6568 2231
rect -6614 2159 -6608 2193
rect -6574 2159 -6568 2193
rect -6614 2121 -6568 2159
rect -6614 2087 -6608 2121
rect -6574 2087 -6568 2121
rect -6614 2049 -6568 2087
rect -6614 2015 -6608 2049
rect -6574 2015 -6568 2049
rect -6614 1977 -6568 2015
rect -6614 1943 -6608 1977
rect -6574 1943 -6568 1977
rect -6614 1905 -6568 1943
rect -6614 1871 -6608 1905
rect -6574 1871 -6568 1905
rect -6614 1856 -6568 1871
rect -6376 2845 -6330 2860
rect -6376 2811 -6370 2845
rect -6336 2811 -6330 2845
rect -6376 2773 -6330 2811
rect -6376 2739 -6370 2773
rect -6336 2739 -6330 2773
rect -6376 2701 -6330 2739
rect -6376 2667 -6370 2701
rect -6336 2667 -6330 2701
rect -6376 2629 -6330 2667
rect -6376 2595 -6370 2629
rect -6336 2595 -6330 2629
rect -6376 2557 -6330 2595
rect -6376 2523 -6370 2557
rect -6336 2523 -6330 2557
rect -6376 2485 -6330 2523
rect -6376 2451 -6370 2485
rect -6336 2451 -6330 2485
rect -6376 2413 -6330 2451
rect -6376 2379 -6370 2413
rect -6336 2379 -6330 2413
rect -6376 2341 -6330 2379
rect -6376 2307 -6370 2341
rect -6336 2307 -6330 2341
rect -6376 2269 -6330 2307
rect -6376 2235 -6370 2269
rect -6336 2235 -6330 2269
rect -6376 2197 -6330 2235
rect -6376 2163 -6370 2197
rect -6336 2163 -6330 2197
rect -6376 2125 -6330 2163
rect -6376 2091 -6370 2125
rect -6336 2091 -6330 2125
rect -6376 2053 -6330 2091
rect -6376 2019 -6370 2053
rect -6336 2019 -6330 2053
rect -6376 1981 -6330 2019
rect -6376 1947 -6370 1981
rect -6336 1947 -6330 1981
rect -6376 1909 -6330 1947
rect -6376 1875 -6370 1909
rect -6336 1875 -6330 1909
rect -6376 1860 -6330 1875
rect -6280 2845 -6234 2860
rect -6280 2811 -6274 2845
rect -6240 2811 -6234 2845
rect -6280 2773 -6234 2811
rect -6280 2739 -6274 2773
rect -6240 2739 -6234 2773
rect -6280 2701 -6234 2739
rect -6280 2667 -6274 2701
rect -6240 2667 -6234 2701
rect -6280 2629 -6234 2667
rect -6280 2595 -6274 2629
rect -6240 2595 -6234 2629
rect -6280 2557 -6234 2595
rect -6280 2523 -6274 2557
rect -6240 2523 -6234 2557
rect -6280 2485 -6234 2523
rect -6280 2451 -6274 2485
rect -6240 2451 -6234 2485
rect -6280 2413 -6234 2451
rect -6280 2379 -6274 2413
rect -6240 2379 -6234 2413
rect -6280 2341 -6234 2379
rect -6280 2307 -6274 2341
rect -6240 2307 -6234 2341
rect -6280 2269 -6234 2307
rect -6280 2235 -6274 2269
rect -6240 2235 -6234 2269
rect -6280 2197 -6234 2235
rect -6280 2163 -6274 2197
rect -6240 2163 -6234 2197
rect -6280 2125 -6234 2163
rect -6280 2091 -6274 2125
rect -6240 2091 -6234 2125
rect -6280 2053 -6234 2091
rect -6280 2019 -6274 2053
rect -6240 2019 -6234 2053
rect -6280 1981 -6234 2019
rect -6280 1947 -6274 1981
rect -6240 1947 -6234 1981
rect -6280 1909 -6234 1947
rect -6280 1875 -6274 1909
rect -6240 1875 -6234 1909
rect -6280 1860 -6234 1875
rect -6184 2845 -6138 2860
rect -6184 2811 -6178 2845
rect -6144 2811 -6138 2845
rect -6184 2773 -6138 2811
rect -6184 2739 -6178 2773
rect -6144 2739 -6138 2773
rect -6184 2701 -6138 2739
rect -6184 2667 -6178 2701
rect -6144 2667 -6138 2701
rect -6184 2629 -6138 2667
rect -6184 2595 -6178 2629
rect -6144 2595 -6138 2629
rect -6184 2557 -6138 2595
rect -6184 2523 -6178 2557
rect -6144 2523 -6138 2557
rect -6184 2485 -6138 2523
rect -6184 2451 -6178 2485
rect -6144 2451 -6138 2485
rect -6184 2413 -6138 2451
rect -6184 2379 -6178 2413
rect -6144 2379 -6138 2413
rect -6184 2341 -6138 2379
rect -6184 2307 -6178 2341
rect -6144 2307 -6138 2341
rect -6184 2269 -6138 2307
rect -6184 2235 -6178 2269
rect -6144 2235 -6138 2269
rect -6184 2197 -6138 2235
rect -6184 2163 -6178 2197
rect -6144 2163 -6138 2197
rect -6184 2125 -6138 2163
rect -6184 2091 -6178 2125
rect -6144 2091 -6138 2125
rect -6184 2053 -6138 2091
rect -6184 2019 -6178 2053
rect -6144 2019 -6138 2053
rect -6184 1981 -6138 2019
rect -6184 1947 -6178 1981
rect -6144 1947 -6138 1981
rect -6184 1909 -6138 1947
rect -6184 1875 -6178 1909
rect -6144 1875 -6138 1909
rect -6184 1860 -6138 1875
rect -6088 2845 -6042 2860
rect -6088 2811 -6082 2845
rect -6048 2811 -6042 2845
rect -6088 2773 -6042 2811
rect -6088 2739 -6082 2773
rect -6048 2739 -6042 2773
rect -6088 2701 -6042 2739
rect -6088 2667 -6082 2701
rect -6048 2667 -6042 2701
rect -6088 2629 -6042 2667
rect -6088 2595 -6082 2629
rect -6048 2595 -6042 2629
rect -6088 2557 -6042 2595
rect -6088 2523 -6082 2557
rect -6048 2523 -6042 2557
rect -6088 2485 -6042 2523
rect -6088 2451 -6082 2485
rect -6048 2451 -6042 2485
rect -6088 2413 -6042 2451
rect -6088 2379 -6082 2413
rect -6048 2379 -6042 2413
rect -6088 2341 -6042 2379
rect -6088 2307 -6082 2341
rect -6048 2307 -6042 2341
rect -6088 2269 -6042 2307
rect -6088 2235 -6082 2269
rect -6048 2235 -6042 2269
rect -6088 2197 -6042 2235
rect -6088 2163 -6082 2197
rect -6048 2163 -6042 2197
rect -6088 2125 -6042 2163
rect -6088 2091 -6082 2125
rect -6048 2091 -6042 2125
rect -6088 2053 -6042 2091
rect -6088 2019 -6082 2053
rect -6048 2019 -6042 2053
rect -6088 1981 -6042 2019
rect -6088 1947 -6082 1981
rect -6048 1947 -6042 1981
rect -6088 1909 -6042 1947
rect -6088 1875 -6082 1909
rect -6048 1875 -6042 1909
rect -6088 1860 -6042 1875
rect -5992 2845 -5946 2860
rect -5992 2811 -5986 2845
rect -5952 2811 -5946 2845
rect -5992 2773 -5946 2811
rect -5992 2739 -5986 2773
rect -5952 2739 -5946 2773
rect -5992 2701 -5946 2739
rect -5992 2667 -5986 2701
rect -5952 2667 -5946 2701
rect -5992 2629 -5946 2667
rect -5992 2595 -5986 2629
rect -5952 2595 -5946 2629
rect -5992 2557 -5946 2595
rect -5992 2523 -5986 2557
rect -5952 2523 -5946 2557
rect -5992 2485 -5946 2523
rect -5992 2451 -5986 2485
rect -5952 2451 -5946 2485
rect -5992 2413 -5946 2451
rect -5992 2379 -5986 2413
rect -5952 2379 -5946 2413
rect -5992 2341 -5946 2379
rect -5992 2307 -5986 2341
rect -5952 2307 -5946 2341
rect -5992 2269 -5946 2307
rect -5992 2235 -5986 2269
rect -5952 2235 -5946 2269
rect -5992 2197 -5946 2235
rect -5992 2163 -5986 2197
rect -5952 2163 -5946 2197
rect -5992 2125 -5946 2163
rect -5992 2091 -5986 2125
rect -5952 2091 -5946 2125
rect -5992 2053 -5946 2091
rect -5992 2019 -5986 2053
rect -5952 2019 -5946 2053
rect -5992 1981 -5946 2019
rect -5992 1947 -5986 1981
rect -5952 1947 -5946 1981
rect -5992 1909 -5946 1947
rect -5992 1875 -5986 1909
rect -5952 1875 -5946 1909
rect -5992 1860 -5946 1875
rect -5896 2845 -5850 2860
rect -5896 2811 -5890 2845
rect -5856 2811 -5850 2845
rect -5896 2773 -5850 2811
rect -5896 2739 -5890 2773
rect -5856 2739 -5850 2773
rect -5896 2701 -5850 2739
rect -5896 2667 -5890 2701
rect -5856 2667 -5850 2701
rect -5896 2629 -5850 2667
rect -5896 2595 -5890 2629
rect -5856 2595 -5850 2629
rect -5896 2557 -5850 2595
rect -5896 2523 -5890 2557
rect -5856 2523 -5850 2557
rect -5896 2485 -5850 2523
rect -5896 2451 -5890 2485
rect -5856 2451 -5850 2485
rect -5896 2413 -5850 2451
rect -5896 2379 -5890 2413
rect -5856 2379 -5850 2413
rect -5896 2341 -5850 2379
rect -5896 2307 -5890 2341
rect -5856 2307 -5850 2341
rect -5896 2269 -5850 2307
rect -5896 2235 -5890 2269
rect -5856 2235 -5850 2269
rect -5896 2197 -5850 2235
rect -5896 2163 -5890 2197
rect -5856 2163 -5850 2197
rect -5896 2125 -5850 2163
rect -5896 2091 -5890 2125
rect -5856 2091 -5850 2125
rect -5896 2053 -5850 2091
rect -5896 2019 -5890 2053
rect -5856 2019 -5850 2053
rect -5896 1981 -5850 2019
rect -5896 1947 -5890 1981
rect -5856 1947 -5850 1981
rect -5896 1909 -5850 1947
rect -5896 1875 -5890 1909
rect -5856 1875 -5850 1909
rect -5896 1860 -5850 1875
rect -5800 2845 -5754 2860
rect -5800 2811 -5794 2845
rect -5760 2811 -5754 2845
rect -5800 2773 -5754 2811
rect -5800 2739 -5794 2773
rect -5760 2739 -5754 2773
rect -5800 2701 -5754 2739
rect -5800 2667 -5794 2701
rect -5760 2667 -5754 2701
rect -5800 2629 -5754 2667
rect -5800 2595 -5794 2629
rect -5760 2595 -5754 2629
rect -5800 2557 -5754 2595
rect -5800 2523 -5794 2557
rect -5760 2523 -5754 2557
rect -5800 2485 -5754 2523
rect -5800 2451 -5794 2485
rect -5760 2451 -5754 2485
rect -5800 2413 -5754 2451
rect -5800 2379 -5794 2413
rect -5760 2379 -5754 2413
rect -5800 2341 -5754 2379
rect -5800 2307 -5794 2341
rect -5760 2307 -5754 2341
rect -5800 2269 -5754 2307
rect -5800 2235 -5794 2269
rect -5760 2235 -5754 2269
rect -5800 2197 -5754 2235
rect -5800 2163 -5794 2197
rect -5760 2163 -5754 2197
rect -5800 2125 -5754 2163
rect -5800 2091 -5794 2125
rect -5760 2091 -5754 2125
rect -5800 2053 -5754 2091
rect -5800 2019 -5794 2053
rect -5760 2019 -5754 2053
rect -5800 1981 -5754 2019
rect -5800 1947 -5794 1981
rect -5760 1947 -5754 1981
rect -5800 1909 -5754 1947
rect -5800 1875 -5794 1909
rect -5760 1875 -5754 1909
rect -5800 1860 -5754 1875
rect -5704 2845 -5658 2860
rect -5704 2811 -5698 2845
rect -5664 2811 -5658 2845
rect -5704 2773 -5658 2811
rect -5704 2739 -5698 2773
rect -5664 2739 -5658 2773
rect -5704 2701 -5658 2739
rect -5704 2667 -5698 2701
rect -5664 2667 -5658 2701
rect -5704 2629 -5658 2667
rect -5704 2595 -5698 2629
rect -5664 2595 -5658 2629
rect -5704 2557 -5658 2595
rect -5704 2523 -5698 2557
rect -5664 2523 -5658 2557
rect -5704 2485 -5658 2523
rect -5704 2451 -5698 2485
rect -5664 2451 -5658 2485
rect -5704 2413 -5658 2451
rect -5704 2379 -5698 2413
rect -5664 2379 -5658 2413
rect -5704 2341 -5658 2379
rect -5704 2307 -5698 2341
rect -5664 2307 -5658 2341
rect -5704 2269 -5658 2307
rect -5704 2235 -5698 2269
rect -5664 2235 -5658 2269
rect -5704 2197 -5658 2235
rect -5704 2163 -5698 2197
rect -5664 2163 -5658 2197
rect -5704 2125 -5658 2163
rect -5704 2091 -5698 2125
rect -5664 2091 -5658 2125
rect -5704 2053 -5658 2091
rect -5704 2019 -5698 2053
rect -5664 2019 -5658 2053
rect -5704 1981 -5658 2019
rect -5704 1947 -5698 1981
rect -5664 1947 -5658 1981
rect -5704 1909 -5658 1947
rect -5704 1875 -5698 1909
rect -5664 1875 -5658 1909
rect -5704 1860 -5658 1875
rect -5608 2845 -5562 2860
rect -5608 2811 -5602 2845
rect -5568 2811 -5562 2845
rect -5608 2773 -5562 2811
rect -5608 2739 -5602 2773
rect -5568 2739 -5562 2773
rect -5608 2701 -5562 2739
rect -5608 2667 -5602 2701
rect -5568 2667 -5562 2701
rect -5608 2629 -5562 2667
rect -5608 2595 -5602 2629
rect -5568 2595 -5562 2629
rect -5608 2557 -5562 2595
rect -5608 2523 -5602 2557
rect -5568 2523 -5562 2557
rect -5608 2485 -5562 2523
rect -5608 2451 -5602 2485
rect -5568 2451 -5562 2485
rect -5608 2413 -5562 2451
rect -5608 2379 -5602 2413
rect -5568 2379 -5562 2413
rect -5608 2341 -5562 2379
rect -5608 2307 -5602 2341
rect -5568 2307 -5562 2341
rect -5608 2269 -5562 2307
rect -5608 2235 -5602 2269
rect -5568 2235 -5562 2269
rect -5608 2197 -5562 2235
rect -5608 2163 -5602 2197
rect -5568 2163 -5562 2197
rect -5608 2125 -5562 2163
rect -5608 2091 -5602 2125
rect -5568 2091 -5562 2125
rect -5608 2053 -5562 2091
rect -5608 2019 -5602 2053
rect -5568 2019 -5562 2053
rect -5608 1981 -5562 2019
rect -5608 1947 -5602 1981
rect -5568 1947 -5562 1981
rect -5608 1909 -5562 1947
rect -5608 1875 -5602 1909
rect -5568 1875 -5562 1909
rect -5608 1860 -5562 1875
rect -5512 2845 -5466 2860
rect -5512 2811 -5506 2845
rect -5472 2811 -5466 2845
rect -5512 2773 -5466 2811
rect -5512 2739 -5506 2773
rect -5472 2739 -5466 2773
rect -5512 2701 -5466 2739
rect -5512 2667 -5506 2701
rect -5472 2667 -5466 2701
rect -5512 2629 -5466 2667
rect -5512 2595 -5506 2629
rect -5472 2595 -5466 2629
rect -5512 2557 -5466 2595
rect -5512 2523 -5506 2557
rect -5472 2523 -5466 2557
rect -5512 2485 -5466 2523
rect -5512 2451 -5506 2485
rect -5472 2451 -5466 2485
rect -5512 2413 -5466 2451
rect -5512 2379 -5506 2413
rect -5472 2379 -5466 2413
rect -5512 2341 -5466 2379
rect -5512 2307 -5506 2341
rect -5472 2307 -5466 2341
rect -5512 2269 -5466 2307
rect -5512 2235 -5506 2269
rect -5472 2235 -5466 2269
rect -5512 2197 -5466 2235
rect -5512 2163 -5506 2197
rect -5472 2163 -5466 2197
rect -5512 2125 -5466 2163
rect -5512 2091 -5506 2125
rect -5472 2091 -5466 2125
rect -5512 2053 -5466 2091
rect -5512 2019 -5506 2053
rect -5472 2019 -5466 2053
rect -5512 1981 -5466 2019
rect -5512 1947 -5506 1981
rect -5472 1947 -5466 1981
rect -5512 1909 -5466 1947
rect -5512 1875 -5506 1909
rect -5472 1875 -5466 1909
rect -5512 1860 -5466 1875
rect -5416 2845 -5370 2860
rect -5416 2811 -5410 2845
rect -5376 2811 -5370 2845
rect -5416 2773 -5370 2811
rect -5416 2739 -5410 2773
rect -5376 2739 -5370 2773
rect -5416 2701 -5370 2739
rect -5416 2667 -5410 2701
rect -5376 2667 -5370 2701
rect -5416 2629 -5370 2667
rect -5416 2595 -5410 2629
rect -5376 2595 -5370 2629
rect -5416 2557 -5370 2595
rect -5416 2523 -5410 2557
rect -5376 2523 -5370 2557
rect -5416 2485 -5370 2523
rect -5416 2451 -5410 2485
rect -5376 2451 -5370 2485
rect -5416 2413 -5370 2451
rect -5416 2379 -5410 2413
rect -5376 2379 -5370 2413
rect -5416 2341 -5370 2379
rect -5416 2307 -5410 2341
rect -5376 2307 -5370 2341
rect -5416 2269 -5370 2307
rect -5416 2235 -5410 2269
rect -5376 2235 -5370 2269
rect -5416 2197 -5370 2235
rect -5416 2163 -5410 2197
rect -5376 2163 -5370 2197
rect -5416 2125 -5370 2163
rect -5416 2091 -5410 2125
rect -5376 2091 -5370 2125
rect -5416 2053 -5370 2091
rect -5416 2019 -5410 2053
rect -5376 2019 -5370 2053
rect -5416 1981 -5370 2019
rect -5416 1947 -5410 1981
rect -5376 1947 -5370 1981
rect -5416 1909 -5370 1947
rect -5416 1875 -5410 1909
rect -5376 1875 -5370 1909
rect -5416 1860 -5370 1875
rect -5204 2855 -5158 2870
rect -5204 2821 -5198 2855
rect -5164 2821 -5158 2855
rect -5204 2783 -5158 2821
rect -5204 2749 -5198 2783
rect -5164 2749 -5158 2783
rect -5204 2711 -5158 2749
rect -5204 2677 -5198 2711
rect -5164 2677 -5158 2711
rect -5204 2639 -5158 2677
rect -5204 2605 -5198 2639
rect -5164 2605 -5158 2639
rect -5204 2567 -5158 2605
rect -5204 2533 -5198 2567
rect -5164 2533 -5158 2567
rect -5204 2495 -5158 2533
rect -5204 2461 -5198 2495
rect -5164 2461 -5158 2495
rect -5204 2423 -5158 2461
rect -5204 2389 -5198 2423
rect -5164 2389 -5158 2423
rect -5204 2351 -5158 2389
rect -5204 2317 -5198 2351
rect -5164 2317 -5158 2351
rect -5204 2279 -5158 2317
rect -5204 2245 -5198 2279
rect -5164 2245 -5158 2279
rect -5204 2207 -5158 2245
rect -5204 2173 -5198 2207
rect -5164 2173 -5158 2207
rect -5204 2135 -5158 2173
rect -5204 2101 -5198 2135
rect -5164 2101 -5158 2135
rect -5204 2063 -5158 2101
rect -5204 2029 -5198 2063
rect -5164 2029 -5158 2063
rect -5204 1991 -5158 2029
rect -5204 1957 -5198 1991
rect -5164 1957 -5158 1991
rect -5204 1919 -5158 1957
rect -5204 1885 -5198 1919
rect -5164 1885 -5158 1919
rect -5204 1870 -5158 1885
rect -5108 2855 -5062 2870
rect -5108 2821 -5102 2855
rect -5068 2821 -5062 2855
rect -5108 2783 -5062 2821
rect -5108 2749 -5102 2783
rect -5068 2749 -5062 2783
rect -5108 2711 -5062 2749
rect -5108 2677 -5102 2711
rect -5068 2677 -5062 2711
rect -5108 2639 -5062 2677
rect -5108 2605 -5102 2639
rect -5068 2605 -5062 2639
rect -5108 2567 -5062 2605
rect -5108 2533 -5102 2567
rect -5068 2533 -5062 2567
rect -5108 2495 -5062 2533
rect -5108 2461 -5102 2495
rect -5068 2461 -5062 2495
rect -5108 2423 -5062 2461
rect -5108 2389 -5102 2423
rect -5068 2389 -5062 2423
rect -5108 2351 -5062 2389
rect -5108 2317 -5102 2351
rect -5068 2317 -5062 2351
rect -5108 2279 -5062 2317
rect -5108 2245 -5102 2279
rect -5068 2245 -5062 2279
rect -5108 2207 -5062 2245
rect -5108 2173 -5102 2207
rect -5068 2173 -5062 2207
rect -5108 2135 -5062 2173
rect -5108 2101 -5102 2135
rect -5068 2101 -5062 2135
rect -5108 2063 -5062 2101
rect -5108 2029 -5102 2063
rect -5068 2029 -5062 2063
rect -5108 1991 -5062 2029
rect -5108 1957 -5102 1991
rect -5068 1957 -5062 1991
rect -5108 1919 -5062 1957
rect -5108 1885 -5102 1919
rect -5068 1885 -5062 1919
rect -5108 1870 -5062 1885
rect -5012 2855 -4966 2870
rect -5012 2821 -5006 2855
rect -4972 2821 -4966 2855
rect -5012 2783 -4966 2821
rect -5012 2749 -5006 2783
rect -4972 2749 -4966 2783
rect -5012 2711 -4966 2749
rect -5012 2677 -5006 2711
rect -4972 2677 -4966 2711
rect -5012 2639 -4966 2677
rect -5012 2605 -5006 2639
rect -4972 2605 -4966 2639
rect -5012 2567 -4966 2605
rect -5012 2533 -5006 2567
rect -4972 2533 -4966 2567
rect -5012 2495 -4966 2533
rect -5012 2461 -5006 2495
rect -4972 2461 -4966 2495
rect -5012 2423 -4966 2461
rect -5012 2389 -5006 2423
rect -4972 2389 -4966 2423
rect -5012 2351 -4966 2389
rect -5012 2317 -5006 2351
rect -4972 2317 -4966 2351
rect -5012 2279 -4966 2317
rect -5012 2245 -5006 2279
rect -4972 2245 -4966 2279
rect -5012 2207 -4966 2245
rect -5012 2173 -5006 2207
rect -4972 2173 -4966 2207
rect -5012 2135 -4966 2173
rect -5012 2101 -5006 2135
rect -4972 2101 -4966 2135
rect -5012 2063 -4966 2101
rect -5012 2029 -5006 2063
rect -4972 2029 -4966 2063
rect -5012 1991 -4966 2029
rect -5012 1957 -5006 1991
rect -4972 1957 -4966 1991
rect -5012 1919 -4966 1957
rect -5012 1885 -5006 1919
rect -4972 1885 -4966 1919
rect -5012 1870 -4966 1885
rect -4916 2855 -4870 2870
rect -4916 2821 -4910 2855
rect -4876 2821 -4870 2855
rect -4916 2783 -4870 2821
rect -4916 2749 -4910 2783
rect -4876 2749 -4870 2783
rect -4916 2711 -4870 2749
rect -4916 2677 -4910 2711
rect -4876 2677 -4870 2711
rect -4916 2639 -4870 2677
rect -4916 2605 -4910 2639
rect -4876 2605 -4870 2639
rect -4916 2567 -4870 2605
rect -4916 2533 -4910 2567
rect -4876 2533 -4870 2567
rect -4916 2495 -4870 2533
rect -4916 2461 -4910 2495
rect -4876 2461 -4870 2495
rect -4916 2423 -4870 2461
rect -4916 2389 -4910 2423
rect -4876 2389 -4870 2423
rect -4916 2351 -4870 2389
rect -4916 2317 -4910 2351
rect -4876 2317 -4870 2351
rect -4916 2279 -4870 2317
rect -4916 2245 -4910 2279
rect -4876 2245 -4870 2279
rect -4916 2207 -4870 2245
rect -4916 2173 -4910 2207
rect -4876 2173 -4870 2207
rect -4916 2135 -4870 2173
rect -4916 2101 -4910 2135
rect -4876 2101 -4870 2135
rect -4916 2063 -4870 2101
rect -4916 2029 -4910 2063
rect -4876 2029 -4870 2063
rect -4916 1991 -4870 2029
rect -4916 1957 -4910 1991
rect -4876 1957 -4870 1991
rect -4916 1919 -4870 1957
rect -4916 1885 -4910 1919
rect -4876 1885 -4870 1919
rect -4916 1870 -4870 1885
rect -4820 2855 -4774 2870
rect -4820 2821 -4814 2855
rect -4780 2821 -4774 2855
rect -4820 2783 -4774 2821
rect -4820 2749 -4814 2783
rect -4780 2749 -4774 2783
rect -4820 2711 -4774 2749
rect -4820 2677 -4814 2711
rect -4780 2677 -4774 2711
rect -4820 2639 -4774 2677
rect -4820 2605 -4814 2639
rect -4780 2605 -4774 2639
rect -4820 2567 -4774 2605
rect -4820 2533 -4814 2567
rect -4780 2533 -4774 2567
rect -4820 2495 -4774 2533
rect -4820 2461 -4814 2495
rect -4780 2461 -4774 2495
rect -4820 2423 -4774 2461
rect -4820 2389 -4814 2423
rect -4780 2389 -4774 2423
rect -4820 2351 -4774 2389
rect -4820 2317 -4814 2351
rect -4780 2317 -4774 2351
rect -4820 2279 -4774 2317
rect -4820 2245 -4814 2279
rect -4780 2245 -4774 2279
rect -4820 2207 -4774 2245
rect -4820 2173 -4814 2207
rect -4780 2173 -4774 2207
rect -4820 2135 -4774 2173
rect -4820 2101 -4814 2135
rect -4780 2101 -4774 2135
rect -4820 2063 -4774 2101
rect -4820 2029 -4814 2063
rect -4780 2029 -4774 2063
rect -4820 1991 -4774 2029
rect -4820 1957 -4814 1991
rect -4780 1957 -4774 1991
rect -4820 1919 -4774 1957
rect -4820 1885 -4814 1919
rect -4780 1885 -4774 1919
rect -4820 1870 -4774 1885
rect -4724 2855 -4678 2870
rect -4724 2821 -4718 2855
rect -4684 2821 -4678 2855
rect -4724 2783 -4678 2821
rect -4724 2749 -4718 2783
rect -4684 2749 -4678 2783
rect -4724 2711 -4678 2749
rect -4724 2677 -4718 2711
rect -4684 2677 -4678 2711
rect -4724 2639 -4678 2677
rect -4724 2605 -4718 2639
rect -4684 2605 -4678 2639
rect -4724 2567 -4678 2605
rect -4724 2533 -4718 2567
rect -4684 2533 -4678 2567
rect -4724 2495 -4678 2533
rect -2406 2506 -2396 2668
rect -2244 2624 -2234 2668
rect -1932 2624 -1864 3372
rect -1126 3324 -1020 4630
rect 1478 4607 1484 4641
rect 1518 4607 1524 4641
rect 1478 4569 1524 4607
rect 1478 4535 1484 4569
rect 1518 4535 1524 4569
rect 1478 4497 1524 4535
rect 1478 4463 1484 4497
rect 1518 4463 1524 4497
rect 1478 4425 1524 4463
rect 1478 4391 1484 4425
rect 1518 4391 1524 4425
rect 1478 4353 1524 4391
rect 1478 4319 1484 4353
rect 1518 4319 1524 4353
rect 1478 4281 1524 4319
rect 1478 4247 1484 4281
rect 1518 4247 1524 4281
rect 1478 4209 1524 4247
rect 1478 4175 1484 4209
rect 1518 4175 1524 4209
rect 1478 4137 1524 4175
rect 1478 4103 1484 4137
rect 1518 4103 1524 4137
rect 1478 4065 1524 4103
rect 1478 4031 1484 4065
rect 1518 4031 1524 4065
rect 1478 3993 1524 4031
rect 1478 3959 1484 3993
rect 1518 3959 1524 3993
rect 1478 3944 1524 3959
rect 1574 4929 1620 4944
rect 1574 4895 1580 4929
rect 1614 4895 1620 4929
rect 1574 4857 1620 4895
rect 1574 4823 1580 4857
rect 1614 4823 1620 4857
rect 1574 4785 1620 4823
rect 1574 4751 1580 4785
rect 1614 4751 1620 4785
rect 1574 4713 1620 4751
rect 1574 4679 1580 4713
rect 1614 4679 1620 4713
rect 1574 4641 1620 4679
rect 1574 4607 1580 4641
rect 1614 4607 1620 4641
rect 1574 4569 1620 4607
rect 1574 4535 1580 4569
rect 1614 4535 1620 4569
rect 1574 4497 1620 4535
rect 1574 4463 1580 4497
rect 1614 4463 1620 4497
rect 1574 4425 1620 4463
rect 1574 4391 1580 4425
rect 1614 4391 1620 4425
rect 1574 4353 1620 4391
rect 1574 4319 1580 4353
rect 1614 4319 1620 4353
rect 1574 4281 1620 4319
rect 1574 4247 1580 4281
rect 1614 4247 1620 4281
rect 1574 4209 1620 4247
rect 1574 4175 1580 4209
rect 1614 4175 1620 4209
rect 1574 4137 1620 4175
rect 1574 4103 1580 4137
rect 1614 4103 1620 4137
rect 1574 4065 1620 4103
rect 1574 4031 1580 4065
rect 1614 4031 1620 4065
rect 1574 3993 1620 4031
rect 1574 3959 1580 3993
rect 1614 3959 1620 3993
rect 1574 3944 1620 3959
rect 1670 4929 1716 4944
rect 1670 4895 1676 4929
rect 1710 4895 1716 4929
rect 1670 4857 1716 4895
rect 1670 4823 1676 4857
rect 1710 4823 1716 4857
rect 1670 4785 1716 4823
rect 1670 4751 1676 4785
rect 1710 4751 1716 4785
rect 1670 4713 1716 4751
rect 1670 4679 1676 4713
rect 1710 4679 1716 4713
rect 1670 4641 1716 4679
rect 1670 4607 1676 4641
rect 1710 4607 1716 4641
rect 1670 4569 1716 4607
rect 1670 4535 1676 4569
rect 1710 4535 1716 4569
rect 1670 4497 1716 4535
rect 1670 4463 1676 4497
rect 1710 4463 1716 4497
rect 1670 4425 1716 4463
rect 1670 4391 1676 4425
rect 1710 4391 1716 4425
rect 1670 4353 1716 4391
rect 1670 4319 1676 4353
rect 1710 4319 1716 4353
rect 1670 4281 1716 4319
rect 1670 4247 1676 4281
rect 1710 4247 1716 4281
rect 1670 4209 1716 4247
rect 1670 4175 1676 4209
rect 1710 4175 1716 4209
rect 1670 4137 1716 4175
rect 1670 4103 1676 4137
rect 1710 4103 1716 4137
rect 1670 4065 1716 4103
rect 1670 4031 1676 4065
rect 1710 4031 1716 4065
rect 1670 3993 1716 4031
rect 1670 3959 1676 3993
rect 1710 3959 1716 3993
rect 1670 3944 1716 3959
rect 1766 4929 1812 4944
rect 1766 4895 1772 4929
rect 1806 4895 1812 4929
rect 1766 4857 1812 4895
rect 1766 4823 1772 4857
rect 1806 4823 1812 4857
rect 1766 4785 1812 4823
rect 1766 4751 1772 4785
rect 1806 4751 1812 4785
rect 1766 4713 1812 4751
rect 1766 4679 1772 4713
rect 1806 4679 1812 4713
rect 1766 4641 1812 4679
rect 1766 4607 1772 4641
rect 1806 4607 1812 4641
rect 1766 4569 1812 4607
rect 1766 4535 1772 4569
rect 1806 4535 1812 4569
rect 1766 4497 1812 4535
rect 1766 4463 1772 4497
rect 1806 4463 1812 4497
rect 1766 4425 1812 4463
rect 1766 4391 1772 4425
rect 1806 4391 1812 4425
rect 1766 4353 1812 4391
rect 1766 4319 1772 4353
rect 1806 4319 1812 4353
rect 1766 4281 1812 4319
rect 1766 4247 1772 4281
rect 1806 4247 1812 4281
rect 1766 4209 1812 4247
rect 1766 4175 1772 4209
rect 1806 4175 1812 4209
rect 1766 4137 1812 4175
rect 1766 4103 1772 4137
rect 1806 4103 1812 4137
rect 1766 4065 1812 4103
rect 1766 4031 1772 4065
rect 1806 4031 1812 4065
rect 1766 3993 1812 4031
rect 1766 3959 1772 3993
rect 1806 3959 1812 3993
rect 1766 3944 1812 3959
rect 1862 4929 1908 4944
rect 1862 4895 1868 4929
rect 1902 4895 1908 4929
rect 15512 4943 15558 4981
rect 1862 4857 1908 4895
rect 1862 4823 1868 4857
rect 1902 4823 1908 4857
rect 1862 4785 1908 4823
rect 1862 4751 1868 4785
rect 1902 4751 1908 4785
rect 1862 4713 1908 4751
rect 1862 4679 1868 4713
rect 1902 4679 1908 4713
rect 1862 4641 1908 4679
rect 1862 4607 1868 4641
rect 1902 4607 1908 4641
rect 1862 4569 1908 4607
rect 1862 4535 1868 4569
rect 1902 4535 1908 4569
rect 1862 4497 1908 4535
rect 1862 4463 1868 4497
rect 1902 4463 1908 4497
rect 1862 4425 1908 4463
rect 1862 4391 1868 4425
rect 1902 4391 1908 4425
rect 1862 4353 1908 4391
rect 1862 4319 1868 4353
rect 1902 4319 1908 4353
rect 1862 4281 1908 4319
rect 1862 4247 1868 4281
rect 1902 4247 1908 4281
rect 1862 4209 1908 4247
rect 1862 4175 1868 4209
rect 1902 4175 1908 4209
rect 1862 4137 1908 4175
rect 1862 4103 1868 4137
rect 1902 4103 1908 4137
rect 1862 4065 1908 4103
rect 1862 4031 1868 4065
rect 1902 4031 1908 4065
rect 1862 3993 1908 4031
rect 1862 3959 1868 3993
rect 1902 3959 1908 3993
rect 1862 3944 1908 3959
rect 4434 4913 4480 4928
rect 4434 4879 4440 4913
rect 4474 4879 4480 4913
rect 4434 4841 4480 4879
rect 4434 4807 4440 4841
rect 4474 4807 4480 4841
rect 4434 4769 4480 4807
rect 4434 4735 4440 4769
rect 4474 4735 4480 4769
rect 4434 4697 4480 4735
rect 4434 4663 4440 4697
rect 4474 4663 4480 4697
rect 4434 4625 4480 4663
rect 4434 4591 4440 4625
rect 4474 4591 4480 4625
rect 4434 4553 4480 4591
rect 4434 4519 4440 4553
rect 4474 4519 4480 4553
rect 4434 4481 4480 4519
rect 4434 4447 4440 4481
rect 4474 4447 4480 4481
rect 4434 4409 4480 4447
rect 4434 4375 4440 4409
rect 4474 4375 4480 4409
rect 4434 4337 4480 4375
rect 4434 4303 4440 4337
rect 4474 4303 4480 4337
rect 4434 4265 4480 4303
rect 4434 4231 4440 4265
rect 4474 4231 4480 4265
rect 4434 4193 4480 4231
rect 4434 4159 4440 4193
rect 4474 4159 4480 4193
rect 4434 4121 4480 4159
rect 4434 4087 4440 4121
rect 4474 4087 4480 4121
rect 4434 4049 4480 4087
rect 4434 4015 4440 4049
rect 4474 4015 4480 4049
rect 4434 3977 4480 4015
rect 4434 3943 4440 3977
rect 4474 3943 4480 3977
rect 4434 3928 4480 3943
rect 4530 4913 4576 4928
rect 4530 4879 4536 4913
rect 4570 4879 4576 4913
rect 4530 4841 4576 4879
rect 4530 4807 4536 4841
rect 4570 4807 4576 4841
rect 4530 4769 4576 4807
rect 4530 4735 4536 4769
rect 4570 4735 4576 4769
rect 4530 4697 4576 4735
rect 4530 4663 4536 4697
rect 4570 4663 4576 4697
rect 4530 4625 4576 4663
rect 4530 4591 4536 4625
rect 4570 4591 4576 4625
rect 4530 4553 4576 4591
rect 4530 4519 4536 4553
rect 4570 4519 4576 4553
rect 4530 4481 4576 4519
rect 4530 4447 4536 4481
rect 4570 4447 4576 4481
rect 4530 4409 4576 4447
rect 4530 4375 4536 4409
rect 4570 4375 4576 4409
rect 4530 4337 4576 4375
rect 4530 4303 4536 4337
rect 4570 4303 4576 4337
rect 4530 4265 4576 4303
rect 4530 4231 4536 4265
rect 4570 4231 4576 4265
rect 4530 4193 4576 4231
rect 4530 4159 4536 4193
rect 4570 4159 4576 4193
rect 4530 4121 4576 4159
rect 4530 4087 4536 4121
rect 4570 4087 4576 4121
rect 4530 4049 4576 4087
rect 4530 4015 4536 4049
rect 4570 4015 4576 4049
rect 4530 3977 4576 4015
rect 4530 3943 4536 3977
rect 4570 3943 4576 3977
rect 4530 3928 4576 3943
rect 4626 4913 4672 4928
rect 4626 4879 4632 4913
rect 4666 4879 4672 4913
rect 4626 4841 4672 4879
rect 4626 4807 4632 4841
rect 4666 4807 4672 4841
rect 4626 4769 4672 4807
rect 4626 4735 4632 4769
rect 4666 4735 4672 4769
rect 4626 4697 4672 4735
rect 4626 4663 4632 4697
rect 4666 4663 4672 4697
rect 4626 4625 4672 4663
rect 4626 4591 4632 4625
rect 4666 4591 4672 4625
rect 4626 4553 4672 4591
rect 4626 4519 4632 4553
rect 4666 4519 4672 4553
rect 4626 4481 4672 4519
rect 4626 4447 4632 4481
rect 4666 4447 4672 4481
rect 4626 4409 4672 4447
rect 4626 4375 4632 4409
rect 4666 4375 4672 4409
rect 4626 4337 4672 4375
rect 4626 4303 4632 4337
rect 4666 4303 4672 4337
rect 4626 4265 4672 4303
rect 4626 4231 4632 4265
rect 4666 4231 4672 4265
rect 4626 4193 4672 4231
rect 4626 4159 4632 4193
rect 4666 4159 4672 4193
rect 4626 4121 4672 4159
rect 4626 4087 4632 4121
rect 4666 4087 4672 4121
rect 4626 4049 4672 4087
rect 4626 4015 4632 4049
rect 4666 4015 4672 4049
rect 4626 3977 4672 4015
rect 4626 3943 4632 3977
rect 4666 3943 4672 3977
rect 4626 3928 4672 3943
rect 4722 4913 4768 4928
rect 4722 4879 4728 4913
rect 4762 4879 4768 4913
rect 4722 4841 4768 4879
rect 4722 4807 4728 4841
rect 4762 4807 4768 4841
rect 4722 4769 4768 4807
rect 4722 4735 4728 4769
rect 4762 4735 4768 4769
rect 4722 4697 4768 4735
rect 4722 4663 4728 4697
rect 4762 4663 4768 4697
rect 4722 4625 4768 4663
rect 4722 4591 4728 4625
rect 4762 4591 4768 4625
rect 4722 4553 4768 4591
rect 4722 4519 4728 4553
rect 4762 4519 4768 4553
rect 4722 4481 4768 4519
rect 4722 4447 4728 4481
rect 4762 4447 4768 4481
rect 4722 4409 4768 4447
rect 4722 4375 4728 4409
rect 4762 4375 4768 4409
rect 4722 4337 4768 4375
rect 4722 4303 4728 4337
rect 4762 4303 4768 4337
rect 4722 4265 4768 4303
rect 4722 4231 4728 4265
rect 4762 4231 4768 4265
rect 4722 4193 4768 4231
rect 4722 4159 4728 4193
rect 4762 4159 4768 4193
rect 4722 4121 4768 4159
rect 4722 4087 4728 4121
rect 4762 4087 4768 4121
rect 4722 4049 4768 4087
rect 4722 4015 4728 4049
rect 4762 4015 4768 4049
rect 4722 3977 4768 4015
rect 4722 3943 4728 3977
rect 4762 3943 4768 3977
rect 4722 3928 4768 3943
rect 4818 4913 4864 4928
rect 4818 4879 4824 4913
rect 4858 4879 4864 4913
rect 4818 4841 4864 4879
rect 4818 4807 4824 4841
rect 4858 4807 4864 4841
rect 4818 4769 4864 4807
rect 4818 4735 4824 4769
rect 4858 4735 4864 4769
rect 4818 4697 4864 4735
rect 4818 4663 4824 4697
rect 4858 4663 4864 4697
rect 4818 4625 4864 4663
rect 4818 4591 4824 4625
rect 4858 4591 4864 4625
rect 4818 4553 4864 4591
rect 4818 4519 4824 4553
rect 4858 4519 4864 4553
rect 4818 4481 4864 4519
rect 4818 4447 4824 4481
rect 4858 4447 4864 4481
rect 4818 4409 4864 4447
rect 4818 4375 4824 4409
rect 4858 4375 4864 4409
rect 4818 4337 4864 4375
rect 4818 4303 4824 4337
rect 4858 4303 4864 4337
rect 4818 4265 4864 4303
rect 4818 4231 4824 4265
rect 4858 4231 4864 4265
rect 4818 4193 4864 4231
rect 4818 4159 4824 4193
rect 4858 4159 4864 4193
rect 4818 4121 4864 4159
rect 4818 4087 4824 4121
rect 4858 4087 4864 4121
rect 4818 4049 4864 4087
rect 4818 4015 4824 4049
rect 4858 4015 4864 4049
rect 4818 3977 4864 4015
rect 4818 3943 4824 3977
rect 4858 3943 4864 3977
rect 4818 3928 4864 3943
rect 7464 4913 7510 4928
rect 7464 4879 7470 4913
rect 7504 4879 7510 4913
rect 7464 4841 7510 4879
rect 7464 4807 7470 4841
rect 7504 4807 7510 4841
rect 7464 4769 7510 4807
rect 7464 4735 7470 4769
rect 7504 4735 7510 4769
rect 7464 4697 7510 4735
rect 7464 4663 7470 4697
rect 7504 4663 7510 4697
rect 7464 4625 7510 4663
rect 7464 4591 7470 4625
rect 7504 4591 7510 4625
rect 7464 4553 7510 4591
rect 7464 4519 7470 4553
rect 7504 4519 7510 4553
rect 7464 4481 7510 4519
rect 7464 4447 7470 4481
rect 7504 4447 7510 4481
rect 7464 4409 7510 4447
rect 7464 4375 7470 4409
rect 7504 4375 7510 4409
rect 7464 4337 7510 4375
rect 7464 4303 7470 4337
rect 7504 4303 7510 4337
rect 7464 4265 7510 4303
rect 7464 4231 7470 4265
rect 7504 4231 7510 4265
rect 7464 4193 7510 4231
rect 7464 4159 7470 4193
rect 7504 4159 7510 4193
rect 7464 4121 7510 4159
rect 7464 4087 7470 4121
rect 7504 4087 7510 4121
rect 7464 4049 7510 4087
rect 7464 4015 7470 4049
rect 7504 4015 7510 4049
rect 7464 3977 7510 4015
rect 7464 3943 7470 3977
rect 7504 3943 7510 3977
rect 7464 3928 7510 3943
rect 7560 4913 7606 4928
rect 7560 4879 7566 4913
rect 7600 4879 7606 4913
rect 7560 4841 7606 4879
rect 7560 4807 7566 4841
rect 7600 4807 7606 4841
rect 7560 4769 7606 4807
rect 7560 4735 7566 4769
rect 7600 4735 7606 4769
rect 7560 4697 7606 4735
rect 7560 4663 7566 4697
rect 7600 4663 7606 4697
rect 7560 4625 7606 4663
rect 7560 4591 7566 4625
rect 7600 4591 7606 4625
rect 7560 4553 7606 4591
rect 7560 4519 7566 4553
rect 7600 4519 7606 4553
rect 7560 4481 7606 4519
rect 7560 4447 7566 4481
rect 7600 4447 7606 4481
rect 7560 4409 7606 4447
rect 7560 4375 7566 4409
rect 7600 4375 7606 4409
rect 7560 4337 7606 4375
rect 7560 4303 7566 4337
rect 7600 4303 7606 4337
rect 7560 4265 7606 4303
rect 7560 4231 7566 4265
rect 7600 4231 7606 4265
rect 7560 4193 7606 4231
rect 7560 4159 7566 4193
rect 7600 4159 7606 4193
rect 7560 4121 7606 4159
rect 7560 4087 7566 4121
rect 7600 4087 7606 4121
rect 7560 4049 7606 4087
rect 7560 4015 7566 4049
rect 7600 4015 7606 4049
rect 7560 3977 7606 4015
rect 7560 3943 7566 3977
rect 7600 3943 7606 3977
rect 7560 3928 7606 3943
rect 7656 4913 7702 4928
rect 7656 4879 7662 4913
rect 7696 4879 7702 4913
rect 7656 4841 7702 4879
rect 7656 4807 7662 4841
rect 7696 4807 7702 4841
rect 7656 4769 7702 4807
rect 7656 4735 7662 4769
rect 7696 4735 7702 4769
rect 7656 4697 7702 4735
rect 7656 4663 7662 4697
rect 7696 4663 7702 4697
rect 7656 4625 7702 4663
rect 7656 4591 7662 4625
rect 7696 4591 7702 4625
rect 7656 4553 7702 4591
rect 7656 4519 7662 4553
rect 7696 4519 7702 4553
rect 7656 4481 7702 4519
rect 7656 4447 7662 4481
rect 7696 4447 7702 4481
rect 7656 4409 7702 4447
rect 7656 4375 7662 4409
rect 7696 4375 7702 4409
rect 7656 4337 7702 4375
rect 7656 4303 7662 4337
rect 7696 4303 7702 4337
rect 7656 4265 7702 4303
rect 7656 4231 7662 4265
rect 7696 4231 7702 4265
rect 7656 4193 7702 4231
rect 7656 4159 7662 4193
rect 7696 4159 7702 4193
rect 7656 4121 7702 4159
rect 7656 4087 7662 4121
rect 7696 4087 7702 4121
rect 7656 4049 7702 4087
rect 7656 4015 7662 4049
rect 7696 4015 7702 4049
rect 7656 3977 7702 4015
rect 7656 3943 7662 3977
rect 7696 3943 7702 3977
rect 7656 3928 7702 3943
rect 7752 4913 7798 4928
rect 7752 4879 7758 4913
rect 7792 4879 7798 4913
rect 7752 4841 7798 4879
rect 7752 4807 7758 4841
rect 7792 4807 7798 4841
rect 7752 4769 7798 4807
rect 7752 4735 7758 4769
rect 7792 4735 7798 4769
rect 7752 4697 7798 4735
rect 7752 4663 7758 4697
rect 7792 4663 7798 4697
rect 7752 4625 7798 4663
rect 7752 4591 7758 4625
rect 7792 4591 7798 4625
rect 7752 4553 7798 4591
rect 7752 4519 7758 4553
rect 7792 4519 7798 4553
rect 7752 4481 7798 4519
rect 7752 4447 7758 4481
rect 7792 4447 7798 4481
rect 7752 4409 7798 4447
rect 7752 4375 7758 4409
rect 7792 4375 7798 4409
rect 7752 4337 7798 4375
rect 7752 4303 7758 4337
rect 7792 4303 7798 4337
rect 7752 4265 7798 4303
rect 7752 4231 7758 4265
rect 7792 4231 7798 4265
rect 7752 4193 7798 4231
rect 7752 4159 7758 4193
rect 7792 4159 7798 4193
rect 7752 4121 7798 4159
rect 7752 4087 7758 4121
rect 7792 4087 7798 4121
rect 7752 4049 7798 4087
rect 7752 4015 7758 4049
rect 7792 4015 7798 4049
rect 7752 3977 7798 4015
rect 7752 3943 7758 3977
rect 7792 3943 7798 3977
rect 7752 3928 7798 3943
rect 7848 4913 7894 4928
rect 7848 4879 7854 4913
rect 7888 4879 7894 4913
rect 7848 4841 7894 4879
rect 7848 4807 7854 4841
rect 7888 4807 7894 4841
rect 7848 4769 7894 4807
rect 7848 4735 7854 4769
rect 7888 4735 7894 4769
rect 7848 4697 7894 4735
rect 7848 4663 7854 4697
rect 7888 4663 7894 4697
rect 7848 4625 7894 4663
rect 7848 4591 7854 4625
rect 7888 4591 7894 4625
rect 7848 4553 7894 4591
rect 7848 4519 7854 4553
rect 7888 4519 7894 4553
rect 7848 4481 7894 4519
rect 7848 4447 7854 4481
rect 7888 4447 7894 4481
rect 7848 4409 7894 4447
rect 7848 4375 7854 4409
rect 7888 4375 7894 4409
rect 7848 4337 7894 4375
rect 7848 4303 7854 4337
rect 7888 4303 7894 4337
rect 7848 4265 7894 4303
rect 7848 4231 7854 4265
rect 7888 4231 7894 4265
rect 7848 4193 7894 4231
rect 7848 4159 7854 4193
rect 7888 4159 7894 4193
rect 7848 4121 7894 4159
rect 7848 4087 7854 4121
rect 7888 4087 7894 4121
rect 7848 4049 7894 4087
rect 7848 4015 7854 4049
rect 7888 4015 7894 4049
rect 7848 3977 7894 4015
rect 7848 3943 7854 3977
rect 7888 3943 7894 3977
rect 7848 3928 7894 3943
rect 10552 4911 10598 4926
rect 10552 4877 10558 4911
rect 10592 4877 10598 4911
rect 10552 4839 10598 4877
rect 10552 4805 10558 4839
rect 10592 4805 10598 4839
rect 10552 4767 10598 4805
rect 10552 4733 10558 4767
rect 10592 4733 10598 4767
rect 10552 4695 10598 4733
rect 10552 4661 10558 4695
rect 10592 4661 10598 4695
rect 10552 4623 10598 4661
rect 10552 4589 10558 4623
rect 10592 4589 10598 4623
rect 10552 4551 10598 4589
rect 10552 4517 10558 4551
rect 10592 4517 10598 4551
rect 10552 4479 10598 4517
rect 10552 4445 10558 4479
rect 10592 4445 10598 4479
rect 10552 4407 10598 4445
rect 10552 4373 10558 4407
rect 10592 4373 10598 4407
rect 10552 4335 10598 4373
rect 10552 4301 10558 4335
rect 10592 4301 10598 4335
rect 10552 4263 10598 4301
rect 10552 4229 10558 4263
rect 10592 4229 10598 4263
rect 10552 4191 10598 4229
rect 10552 4157 10558 4191
rect 10592 4157 10598 4191
rect 10552 4119 10598 4157
rect 10552 4085 10558 4119
rect 10592 4085 10598 4119
rect 10552 4047 10598 4085
rect 10552 4013 10558 4047
rect 10592 4013 10598 4047
rect 10552 3975 10598 4013
rect 10552 3941 10558 3975
rect 10592 3941 10598 3975
rect 10552 3926 10598 3941
rect 10648 4911 10694 4926
rect 10648 4877 10654 4911
rect 10688 4877 10694 4911
rect 10648 4839 10694 4877
rect 10648 4805 10654 4839
rect 10688 4805 10694 4839
rect 10648 4767 10694 4805
rect 10648 4733 10654 4767
rect 10688 4733 10694 4767
rect 10648 4695 10694 4733
rect 10648 4661 10654 4695
rect 10688 4661 10694 4695
rect 10648 4623 10694 4661
rect 10648 4589 10654 4623
rect 10688 4589 10694 4623
rect 10648 4551 10694 4589
rect 10648 4517 10654 4551
rect 10688 4517 10694 4551
rect 10648 4479 10694 4517
rect 10648 4445 10654 4479
rect 10688 4445 10694 4479
rect 10648 4407 10694 4445
rect 10648 4373 10654 4407
rect 10688 4373 10694 4407
rect 10648 4335 10694 4373
rect 10648 4301 10654 4335
rect 10688 4301 10694 4335
rect 10648 4263 10694 4301
rect 10648 4229 10654 4263
rect 10688 4229 10694 4263
rect 10648 4191 10694 4229
rect 10648 4157 10654 4191
rect 10688 4157 10694 4191
rect 10648 4119 10694 4157
rect 10648 4085 10654 4119
rect 10688 4085 10694 4119
rect 10648 4047 10694 4085
rect 10648 4013 10654 4047
rect 10688 4013 10694 4047
rect 10648 3975 10694 4013
rect 10648 3941 10654 3975
rect 10688 3941 10694 3975
rect 10648 3926 10694 3941
rect 10744 4911 10790 4926
rect 10744 4877 10750 4911
rect 10784 4877 10790 4911
rect 10744 4839 10790 4877
rect 10744 4805 10750 4839
rect 10784 4805 10790 4839
rect 10744 4767 10790 4805
rect 10744 4733 10750 4767
rect 10784 4733 10790 4767
rect 10744 4695 10790 4733
rect 10744 4661 10750 4695
rect 10784 4661 10790 4695
rect 10744 4623 10790 4661
rect 10744 4589 10750 4623
rect 10784 4589 10790 4623
rect 10744 4551 10790 4589
rect 10744 4517 10750 4551
rect 10784 4517 10790 4551
rect 10744 4479 10790 4517
rect 10744 4445 10750 4479
rect 10784 4445 10790 4479
rect 10744 4407 10790 4445
rect 10744 4373 10750 4407
rect 10784 4373 10790 4407
rect 10744 4335 10790 4373
rect 10744 4301 10750 4335
rect 10784 4301 10790 4335
rect 10744 4263 10790 4301
rect 10744 4229 10750 4263
rect 10784 4229 10790 4263
rect 10744 4191 10790 4229
rect 10744 4157 10750 4191
rect 10784 4157 10790 4191
rect 10744 4119 10790 4157
rect 10744 4085 10750 4119
rect 10784 4085 10790 4119
rect 10744 4047 10790 4085
rect 10744 4013 10750 4047
rect 10784 4013 10790 4047
rect 10744 3975 10790 4013
rect 10744 3941 10750 3975
rect 10784 3941 10790 3975
rect 10744 3926 10790 3941
rect 10840 4911 10886 4926
rect 10840 4877 10846 4911
rect 10880 4877 10886 4911
rect 10840 4839 10886 4877
rect 10840 4805 10846 4839
rect 10880 4805 10886 4839
rect 10840 4767 10886 4805
rect 10840 4733 10846 4767
rect 10880 4733 10886 4767
rect 10840 4695 10886 4733
rect 10840 4661 10846 4695
rect 10880 4661 10886 4695
rect 10840 4623 10886 4661
rect 10840 4589 10846 4623
rect 10880 4589 10886 4623
rect 10840 4551 10886 4589
rect 10840 4517 10846 4551
rect 10880 4517 10886 4551
rect 10840 4479 10886 4517
rect 10840 4445 10846 4479
rect 10880 4445 10886 4479
rect 10840 4407 10886 4445
rect 10840 4373 10846 4407
rect 10880 4373 10886 4407
rect 10840 4335 10886 4373
rect 10840 4301 10846 4335
rect 10880 4301 10886 4335
rect 10840 4263 10886 4301
rect 10840 4229 10846 4263
rect 10880 4229 10886 4263
rect 10840 4191 10886 4229
rect 10840 4157 10846 4191
rect 10880 4157 10886 4191
rect 10840 4119 10886 4157
rect 10840 4085 10846 4119
rect 10880 4085 10886 4119
rect 10840 4047 10886 4085
rect 10840 4013 10846 4047
rect 10880 4013 10886 4047
rect 10840 3975 10886 4013
rect 10840 3941 10846 3975
rect 10880 3941 10886 3975
rect 10840 3926 10886 3941
rect 10936 4911 10982 4926
rect 10936 4877 10942 4911
rect 10976 4877 10982 4911
rect 15512 4909 15518 4943
rect 15552 4909 15558 4943
rect 10936 4839 10982 4877
rect 10936 4805 10942 4839
rect 10976 4805 10982 4839
rect 10936 4767 10982 4805
rect 10936 4733 10942 4767
rect 10976 4733 10982 4767
rect 10936 4695 10982 4733
rect 10936 4661 10942 4695
rect 10976 4661 10982 4695
rect 10936 4623 10982 4661
rect 10936 4589 10942 4623
rect 10976 4589 10982 4623
rect 10936 4551 10982 4589
rect 10936 4517 10942 4551
rect 10976 4517 10982 4551
rect 10936 4479 10982 4517
rect 10936 4445 10942 4479
rect 10976 4445 10982 4479
rect 10936 4407 10982 4445
rect 10936 4373 10942 4407
rect 10976 4373 10982 4407
rect 10936 4335 10982 4373
rect 10936 4301 10942 4335
rect 10976 4301 10982 4335
rect 10936 4263 10982 4301
rect 10936 4229 10942 4263
rect 10976 4229 10982 4263
rect 10936 4191 10982 4229
rect 10936 4157 10942 4191
rect 10976 4157 10982 4191
rect 10936 4119 10982 4157
rect 10936 4085 10942 4119
rect 10976 4085 10982 4119
rect 10936 4047 10982 4085
rect 10936 4013 10942 4047
rect 10976 4013 10982 4047
rect 10936 3975 10982 4013
rect 10936 3941 10942 3975
rect 10976 3941 10982 3975
rect 10936 3926 10982 3941
rect 13708 4885 13754 4900
rect 13708 4851 13714 4885
rect 13748 4851 13754 4885
rect 13708 4813 13754 4851
rect 13708 4779 13714 4813
rect 13748 4779 13754 4813
rect 13708 4741 13754 4779
rect 13708 4707 13714 4741
rect 13748 4707 13754 4741
rect 13708 4669 13754 4707
rect 13708 4635 13714 4669
rect 13748 4635 13754 4669
rect 13708 4597 13754 4635
rect 13708 4563 13714 4597
rect 13748 4563 13754 4597
rect 13708 4525 13754 4563
rect 13708 4491 13714 4525
rect 13748 4491 13754 4525
rect 13708 4453 13754 4491
rect 13708 4419 13714 4453
rect 13748 4419 13754 4453
rect 13708 4381 13754 4419
rect 13708 4347 13714 4381
rect 13748 4347 13754 4381
rect 13708 4309 13754 4347
rect 13708 4275 13714 4309
rect 13748 4275 13754 4309
rect 13708 4237 13754 4275
rect 13708 4203 13714 4237
rect 13748 4203 13754 4237
rect 13708 4165 13754 4203
rect 13708 4131 13714 4165
rect 13748 4131 13754 4165
rect 13708 4093 13754 4131
rect 13708 4059 13714 4093
rect 13748 4059 13754 4093
rect 13708 4021 13754 4059
rect 13708 3987 13714 4021
rect 13748 3987 13754 4021
rect 13708 3949 13754 3987
rect 13708 3915 13714 3949
rect 13748 3915 13754 3949
rect 13708 3900 13754 3915
rect 13804 4885 13850 4900
rect 13804 4851 13810 4885
rect 13844 4851 13850 4885
rect 13804 4813 13850 4851
rect 13804 4779 13810 4813
rect 13844 4779 13850 4813
rect 13804 4741 13850 4779
rect 13804 4707 13810 4741
rect 13844 4707 13850 4741
rect 13804 4669 13850 4707
rect 13804 4635 13810 4669
rect 13844 4635 13850 4669
rect 13804 4597 13850 4635
rect 13804 4563 13810 4597
rect 13844 4563 13850 4597
rect 13804 4525 13850 4563
rect 13804 4491 13810 4525
rect 13844 4491 13850 4525
rect 13804 4453 13850 4491
rect 13804 4419 13810 4453
rect 13844 4419 13850 4453
rect 13804 4381 13850 4419
rect 13804 4347 13810 4381
rect 13844 4347 13850 4381
rect 13804 4309 13850 4347
rect 13804 4275 13810 4309
rect 13844 4275 13850 4309
rect 13804 4237 13850 4275
rect 13804 4203 13810 4237
rect 13844 4203 13850 4237
rect 13804 4165 13850 4203
rect 13804 4131 13810 4165
rect 13844 4131 13850 4165
rect 13804 4093 13850 4131
rect 13804 4059 13810 4093
rect 13844 4059 13850 4093
rect 13804 4021 13850 4059
rect 13804 3987 13810 4021
rect 13844 3987 13850 4021
rect 13804 3949 13850 3987
rect 13804 3915 13810 3949
rect 13844 3915 13850 3949
rect 13804 3900 13850 3915
rect 13900 4885 13946 4900
rect 13900 4851 13906 4885
rect 13940 4851 13946 4885
rect 13900 4813 13946 4851
rect 13900 4779 13906 4813
rect 13940 4779 13946 4813
rect 13900 4741 13946 4779
rect 13900 4707 13906 4741
rect 13940 4707 13946 4741
rect 13900 4669 13946 4707
rect 13900 4635 13906 4669
rect 13940 4635 13946 4669
rect 13900 4597 13946 4635
rect 13900 4563 13906 4597
rect 13940 4563 13946 4597
rect 13900 4525 13946 4563
rect 13900 4491 13906 4525
rect 13940 4491 13946 4525
rect 13900 4453 13946 4491
rect 13900 4419 13906 4453
rect 13940 4419 13946 4453
rect 13900 4381 13946 4419
rect 13900 4347 13906 4381
rect 13940 4347 13946 4381
rect 13900 4309 13946 4347
rect 13900 4275 13906 4309
rect 13940 4275 13946 4309
rect 13900 4237 13946 4275
rect 13900 4203 13906 4237
rect 13940 4203 13946 4237
rect 13900 4165 13946 4203
rect 13900 4131 13906 4165
rect 13940 4131 13946 4165
rect 13900 4093 13946 4131
rect 13900 4059 13906 4093
rect 13940 4059 13946 4093
rect 13900 4021 13946 4059
rect 13900 3987 13906 4021
rect 13940 3987 13946 4021
rect 13900 3949 13946 3987
rect 13900 3915 13906 3949
rect 13940 3915 13946 3949
rect 13900 3900 13946 3915
rect 13996 4885 14042 4900
rect 13996 4851 14002 4885
rect 14036 4851 14042 4885
rect 13996 4813 14042 4851
rect 13996 4779 14002 4813
rect 14036 4779 14042 4813
rect 13996 4741 14042 4779
rect 13996 4707 14002 4741
rect 14036 4707 14042 4741
rect 13996 4669 14042 4707
rect 13996 4635 14002 4669
rect 14036 4635 14042 4669
rect 13996 4597 14042 4635
rect 13996 4563 14002 4597
rect 14036 4563 14042 4597
rect 13996 4525 14042 4563
rect 13996 4491 14002 4525
rect 14036 4491 14042 4525
rect 13996 4453 14042 4491
rect 13996 4419 14002 4453
rect 14036 4419 14042 4453
rect 13996 4381 14042 4419
rect 13996 4347 14002 4381
rect 14036 4347 14042 4381
rect 13996 4309 14042 4347
rect 13996 4275 14002 4309
rect 14036 4275 14042 4309
rect 13996 4237 14042 4275
rect 13996 4203 14002 4237
rect 14036 4203 14042 4237
rect 13996 4165 14042 4203
rect 13996 4131 14002 4165
rect 14036 4131 14042 4165
rect 13996 4093 14042 4131
rect 13996 4059 14002 4093
rect 14036 4059 14042 4093
rect 13996 4021 14042 4059
rect 13996 3987 14002 4021
rect 14036 3987 14042 4021
rect 13996 3949 14042 3987
rect 13996 3915 14002 3949
rect 14036 3915 14042 3949
rect 13996 3900 14042 3915
rect 14092 4885 14138 4900
rect 14092 4851 14098 4885
rect 14132 4851 14138 4885
rect 14092 4813 14138 4851
rect 14092 4779 14098 4813
rect 14132 4779 14138 4813
rect 14092 4741 14138 4779
rect 14092 4707 14098 4741
rect 14132 4707 14138 4741
rect 14092 4669 14138 4707
rect 14092 4635 14098 4669
rect 14132 4635 14138 4669
rect 14092 4597 14138 4635
rect 14092 4563 14098 4597
rect 14132 4563 14138 4597
rect 14092 4525 14138 4563
rect 14092 4491 14098 4525
rect 14132 4491 14138 4525
rect 14092 4453 14138 4491
rect 14092 4419 14098 4453
rect 14132 4419 14138 4453
rect 14092 4381 14138 4419
rect 14092 4347 14098 4381
rect 14132 4347 14138 4381
rect 14092 4309 14138 4347
rect 14092 4275 14098 4309
rect 14132 4275 14138 4309
rect 14092 4237 14138 4275
rect 14092 4203 14098 4237
rect 14132 4203 14138 4237
rect 14092 4165 14138 4203
rect 14092 4131 14098 4165
rect 14132 4131 14138 4165
rect 14092 4093 14138 4131
rect 14092 4059 14098 4093
rect 14132 4059 14138 4093
rect 14092 4021 14138 4059
rect 14092 3987 14098 4021
rect 14132 3987 14138 4021
rect 14092 3949 14138 3987
rect 14092 3915 14098 3949
rect 14132 3915 14138 3949
rect 15512 4871 15558 4909
rect 15512 4837 15518 4871
rect 15552 4837 15558 4871
rect 15512 4799 15558 4837
rect 15512 4765 15518 4799
rect 15552 4765 15558 4799
rect 15512 4727 15558 4765
rect 15512 4693 15518 4727
rect 15552 4693 15558 4727
rect 15512 4655 15558 4693
rect 15512 4621 15518 4655
rect 15552 4621 15558 4655
rect 15512 4583 15558 4621
rect 15512 4549 15518 4583
rect 15552 4549 15558 4583
rect 15512 4511 15558 4549
rect 15512 4477 15518 4511
rect 15552 4477 15558 4511
rect 15512 4439 15558 4477
rect 15512 4405 15518 4439
rect 15552 4405 15558 4439
rect 15512 4367 15558 4405
rect 15512 4333 15518 4367
rect 15552 4333 15558 4367
rect 15512 4295 15558 4333
rect 15512 4261 15518 4295
rect 15552 4261 15558 4295
rect 15512 4223 15558 4261
rect 15512 4189 15518 4223
rect 15552 4189 15558 4223
rect 15512 4151 15558 4189
rect 15512 4117 15518 4151
rect 15552 4117 15558 4151
rect 15512 4079 15558 4117
rect 15512 4045 15518 4079
rect 15552 4045 15558 4079
rect 15512 4007 15558 4045
rect 15512 3973 15518 4007
rect 15552 3973 15558 4007
rect 15512 3926 15558 3973
rect 15608 5879 15654 5926
rect 15608 5845 15614 5879
rect 15648 5845 15654 5879
rect 15608 5807 15654 5845
rect 15608 5773 15614 5807
rect 15648 5773 15654 5807
rect 15608 5735 15654 5773
rect 15608 5701 15614 5735
rect 15648 5701 15654 5735
rect 15608 5663 15654 5701
rect 15608 5629 15614 5663
rect 15648 5629 15654 5663
rect 15608 5591 15654 5629
rect 15608 5557 15614 5591
rect 15648 5557 15654 5591
rect 15608 5519 15654 5557
rect 15608 5485 15614 5519
rect 15648 5485 15654 5519
rect 15608 5447 15654 5485
rect 15608 5413 15614 5447
rect 15648 5413 15654 5447
rect 15608 5375 15654 5413
rect 15608 5341 15614 5375
rect 15648 5341 15654 5375
rect 15608 5303 15654 5341
rect 15608 5269 15614 5303
rect 15648 5269 15654 5303
rect 15608 5231 15654 5269
rect 15608 5197 15614 5231
rect 15648 5197 15654 5231
rect 15608 5159 15654 5197
rect 15608 5125 15614 5159
rect 15648 5125 15654 5159
rect 15608 5087 15654 5125
rect 15608 5053 15614 5087
rect 15648 5053 15654 5087
rect 15608 5015 15654 5053
rect 15608 4981 15614 5015
rect 15648 4981 15654 5015
rect 15608 4943 15654 4981
rect 15608 4909 15614 4943
rect 15648 4909 15654 4943
rect 15608 4871 15654 4909
rect 15608 4837 15614 4871
rect 15648 4837 15654 4871
rect 15608 4799 15654 4837
rect 15608 4765 15614 4799
rect 15648 4765 15654 4799
rect 15608 4727 15654 4765
rect 15608 4693 15614 4727
rect 15648 4693 15654 4727
rect 15608 4655 15654 4693
rect 15608 4621 15614 4655
rect 15648 4621 15654 4655
rect 15608 4583 15654 4621
rect 15608 4549 15614 4583
rect 15648 4549 15654 4583
rect 15608 4511 15654 4549
rect 15608 4477 15614 4511
rect 15648 4477 15654 4511
rect 15608 4439 15654 4477
rect 15608 4405 15614 4439
rect 15648 4405 15654 4439
rect 15608 4367 15654 4405
rect 15608 4333 15614 4367
rect 15648 4333 15654 4367
rect 15608 4295 15654 4333
rect 15608 4261 15614 4295
rect 15648 4261 15654 4295
rect 15608 4223 15654 4261
rect 15608 4189 15614 4223
rect 15648 4189 15654 4223
rect 15608 4151 15654 4189
rect 15608 4117 15614 4151
rect 15648 4117 15654 4151
rect 15608 4079 15654 4117
rect 15608 4045 15614 4079
rect 15648 4045 15654 4079
rect 15608 4007 15654 4045
rect 15608 3973 15614 4007
rect 15648 3973 15654 4007
rect 15608 3926 15654 3973
rect 15704 5879 15750 5926
rect 15704 5845 15710 5879
rect 15744 5845 15750 5879
rect 15704 5807 15750 5845
rect 15704 5773 15710 5807
rect 15744 5773 15750 5807
rect 15704 5735 15750 5773
rect 15704 5701 15710 5735
rect 15744 5701 15750 5735
rect 15704 5663 15750 5701
rect 15704 5629 15710 5663
rect 15744 5629 15750 5663
rect 15704 5591 15750 5629
rect 15704 5557 15710 5591
rect 15744 5557 15750 5591
rect 15704 5519 15750 5557
rect 15704 5485 15710 5519
rect 15744 5485 15750 5519
rect 15704 5447 15750 5485
rect 15704 5413 15710 5447
rect 15744 5413 15750 5447
rect 15704 5375 15750 5413
rect 15704 5341 15710 5375
rect 15744 5341 15750 5375
rect 15704 5303 15750 5341
rect 15704 5269 15710 5303
rect 15744 5269 15750 5303
rect 16962 5487 17252 5500
rect 16962 5307 16985 5487
rect 17229 5307 17252 5487
rect 16962 5294 17252 5307
rect 18960 5484 19252 5500
rect 18960 5304 18984 5484
rect 19228 5304 19252 5484
rect 18960 5288 19252 5304
rect 20962 5484 21252 5500
rect 20962 5304 20985 5484
rect 21229 5304 21252 5484
rect 20962 5288 21252 5304
rect 23508 5483 23796 5498
rect 23508 5303 23530 5483
rect 23774 5303 23796 5483
rect 23508 5288 23796 5303
rect 25508 5484 25798 5500
rect 25508 5304 25531 5484
rect 25775 5304 25798 5484
rect 25508 5288 25798 5304
rect 27508 5483 27798 5498
rect 27508 5303 27531 5483
rect 27775 5303 27798 5483
rect 27508 5288 27798 5303
rect 15704 5231 15750 5269
rect 15704 5197 15710 5231
rect 15744 5197 15750 5231
rect 15704 5159 15750 5197
rect 15704 5125 15710 5159
rect 15744 5125 15750 5159
rect 15704 5087 15750 5125
rect 15704 5053 15710 5087
rect 15744 5053 15750 5087
rect 15704 5015 15750 5053
rect 15704 4981 15710 5015
rect 15744 4981 15750 5015
rect 15704 4943 15750 4981
rect 15704 4909 15710 4943
rect 15744 4909 15750 4943
rect 15704 4871 15750 4909
rect 15704 4837 15710 4871
rect 15744 4837 15750 4871
rect 15704 4799 15750 4837
rect 15704 4765 15710 4799
rect 15744 4765 15750 4799
rect 15704 4727 15750 4765
rect 15704 4693 15710 4727
rect 15744 4693 15750 4727
rect 15704 4655 15750 4693
rect 15704 4621 15710 4655
rect 15744 4621 15750 4655
rect 15704 4583 15750 4621
rect 15704 4549 15710 4583
rect 15744 4549 15750 4583
rect 15704 4511 15750 4549
rect 15704 4477 15710 4511
rect 15744 4477 15750 4511
rect 15704 4439 15750 4477
rect 15704 4405 15710 4439
rect 15744 4405 15750 4439
rect 15704 4367 15750 4405
rect 15704 4333 15710 4367
rect 15744 4333 15750 4367
rect 15704 4295 15750 4333
rect 15704 4261 15710 4295
rect 15744 4261 15750 4295
rect 15704 4223 15750 4261
rect 15704 4189 15710 4223
rect 15744 4189 15750 4223
rect 15704 4151 15750 4189
rect 15704 4117 15710 4151
rect 15744 4117 15750 4151
rect 16776 5115 16822 5130
rect 16776 5081 16782 5115
rect 16816 5081 16822 5115
rect 16776 5043 16822 5081
rect 16776 5009 16782 5043
rect 16816 5009 16822 5043
rect 16776 4971 16822 5009
rect 16776 4937 16782 4971
rect 16816 4937 16822 4971
rect 16776 4899 16822 4937
rect 16776 4865 16782 4899
rect 16816 4865 16822 4899
rect 16776 4827 16822 4865
rect 16776 4793 16782 4827
rect 16816 4793 16822 4827
rect 16776 4755 16822 4793
rect 16776 4721 16782 4755
rect 16816 4721 16822 4755
rect 16776 4683 16822 4721
rect 16776 4649 16782 4683
rect 16816 4649 16822 4683
rect 16776 4611 16822 4649
rect 16776 4577 16782 4611
rect 16816 4577 16822 4611
rect 16776 4539 16822 4577
rect 16776 4505 16782 4539
rect 16816 4505 16822 4539
rect 16776 4467 16822 4505
rect 16776 4433 16782 4467
rect 16816 4433 16822 4467
rect 16776 4395 16822 4433
rect 16776 4361 16782 4395
rect 16816 4361 16822 4395
rect 16776 4323 16822 4361
rect 16776 4289 16782 4323
rect 16816 4289 16822 4323
rect 16776 4251 16822 4289
rect 16776 4217 16782 4251
rect 16816 4217 16822 4251
rect 16776 4179 16822 4217
rect 16776 4145 16782 4179
rect 16816 4145 16822 4179
rect 16776 4130 16822 4145
rect 16872 5115 16918 5130
rect 16872 5081 16878 5115
rect 16912 5081 16918 5115
rect 16872 5043 16918 5081
rect 16872 5009 16878 5043
rect 16912 5009 16918 5043
rect 16872 4971 16918 5009
rect 16872 4937 16878 4971
rect 16912 4937 16918 4971
rect 16872 4899 16918 4937
rect 16872 4865 16878 4899
rect 16912 4865 16918 4899
rect 16872 4827 16918 4865
rect 16872 4793 16878 4827
rect 16912 4793 16918 4827
rect 16872 4755 16918 4793
rect 16872 4721 16878 4755
rect 16912 4721 16918 4755
rect 16872 4683 16918 4721
rect 16872 4649 16878 4683
rect 16912 4649 16918 4683
rect 16872 4611 16918 4649
rect 16872 4577 16878 4611
rect 16912 4577 16918 4611
rect 16872 4539 16918 4577
rect 16872 4505 16878 4539
rect 16912 4505 16918 4539
rect 16872 4467 16918 4505
rect 16872 4433 16878 4467
rect 16912 4433 16918 4467
rect 16872 4395 16918 4433
rect 16872 4361 16878 4395
rect 16912 4361 16918 4395
rect 16872 4323 16918 4361
rect 16872 4289 16878 4323
rect 16912 4289 16918 4323
rect 16872 4251 16918 4289
rect 16872 4217 16878 4251
rect 16912 4217 16918 4251
rect 16872 4179 16918 4217
rect 16872 4145 16878 4179
rect 16912 4145 16918 4179
rect 16872 4130 16918 4145
rect 16968 5115 17014 5130
rect 16968 5081 16974 5115
rect 17008 5081 17014 5115
rect 16968 5043 17014 5081
rect 16968 5009 16974 5043
rect 17008 5009 17014 5043
rect 16968 4971 17014 5009
rect 16968 4937 16974 4971
rect 17008 4937 17014 4971
rect 16968 4899 17014 4937
rect 16968 4865 16974 4899
rect 17008 4865 17014 4899
rect 16968 4827 17014 4865
rect 16968 4793 16974 4827
rect 17008 4793 17014 4827
rect 16968 4755 17014 4793
rect 16968 4721 16974 4755
rect 17008 4721 17014 4755
rect 16968 4683 17014 4721
rect 16968 4649 16974 4683
rect 17008 4649 17014 4683
rect 16968 4611 17014 4649
rect 16968 4577 16974 4611
rect 17008 4577 17014 4611
rect 16968 4539 17014 4577
rect 16968 4505 16974 4539
rect 17008 4505 17014 4539
rect 16968 4467 17014 4505
rect 16968 4433 16974 4467
rect 17008 4433 17014 4467
rect 16968 4395 17014 4433
rect 16968 4361 16974 4395
rect 17008 4361 17014 4395
rect 16968 4323 17014 4361
rect 16968 4289 16974 4323
rect 17008 4289 17014 4323
rect 16968 4251 17014 4289
rect 16968 4217 16974 4251
rect 17008 4217 17014 4251
rect 16968 4179 17014 4217
rect 16968 4145 16974 4179
rect 17008 4145 17014 4179
rect 16968 4130 17014 4145
rect 17064 5115 17110 5130
rect 17064 5081 17070 5115
rect 17104 5081 17110 5115
rect 17064 5043 17110 5081
rect 17064 5009 17070 5043
rect 17104 5009 17110 5043
rect 17064 4971 17110 5009
rect 17064 4937 17070 4971
rect 17104 4937 17110 4971
rect 17064 4899 17110 4937
rect 17064 4865 17070 4899
rect 17104 4865 17110 4899
rect 17064 4827 17110 4865
rect 17064 4793 17070 4827
rect 17104 4793 17110 4827
rect 17064 4755 17110 4793
rect 17064 4721 17070 4755
rect 17104 4721 17110 4755
rect 17064 4683 17110 4721
rect 17064 4649 17070 4683
rect 17104 4649 17110 4683
rect 17064 4611 17110 4649
rect 17064 4577 17070 4611
rect 17104 4577 17110 4611
rect 17064 4539 17110 4577
rect 17064 4505 17070 4539
rect 17104 4505 17110 4539
rect 17064 4467 17110 4505
rect 17064 4433 17070 4467
rect 17104 4433 17110 4467
rect 17064 4395 17110 4433
rect 17064 4361 17070 4395
rect 17104 4361 17110 4395
rect 17064 4323 17110 4361
rect 17064 4289 17070 4323
rect 17104 4289 17110 4323
rect 17064 4251 17110 4289
rect 17064 4217 17070 4251
rect 17104 4217 17110 4251
rect 17064 4179 17110 4217
rect 17064 4145 17070 4179
rect 17104 4145 17110 4179
rect 17064 4130 17110 4145
rect 17160 5115 17206 5130
rect 17160 5081 17166 5115
rect 17200 5081 17206 5115
rect 17160 5043 17206 5081
rect 17160 5009 17166 5043
rect 17200 5009 17206 5043
rect 17160 4971 17206 5009
rect 17160 4937 17166 4971
rect 17200 4937 17206 4971
rect 17160 4899 17206 4937
rect 17160 4865 17166 4899
rect 17200 4865 17206 4899
rect 17160 4827 17206 4865
rect 17160 4793 17166 4827
rect 17200 4793 17206 4827
rect 17160 4755 17206 4793
rect 17160 4721 17166 4755
rect 17200 4721 17206 4755
rect 17160 4683 17206 4721
rect 17160 4649 17166 4683
rect 17200 4649 17206 4683
rect 17160 4611 17206 4649
rect 17160 4577 17166 4611
rect 17200 4577 17206 4611
rect 17160 4539 17206 4577
rect 17160 4505 17166 4539
rect 17200 4505 17206 4539
rect 17160 4467 17206 4505
rect 17160 4433 17166 4467
rect 17200 4433 17206 4467
rect 17160 4395 17206 4433
rect 17160 4361 17166 4395
rect 17200 4361 17206 4395
rect 17160 4323 17206 4361
rect 17160 4289 17166 4323
rect 17200 4289 17206 4323
rect 17160 4251 17206 4289
rect 17160 4217 17166 4251
rect 17200 4217 17206 4251
rect 17160 4179 17206 4217
rect 17160 4145 17166 4179
rect 17200 4145 17206 4179
rect 17160 4130 17206 4145
rect 17256 5115 17302 5130
rect 17256 5081 17262 5115
rect 17296 5081 17302 5115
rect 17256 5043 17302 5081
rect 17256 5009 17262 5043
rect 17296 5009 17302 5043
rect 17256 4971 17302 5009
rect 17256 4937 17262 4971
rect 17296 4937 17302 4971
rect 17256 4899 17302 4937
rect 17256 4865 17262 4899
rect 17296 4865 17302 4899
rect 17256 4827 17302 4865
rect 17256 4793 17262 4827
rect 17296 4793 17302 4827
rect 17256 4755 17302 4793
rect 17256 4721 17262 4755
rect 17296 4721 17302 4755
rect 17256 4683 17302 4721
rect 17256 4649 17262 4683
rect 17296 4649 17302 4683
rect 17256 4611 17302 4649
rect 17256 4577 17262 4611
rect 17296 4577 17302 4611
rect 17256 4539 17302 4577
rect 17256 4505 17262 4539
rect 17296 4505 17302 4539
rect 17256 4467 17302 4505
rect 17256 4433 17262 4467
rect 17296 4433 17302 4467
rect 17256 4395 17302 4433
rect 17256 4361 17262 4395
rect 17296 4361 17302 4395
rect 17256 4323 17302 4361
rect 17256 4289 17262 4323
rect 17296 4289 17302 4323
rect 17256 4251 17302 4289
rect 17256 4217 17262 4251
rect 17296 4217 17302 4251
rect 17256 4179 17302 4217
rect 17256 4145 17262 4179
rect 17296 4145 17302 4179
rect 17256 4130 17302 4145
rect 17464 5113 17510 5128
rect 17464 5079 17470 5113
rect 17504 5079 17510 5113
rect 17464 5041 17510 5079
rect 17464 5007 17470 5041
rect 17504 5007 17510 5041
rect 17464 4969 17510 5007
rect 17464 4935 17470 4969
rect 17504 4935 17510 4969
rect 17464 4897 17510 4935
rect 17464 4863 17470 4897
rect 17504 4863 17510 4897
rect 17464 4825 17510 4863
rect 17464 4791 17470 4825
rect 17504 4791 17510 4825
rect 17464 4753 17510 4791
rect 17464 4719 17470 4753
rect 17504 4719 17510 4753
rect 17464 4681 17510 4719
rect 17464 4647 17470 4681
rect 17504 4647 17510 4681
rect 17464 4609 17510 4647
rect 17464 4575 17470 4609
rect 17504 4575 17510 4609
rect 17464 4537 17510 4575
rect 17464 4503 17470 4537
rect 17504 4503 17510 4537
rect 17464 4465 17510 4503
rect 17464 4431 17470 4465
rect 17504 4431 17510 4465
rect 17464 4393 17510 4431
rect 17464 4359 17470 4393
rect 17504 4359 17510 4393
rect 17464 4321 17510 4359
rect 17464 4287 17470 4321
rect 17504 4287 17510 4321
rect 17464 4249 17510 4287
rect 17464 4215 17470 4249
rect 17504 4215 17510 4249
rect 17464 4177 17510 4215
rect 17464 4143 17470 4177
rect 17504 4143 17510 4177
rect 17464 4128 17510 4143
rect 17560 5113 17606 5128
rect 17560 5079 17566 5113
rect 17600 5079 17606 5113
rect 17560 5041 17606 5079
rect 17560 5007 17566 5041
rect 17600 5007 17606 5041
rect 17560 4969 17606 5007
rect 17560 4935 17566 4969
rect 17600 4935 17606 4969
rect 17560 4897 17606 4935
rect 17560 4863 17566 4897
rect 17600 4863 17606 4897
rect 17560 4825 17606 4863
rect 17560 4791 17566 4825
rect 17600 4791 17606 4825
rect 17560 4753 17606 4791
rect 17560 4719 17566 4753
rect 17600 4719 17606 4753
rect 17560 4681 17606 4719
rect 17560 4647 17566 4681
rect 17600 4647 17606 4681
rect 17560 4609 17606 4647
rect 17560 4575 17566 4609
rect 17600 4575 17606 4609
rect 17560 4537 17606 4575
rect 17560 4503 17566 4537
rect 17600 4503 17606 4537
rect 17560 4465 17606 4503
rect 17560 4431 17566 4465
rect 17600 4431 17606 4465
rect 17560 4393 17606 4431
rect 17560 4359 17566 4393
rect 17600 4359 17606 4393
rect 17560 4321 17606 4359
rect 17560 4287 17566 4321
rect 17600 4287 17606 4321
rect 17560 4249 17606 4287
rect 17560 4215 17566 4249
rect 17600 4215 17606 4249
rect 17560 4177 17606 4215
rect 17560 4143 17566 4177
rect 17600 4143 17606 4177
rect 17560 4128 17606 4143
rect 17656 5113 17702 5128
rect 17656 5079 17662 5113
rect 17696 5079 17702 5113
rect 17656 5041 17702 5079
rect 17656 5007 17662 5041
rect 17696 5007 17702 5041
rect 17656 4969 17702 5007
rect 17656 4935 17662 4969
rect 17696 4935 17702 4969
rect 17656 4897 17702 4935
rect 17656 4863 17662 4897
rect 17696 4863 17702 4897
rect 17656 4825 17702 4863
rect 17656 4791 17662 4825
rect 17696 4791 17702 4825
rect 17656 4753 17702 4791
rect 17656 4719 17662 4753
rect 17696 4719 17702 4753
rect 17656 4681 17702 4719
rect 17656 4647 17662 4681
rect 17696 4647 17702 4681
rect 17656 4609 17702 4647
rect 17656 4575 17662 4609
rect 17696 4575 17702 4609
rect 17656 4537 17702 4575
rect 17656 4503 17662 4537
rect 17696 4503 17702 4537
rect 17656 4465 17702 4503
rect 17656 4431 17662 4465
rect 17696 4431 17702 4465
rect 17656 4393 17702 4431
rect 17656 4359 17662 4393
rect 17696 4359 17702 4393
rect 17656 4321 17702 4359
rect 17656 4287 17662 4321
rect 17696 4287 17702 4321
rect 17656 4249 17702 4287
rect 17656 4215 17662 4249
rect 17696 4215 17702 4249
rect 17656 4177 17702 4215
rect 17656 4143 17662 4177
rect 17696 4143 17702 4177
rect 17656 4128 17702 4143
rect 17752 5113 17798 5128
rect 17752 5079 17758 5113
rect 17792 5079 17798 5113
rect 17752 5041 17798 5079
rect 17752 5007 17758 5041
rect 17792 5007 17798 5041
rect 17752 4969 17798 5007
rect 17752 4935 17758 4969
rect 17792 4935 17798 4969
rect 17752 4897 17798 4935
rect 17752 4863 17758 4897
rect 17792 4863 17798 4897
rect 17752 4825 17798 4863
rect 17752 4791 17758 4825
rect 17792 4791 17798 4825
rect 17752 4753 17798 4791
rect 17752 4719 17758 4753
rect 17792 4719 17798 4753
rect 17752 4681 17798 4719
rect 17752 4647 17758 4681
rect 17792 4647 17798 4681
rect 17752 4609 17798 4647
rect 17752 4575 17758 4609
rect 17792 4575 17798 4609
rect 17752 4537 17798 4575
rect 17752 4503 17758 4537
rect 17792 4503 17798 4537
rect 17752 4465 17798 4503
rect 17752 4431 17758 4465
rect 17792 4431 17798 4465
rect 17752 4393 17798 4431
rect 17752 4359 17758 4393
rect 17792 4359 17798 4393
rect 17752 4321 17798 4359
rect 17752 4287 17758 4321
rect 17792 4287 17798 4321
rect 17752 4249 17798 4287
rect 17752 4215 17758 4249
rect 17792 4215 17798 4249
rect 17752 4177 17798 4215
rect 17752 4143 17758 4177
rect 17792 4143 17798 4177
rect 17752 4128 17798 4143
rect 17848 5113 17894 5128
rect 17848 5079 17854 5113
rect 17888 5079 17894 5113
rect 17848 5041 17894 5079
rect 17848 5007 17854 5041
rect 17888 5007 17894 5041
rect 17848 4969 17894 5007
rect 17848 4935 17854 4969
rect 17888 4935 17894 4969
rect 17848 4897 17894 4935
rect 17848 4863 17854 4897
rect 17888 4863 17894 4897
rect 17848 4825 17894 4863
rect 17848 4791 17854 4825
rect 17888 4791 17894 4825
rect 17848 4753 17894 4791
rect 17848 4719 17854 4753
rect 17888 4719 17894 4753
rect 17848 4681 17894 4719
rect 17848 4647 17854 4681
rect 17888 4647 17894 4681
rect 17848 4609 17894 4647
rect 17848 4575 17854 4609
rect 17888 4575 17894 4609
rect 17848 4537 17894 4575
rect 17848 4503 17854 4537
rect 17888 4503 17894 4537
rect 17848 4465 17894 4503
rect 17848 4431 17854 4465
rect 17888 4431 17894 4465
rect 17848 4393 17894 4431
rect 17848 4359 17854 4393
rect 17888 4359 17894 4393
rect 17848 4321 17894 4359
rect 17848 4287 17854 4321
rect 17888 4287 17894 4321
rect 17848 4249 17894 4287
rect 17848 4215 17854 4249
rect 17888 4215 17894 4249
rect 17848 4177 17894 4215
rect 17848 4143 17854 4177
rect 17888 4143 17894 4177
rect 17848 4128 17894 4143
rect 17944 5113 17990 5128
rect 17944 5079 17950 5113
rect 17984 5079 17990 5113
rect 17944 5041 17990 5079
rect 17944 5007 17950 5041
rect 17984 5007 17990 5041
rect 17944 4969 17990 5007
rect 17944 4935 17950 4969
rect 17984 4935 17990 4969
rect 17944 4897 17990 4935
rect 17944 4863 17950 4897
rect 17984 4863 17990 4897
rect 17944 4825 17990 4863
rect 17944 4791 17950 4825
rect 17984 4791 17990 4825
rect 17944 4753 17990 4791
rect 17944 4719 17950 4753
rect 17984 4719 17990 4753
rect 17944 4681 17990 4719
rect 17944 4647 17950 4681
rect 17984 4647 17990 4681
rect 17944 4609 17990 4647
rect 17944 4575 17950 4609
rect 17984 4575 17990 4609
rect 17944 4537 17990 4575
rect 17944 4503 17950 4537
rect 17984 4503 17990 4537
rect 17944 4465 17990 4503
rect 17944 4431 17950 4465
rect 17984 4431 17990 4465
rect 17944 4393 17990 4431
rect 17944 4359 17950 4393
rect 17984 4359 17990 4393
rect 17944 4321 17990 4359
rect 17944 4287 17950 4321
rect 17984 4287 17990 4321
rect 17944 4249 17990 4287
rect 17944 4215 17950 4249
rect 17984 4215 17990 4249
rect 17944 4177 17990 4215
rect 17944 4143 17950 4177
rect 17984 4143 17990 4177
rect 17944 4128 17990 4143
rect 18040 5113 18086 5128
rect 18040 5079 18046 5113
rect 18080 5079 18086 5113
rect 18040 5041 18086 5079
rect 18040 5007 18046 5041
rect 18080 5007 18086 5041
rect 18040 4969 18086 5007
rect 18040 4935 18046 4969
rect 18080 4935 18086 4969
rect 18040 4897 18086 4935
rect 18040 4863 18046 4897
rect 18080 4863 18086 4897
rect 18040 4825 18086 4863
rect 18040 4791 18046 4825
rect 18080 4791 18086 4825
rect 18040 4753 18086 4791
rect 18040 4719 18046 4753
rect 18080 4719 18086 4753
rect 18040 4681 18086 4719
rect 18040 4647 18046 4681
rect 18080 4647 18086 4681
rect 18040 4609 18086 4647
rect 18040 4575 18046 4609
rect 18080 4575 18086 4609
rect 18040 4537 18086 4575
rect 18040 4503 18046 4537
rect 18080 4503 18086 4537
rect 18040 4465 18086 4503
rect 18040 4431 18046 4465
rect 18080 4431 18086 4465
rect 18040 4393 18086 4431
rect 18040 4359 18046 4393
rect 18080 4359 18086 4393
rect 18040 4321 18086 4359
rect 18040 4287 18046 4321
rect 18080 4287 18086 4321
rect 18040 4249 18086 4287
rect 18040 4215 18046 4249
rect 18080 4215 18086 4249
rect 18040 4177 18086 4215
rect 18040 4143 18046 4177
rect 18080 4143 18086 4177
rect 18040 4128 18086 4143
rect 18136 5113 18182 5128
rect 18136 5079 18142 5113
rect 18176 5079 18182 5113
rect 18136 5041 18182 5079
rect 18136 5007 18142 5041
rect 18176 5007 18182 5041
rect 18136 4969 18182 5007
rect 18136 4935 18142 4969
rect 18176 4935 18182 4969
rect 18136 4897 18182 4935
rect 18136 4863 18142 4897
rect 18176 4863 18182 4897
rect 18136 4825 18182 4863
rect 18136 4791 18142 4825
rect 18176 4791 18182 4825
rect 18136 4753 18182 4791
rect 18136 4719 18142 4753
rect 18176 4719 18182 4753
rect 18136 4681 18182 4719
rect 18136 4647 18142 4681
rect 18176 4647 18182 4681
rect 18136 4609 18182 4647
rect 18136 4575 18142 4609
rect 18176 4575 18182 4609
rect 18136 4537 18182 4575
rect 18136 4503 18142 4537
rect 18176 4503 18182 4537
rect 18136 4465 18182 4503
rect 18136 4431 18142 4465
rect 18176 4431 18182 4465
rect 18136 4393 18182 4431
rect 18136 4359 18142 4393
rect 18176 4359 18182 4393
rect 18136 4321 18182 4359
rect 18136 4287 18142 4321
rect 18176 4287 18182 4321
rect 18136 4249 18182 4287
rect 18136 4215 18142 4249
rect 18176 4215 18182 4249
rect 18136 4177 18182 4215
rect 18136 4143 18142 4177
rect 18176 4143 18182 4177
rect 18136 4128 18182 4143
rect 18232 5113 18278 5128
rect 18232 5079 18238 5113
rect 18272 5079 18278 5113
rect 18232 5041 18278 5079
rect 18232 5007 18238 5041
rect 18272 5007 18278 5041
rect 18232 4969 18278 5007
rect 18232 4935 18238 4969
rect 18272 4935 18278 4969
rect 18232 4897 18278 4935
rect 18232 4863 18238 4897
rect 18272 4863 18278 4897
rect 18232 4825 18278 4863
rect 18232 4791 18238 4825
rect 18272 4791 18278 4825
rect 18232 4753 18278 4791
rect 18232 4719 18238 4753
rect 18272 4719 18278 4753
rect 18232 4681 18278 4719
rect 18232 4647 18238 4681
rect 18272 4647 18278 4681
rect 18232 4609 18278 4647
rect 18232 4575 18238 4609
rect 18272 4575 18278 4609
rect 18232 4537 18278 4575
rect 18232 4503 18238 4537
rect 18272 4503 18278 4537
rect 18232 4465 18278 4503
rect 18232 4431 18238 4465
rect 18272 4431 18278 4465
rect 18232 4393 18278 4431
rect 18232 4359 18238 4393
rect 18272 4359 18278 4393
rect 18232 4321 18278 4359
rect 18232 4287 18238 4321
rect 18272 4287 18278 4321
rect 18232 4249 18278 4287
rect 18232 4215 18238 4249
rect 18272 4215 18278 4249
rect 18232 4177 18278 4215
rect 18232 4143 18238 4177
rect 18272 4143 18278 4177
rect 18232 4128 18278 4143
rect 18328 5113 18374 5128
rect 18328 5079 18334 5113
rect 18368 5079 18374 5113
rect 18328 5041 18374 5079
rect 18328 5007 18334 5041
rect 18368 5007 18374 5041
rect 18328 4969 18374 5007
rect 18328 4935 18334 4969
rect 18368 4935 18374 4969
rect 18328 4897 18374 4935
rect 18328 4863 18334 4897
rect 18368 4863 18374 4897
rect 18328 4825 18374 4863
rect 18328 4791 18334 4825
rect 18368 4791 18374 4825
rect 18328 4753 18374 4791
rect 18328 4719 18334 4753
rect 18368 4719 18374 4753
rect 18328 4681 18374 4719
rect 18328 4647 18334 4681
rect 18368 4647 18374 4681
rect 18328 4609 18374 4647
rect 18328 4575 18334 4609
rect 18368 4575 18374 4609
rect 18328 4537 18374 4575
rect 18328 4503 18334 4537
rect 18368 4503 18374 4537
rect 18328 4465 18374 4503
rect 18328 4431 18334 4465
rect 18368 4431 18374 4465
rect 18328 4393 18374 4431
rect 18328 4359 18334 4393
rect 18368 4359 18374 4393
rect 18328 4321 18374 4359
rect 18328 4287 18334 4321
rect 18368 4287 18374 4321
rect 18328 4249 18374 4287
rect 18328 4215 18334 4249
rect 18368 4215 18374 4249
rect 18328 4177 18374 4215
rect 18328 4143 18334 4177
rect 18368 4143 18374 4177
rect 18328 4128 18374 4143
rect 18424 5113 18470 5128
rect 18424 5079 18430 5113
rect 18464 5079 18470 5113
rect 18424 5041 18470 5079
rect 18424 5007 18430 5041
rect 18464 5007 18470 5041
rect 18424 4969 18470 5007
rect 18424 4935 18430 4969
rect 18464 4935 18470 4969
rect 18424 4897 18470 4935
rect 18424 4863 18430 4897
rect 18464 4863 18470 4897
rect 18424 4825 18470 4863
rect 18424 4791 18430 4825
rect 18464 4791 18470 4825
rect 18424 4753 18470 4791
rect 18424 4719 18430 4753
rect 18464 4719 18470 4753
rect 18424 4681 18470 4719
rect 18424 4647 18430 4681
rect 18464 4647 18470 4681
rect 18424 4609 18470 4647
rect 18424 4575 18430 4609
rect 18464 4575 18470 4609
rect 18424 4537 18470 4575
rect 18424 4503 18430 4537
rect 18464 4503 18470 4537
rect 18424 4465 18470 4503
rect 18424 4431 18430 4465
rect 18464 4431 18470 4465
rect 18424 4393 18470 4431
rect 18424 4359 18430 4393
rect 18464 4359 18470 4393
rect 18424 4321 18470 4359
rect 18424 4287 18430 4321
rect 18464 4287 18470 4321
rect 18424 4249 18470 4287
rect 18424 4215 18430 4249
rect 18464 4215 18470 4249
rect 18424 4177 18470 4215
rect 18424 4143 18430 4177
rect 18464 4143 18470 4177
rect 18424 4128 18470 4143
rect 18668 5107 18714 5122
rect 18668 5073 18674 5107
rect 18708 5073 18714 5107
rect 18668 5035 18714 5073
rect 18668 5001 18674 5035
rect 18708 5001 18714 5035
rect 18668 4963 18714 5001
rect 18668 4929 18674 4963
rect 18708 4929 18714 4963
rect 18668 4891 18714 4929
rect 18668 4857 18674 4891
rect 18708 4857 18714 4891
rect 18668 4819 18714 4857
rect 18668 4785 18674 4819
rect 18708 4785 18714 4819
rect 18668 4747 18714 4785
rect 18668 4713 18674 4747
rect 18708 4713 18714 4747
rect 18668 4675 18714 4713
rect 18668 4641 18674 4675
rect 18708 4641 18714 4675
rect 18668 4603 18714 4641
rect 18668 4569 18674 4603
rect 18708 4569 18714 4603
rect 18668 4531 18714 4569
rect 18668 4497 18674 4531
rect 18708 4497 18714 4531
rect 18668 4459 18714 4497
rect 18668 4425 18674 4459
rect 18708 4425 18714 4459
rect 18668 4387 18714 4425
rect 18668 4353 18674 4387
rect 18708 4353 18714 4387
rect 18668 4315 18714 4353
rect 18668 4281 18674 4315
rect 18708 4281 18714 4315
rect 18668 4243 18714 4281
rect 18668 4209 18674 4243
rect 18708 4209 18714 4243
rect 18668 4171 18714 4209
rect 18668 4137 18674 4171
rect 18708 4137 18714 4171
rect 18668 4122 18714 4137
rect 18764 5107 18810 5122
rect 18764 5073 18770 5107
rect 18804 5073 18810 5107
rect 18764 5035 18810 5073
rect 18764 5001 18770 5035
rect 18804 5001 18810 5035
rect 18764 4963 18810 5001
rect 18764 4929 18770 4963
rect 18804 4929 18810 4963
rect 18764 4891 18810 4929
rect 18764 4857 18770 4891
rect 18804 4857 18810 4891
rect 18764 4819 18810 4857
rect 18764 4785 18770 4819
rect 18804 4785 18810 4819
rect 18764 4747 18810 4785
rect 18764 4713 18770 4747
rect 18804 4713 18810 4747
rect 18764 4675 18810 4713
rect 18764 4641 18770 4675
rect 18804 4641 18810 4675
rect 18764 4603 18810 4641
rect 18764 4569 18770 4603
rect 18804 4569 18810 4603
rect 18764 4531 18810 4569
rect 18764 4497 18770 4531
rect 18804 4497 18810 4531
rect 18764 4459 18810 4497
rect 18764 4425 18770 4459
rect 18804 4425 18810 4459
rect 18764 4387 18810 4425
rect 18764 4353 18770 4387
rect 18804 4353 18810 4387
rect 18764 4315 18810 4353
rect 18764 4281 18770 4315
rect 18804 4281 18810 4315
rect 18764 4243 18810 4281
rect 18764 4209 18770 4243
rect 18804 4209 18810 4243
rect 18764 4171 18810 4209
rect 18764 4137 18770 4171
rect 18804 4137 18810 4171
rect 18764 4122 18810 4137
rect 18860 5107 18906 5122
rect 18860 5073 18866 5107
rect 18900 5073 18906 5107
rect 18860 5035 18906 5073
rect 18860 5001 18866 5035
rect 18900 5001 18906 5035
rect 18860 4963 18906 5001
rect 18860 4929 18866 4963
rect 18900 4929 18906 4963
rect 18860 4891 18906 4929
rect 18860 4857 18866 4891
rect 18900 4857 18906 4891
rect 18860 4819 18906 4857
rect 18860 4785 18866 4819
rect 18900 4785 18906 4819
rect 18860 4747 18906 4785
rect 18860 4713 18866 4747
rect 18900 4713 18906 4747
rect 18860 4675 18906 4713
rect 18860 4641 18866 4675
rect 18900 4641 18906 4675
rect 18860 4603 18906 4641
rect 18860 4569 18866 4603
rect 18900 4569 18906 4603
rect 18860 4531 18906 4569
rect 18860 4497 18866 4531
rect 18900 4497 18906 4531
rect 18860 4459 18906 4497
rect 18860 4425 18866 4459
rect 18900 4425 18906 4459
rect 18860 4387 18906 4425
rect 18860 4353 18866 4387
rect 18900 4353 18906 4387
rect 18860 4315 18906 4353
rect 18860 4281 18866 4315
rect 18900 4281 18906 4315
rect 18860 4243 18906 4281
rect 18860 4209 18866 4243
rect 18900 4209 18906 4243
rect 18860 4171 18906 4209
rect 18860 4137 18866 4171
rect 18900 4137 18906 4171
rect 18860 4122 18906 4137
rect 18956 5107 19002 5122
rect 18956 5073 18962 5107
rect 18996 5073 19002 5107
rect 18956 5035 19002 5073
rect 18956 5001 18962 5035
rect 18996 5001 19002 5035
rect 18956 4963 19002 5001
rect 18956 4929 18962 4963
rect 18996 4929 19002 4963
rect 18956 4891 19002 4929
rect 18956 4857 18962 4891
rect 18996 4857 19002 4891
rect 18956 4819 19002 4857
rect 18956 4785 18962 4819
rect 18996 4785 19002 4819
rect 18956 4747 19002 4785
rect 18956 4713 18962 4747
rect 18996 4713 19002 4747
rect 18956 4675 19002 4713
rect 18956 4641 18962 4675
rect 18996 4641 19002 4675
rect 18956 4603 19002 4641
rect 18956 4569 18962 4603
rect 18996 4569 19002 4603
rect 18956 4531 19002 4569
rect 18956 4497 18962 4531
rect 18996 4497 19002 4531
rect 18956 4459 19002 4497
rect 18956 4425 18962 4459
rect 18996 4425 19002 4459
rect 18956 4387 19002 4425
rect 18956 4353 18962 4387
rect 18996 4353 19002 4387
rect 18956 4315 19002 4353
rect 18956 4281 18962 4315
rect 18996 4281 19002 4315
rect 18956 4243 19002 4281
rect 18956 4209 18962 4243
rect 18996 4209 19002 4243
rect 18956 4171 19002 4209
rect 18956 4137 18962 4171
rect 18996 4137 19002 4171
rect 18956 4122 19002 4137
rect 19052 5107 19098 5122
rect 19052 5073 19058 5107
rect 19092 5073 19098 5107
rect 19052 5035 19098 5073
rect 19052 5001 19058 5035
rect 19092 5001 19098 5035
rect 19052 4963 19098 5001
rect 19052 4929 19058 4963
rect 19092 4929 19098 4963
rect 19052 4891 19098 4929
rect 19052 4857 19058 4891
rect 19092 4857 19098 4891
rect 19052 4819 19098 4857
rect 19052 4785 19058 4819
rect 19092 4785 19098 4819
rect 19052 4747 19098 4785
rect 19052 4713 19058 4747
rect 19092 4713 19098 4747
rect 19052 4675 19098 4713
rect 19052 4641 19058 4675
rect 19092 4641 19098 4675
rect 19052 4603 19098 4641
rect 19052 4569 19058 4603
rect 19092 4569 19098 4603
rect 19052 4531 19098 4569
rect 19052 4497 19058 4531
rect 19092 4497 19098 4531
rect 19052 4459 19098 4497
rect 19052 4425 19058 4459
rect 19092 4425 19098 4459
rect 19052 4387 19098 4425
rect 19052 4353 19058 4387
rect 19092 4353 19098 4387
rect 19052 4315 19098 4353
rect 19052 4281 19058 4315
rect 19092 4281 19098 4315
rect 19052 4243 19098 4281
rect 19052 4209 19058 4243
rect 19092 4209 19098 4243
rect 19052 4171 19098 4209
rect 19052 4137 19058 4171
rect 19092 4137 19098 4171
rect 19052 4122 19098 4137
rect 19148 5107 19194 5122
rect 19148 5073 19154 5107
rect 19188 5073 19194 5107
rect 19148 5035 19194 5073
rect 19148 5001 19154 5035
rect 19188 5001 19194 5035
rect 19148 4963 19194 5001
rect 19148 4929 19154 4963
rect 19188 4929 19194 4963
rect 19148 4891 19194 4929
rect 19148 4857 19154 4891
rect 19188 4857 19194 4891
rect 19148 4819 19194 4857
rect 19148 4785 19154 4819
rect 19188 4785 19194 4819
rect 19148 4747 19194 4785
rect 19148 4713 19154 4747
rect 19188 4713 19194 4747
rect 19148 4675 19194 4713
rect 19148 4641 19154 4675
rect 19188 4641 19194 4675
rect 19148 4603 19194 4641
rect 19148 4569 19154 4603
rect 19188 4569 19194 4603
rect 19148 4531 19194 4569
rect 19148 4497 19154 4531
rect 19188 4497 19194 4531
rect 19148 4459 19194 4497
rect 19148 4425 19154 4459
rect 19188 4425 19194 4459
rect 19148 4387 19194 4425
rect 19148 4353 19154 4387
rect 19188 4353 19194 4387
rect 19148 4315 19194 4353
rect 19148 4281 19154 4315
rect 19188 4281 19194 4315
rect 19148 4243 19194 4281
rect 19148 4209 19154 4243
rect 19188 4209 19194 4243
rect 19148 4171 19194 4209
rect 19148 4137 19154 4171
rect 19188 4137 19194 4171
rect 19148 4122 19194 4137
rect 19244 5107 19290 5122
rect 19244 5073 19250 5107
rect 19284 5073 19290 5107
rect 19244 5035 19290 5073
rect 19244 5001 19250 5035
rect 19284 5001 19290 5035
rect 19244 4963 19290 5001
rect 19244 4929 19250 4963
rect 19284 4929 19290 4963
rect 19244 4891 19290 4929
rect 19244 4857 19250 4891
rect 19284 4857 19290 4891
rect 19244 4819 19290 4857
rect 19244 4785 19250 4819
rect 19284 4785 19290 4819
rect 19244 4747 19290 4785
rect 19244 4713 19250 4747
rect 19284 4713 19290 4747
rect 19244 4675 19290 4713
rect 19244 4641 19250 4675
rect 19284 4641 19290 4675
rect 19244 4603 19290 4641
rect 19244 4569 19250 4603
rect 19284 4569 19290 4603
rect 19244 4531 19290 4569
rect 19244 4497 19250 4531
rect 19284 4497 19290 4531
rect 19244 4459 19290 4497
rect 19244 4425 19250 4459
rect 19284 4425 19290 4459
rect 19244 4387 19290 4425
rect 19244 4353 19250 4387
rect 19284 4353 19290 4387
rect 19244 4315 19290 4353
rect 19244 4281 19250 4315
rect 19284 4281 19290 4315
rect 19244 4243 19290 4281
rect 19244 4209 19250 4243
rect 19284 4209 19290 4243
rect 19244 4171 19290 4209
rect 19244 4137 19250 4171
rect 19284 4137 19290 4171
rect 19244 4122 19290 4137
rect 19340 5107 19386 5122
rect 19340 5073 19346 5107
rect 19380 5073 19386 5107
rect 19340 5035 19386 5073
rect 19340 5001 19346 5035
rect 19380 5001 19386 5035
rect 19340 4963 19386 5001
rect 19340 4929 19346 4963
rect 19380 4929 19386 4963
rect 19340 4891 19386 4929
rect 19340 4857 19346 4891
rect 19380 4857 19386 4891
rect 19340 4819 19386 4857
rect 19340 4785 19346 4819
rect 19380 4785 19386 4819
rect 19340 4747 19386 4785
rect 19340 4713 19346 4747
rect 19380 4713 19386 4747
rect 19340 4675 19386 4713
rect 19340 4641 19346 4675
rect 19380 4641 19386 4675
rect 19340 4603 19386 4641
rect 19340 4569 19346 4603
rect 19380 4569 19386 4603
rect 19340 4531 19386 4569
rect 19340 4497 19346 4531
rect 19380 4497 19386 4531
rect 19340 4459 19386 4497
rect 19340 4425 19346 4459
rect 19380 4425 19386 4459
rect 19340 4387 19386 4425
rect 19340 4353 19346 4387
rect 19380 4353 19386 4387
rect 19340 4315 19386 4353
rect 19340 4281 19346 4315
rect 19380 4281 19386 4315
rect 19340 4243 19386 4281
rect 19340 4209 19346 4243
rect 19380 4209 19386 4243
rect 19340 4171 19386 4209
rect 19340 4137 19346 4171
rect 19380 4137 19386 4171
rect 19340 4122 19386 4137
rect 19436 5107 19482 5122
rect 19436 5073 19442 5107
rect 19476 5073 19482 5107
rect 19436 5035 19482 5073
rect 19436 5001 19442 5035
rect 19476 5001 19482 5035
rect 19436 4963 19482 5001
rect 19436 4929 19442 4963
rect 19476 4929 19482 4963
rect 19436 4891 19482 4929
rect 19436 4857 19442 4891
rect 19476 4857 19482 4891
rect 19436 4819 19482 4857
rect 19436 4785 19442 4819
rect 19476 4785 19482 4819
rect 19436 4747 19482 4785
rect 19436 4713 19442 4747
rect 19476 4713 19482 4747
rect 19436 4675 19482 4713
rect 19436 4641 19442 4675
rect 19476 4641 19482 4675
rect 19436 4603 19482 4641
rect 19436 4569 19442 4603
rect 19476 4569 19482 4603
rect 19436 4531 19482 4569
rect 19436 4497 19442 4531
rect 19476 4497 19482 4531
rect 19436 4459 19482 4497
rect 19436 4425 19442 4459
rect 19476 4425 19482 4459
rect 19436 4387 19482 4425
rect 19436 4353 19442 4387
rect 19476 4353 19482 4387
rect 19436 4315 19482 4353
rect 19436 4281 19442 4315
rect 19476 4281 19482 4315
rect 19436 4243 19482 4281
rect 19436 4209 19442 4243
rect 19476 4209 19482 4243
rect 19436 4171 19482 4209
rect 19436 4137 19442 4171
rect 19476 4137 19482 4171
rect 19436 4122 19482 4137
rect 19532 5107 19578 5122
rect 19532 5073 19538 5107
rect 19572 5073 19578 5107
rect 19532 5035 19578 5073
rect 19532 5001 19538 5035
rect 19572 5001 19578 5035
rect 19532 4963 19578 5001
rect 19532 4929 19538 4963
rect 19572 4929 19578 4963
rect 19532 4891 19578 4929
rect 19532 4857 19538 4891
rect 19572 4857 19578 4891
rect 19532 4819 19578 4857
rect 19532 4785 19538 4819
rect 19572 4785 19578 4819
rect 19532 4747 19578 4785
rect 19532 4713 19538 4747
rect 19572 4713 19578 4747
rect 19532 4675 19578 4713
rect 19532 4641 19538 4675
rect 19572 4641 19578 4675
rect 19532 4603 19578 4641
rect 19532 4569 19538 4603
rect 19572 4569 19578 4603
rect 19532 4531 19578 4569
rect 19532 4497 19538 4531
rect 19572 4497 19578 4531
rect 19532 4459 19578 4497
rect 19532 4425 19538 4459
rect 19572 4425 19578 4459
rect 19532 4387 19578 4425
rect 19532 4353 19538 4387
rect 19572 4353 19578 4387
rect 19532 4315 19578 4353
rect 19532 4281 19538 4315
rect 19572 4281 19578 4315
rect 19532 4243 19578 4281
rect 19532 4209 19538 4243
rect 19572 4209 19578 4243
rect 19532 4171 19578 4209
rect 19532 4137 19538 4171
rect 19572 4137 19578 4171
rect 19532 4122 19578 4137
rect 19628 5107 19674 5122
rect 19628 5073 19634 5107
rect 19668 5073 19674 5107
rect 19628 5035 19674 5073
rect 19628 5001 19634 5035
rect 19668 5001 19674 5035
rect 19628 4963 19674 5001
rect 19628 4929 19634 4963
rect 19668 4929 19674 4963
rect 19628 4891 19674 4929
rect 19628 4857 19634 4891
rect 19668 4857 19674 4891
rect 19628 4819 19674 4857
rect 19628 4785 19634 4819
rect 19668 4785 19674 4819
rect 19628 4747 19674 4785
rect 19628 4713 19634 4747
rect 19668 4713 19674 4747
rect 19628 4675 19674 4713
rect 19628 4641 19634 4675
rect 19668 4641 19674 4675
rect 19628 4603 19674 4641
rect 19628 4569 19634 4603
rect 19668 4569 19674 4603
rect 19628 4531 19674 4569
rect 19628 4497 19634 4531
rect 19668 4497 19674 4531
rect 19628 4459 19674 4497
rect 19628 4425 19634 4459
rect 19668 4425 19674 4459
rect 19628 4387 19674 4425
rect 19628 4353 19634 4387
rect 19668 4353 19674 4387
rect 19628 4315 19674 4353
rect 19628 4281 19634 4315
rect 19668 4281 19674 4315
rect 19628 4243 19674 4281
rect 19628 4209 19634 4243
rect 19668 4209 19674 4243
rect 19628 4171 19674 4209
rect 19628 4137 19634 4171
rect 19668 4137 19674 4171
rect 19628 4122 19674 4137
rect 19724 5107 19770 5122
rect 19724 5073 19730 5107
rect 19764 5073 19770 5107
rect 19724 5035 19770 5073
rect 19724 5001 19730 5035
rect 19764 5001 19770 5035
rect 19724 4963 19770 5001
rect 19724 4929 19730 4963
rect 19764 4929 19770 4963
rect 19724 4891 19770 4929
rect 19724 4857 19730 4891
rect 19764 4857 19770 4891
rect 19724 4819 19770 4857
rect 19724 4785 19730 4819
rect 19764 4785 19770 4819
rect 19724 4747 19770 4785
rect 19724 4713 19730 4747
rect 19764 4713 19770 4747
rect 19724 4675 19770 4713
rect 19724 4641 19730 4675
rect 19764 4641 19770 4675
rect 19724 4603 19770 4641
rect 19724 4569 19730 4603
rect 19764 4569 19770 4603
rect 19724 4531 19770 4569
rect 19724 4497 19730 4531
rect 19764 4497 19770 4531
rect 19724 4459 19770 4497
rect 19724 4425 19730 4459
rect 19764 4425 19770 4459
rect 19724 4387 19770 4425
rect 19724 4353 19730 4387
rect 19764 4353 19770 4387
rect 19724 4315 19770 4353
rect 19724 4281 19730 4315
rect 19764 4281 19770 4315
rect 19724 4243 19770 4281
rect 19724 4209 19730 4243
rect 19764 4209 19770 4243
rect 19724 4171 19770 4209
rect 19724 4137 19730 4171
rect 19764 4137 19770 4171
rect 19724 4122 19770 4137
rect 19820 5107 19866 5122
rect 19820 5073 19826 5107
rect 19860 5073 19866 5107
rect 19820 5035 19866 5073
rect 19820 5001 19826 5035
rect 19860 5001 19866 5035
rect 19820 4963 19866 5001
rect 19820 4929 19826 4963
rect 19860 4929 19866 4963
rect 19820 4891 19866 4929
rect 19820 4857 19826 4891
rect 19860 4857 19866 4891
rect 19820 4819 19866 4857
rect 19820 4785 19826 4819
rect 19860 4785 19866 4819
rect 19820 4747 19866 4785
rect 19820 4713 19826 4747
rect 19860 4713 19866 4747
rect 19820 4675 19866 4713
rect 19820 4641 19826 4675
rect 19860 4641 19866 4675
rect 19820 4603 19866 4641
rect 19820 4569 19826 4603
rect 19860 4569 19866 4603
rect 19820 4531 19866 4569
rect 19820 4497 19826 4531
rect 19860 4497 19866 4531
rect 19820 4459 19866 4497
rect 19820 4425 19826 4459
rect 19860 4425 19866 4459
rect 19820 4387 19866 4425
rect 19820 4353 19826 4387
rect 19860 4353 19866 4387
rect 19820 4315 19866 4353
rect 19820 4281 19826 4315
rect 19860 4281 19866 4315
rect 19820 4243 19866 4281
rect 19820 4209 19826 4243
rect 19860 4209 19866 4243
rect 19820 4171 19866 4209
rect 19820 4137 19826 4171
rect 19860 4137 19866 4171
rect 19820 4122 19866 4137
rect 19916 5107 19962 5122
rect 19916 5073 19922 5107
rect 19956 5073 19962 5107
rect 19916 5035 19962 5073
rect 19916 5001 19922 5035
rect 19956 5001 19962 5035
rect 19916 4963 19962 5001
rect 19916 4929 19922 4963
rect 19956 4929 19962 4963
rect 19916 4891 19962 4929
rect 19916 4857 19922 4891
rect 19956 4857 19962 4891
rect 19916 4819 19962 4857
rect 19916 4785 19922 4819
rect 19956 4785 19962 4819
rect 19916 4747 19962 4785
rect 19916 4713 19922 4747
rect 19956 4713 19962 4747
rect 19916 4675 19962 4713
rect 19916 4641 19922 4675
rect 19956 4641 19962 4675
rect 19916 4603 19962 4641
rect 19916 4569 19922 4603
rect 19956 4569 19962 4603
rect 19916 4531 19962 4569
rect 19916 4497 19922 4531
rect 19956 4497 19962 4531
rect 19916 4459 19962 4497
rect 19916 4425 19922 4459
rect 19956 4425 19962 4459
rect 19916 4387 19962 4425
rect 19916 4353 19922 4387
rect 19956 4353 19962 4387
rect 19916 4315 19962 4353
rect 19916 4281 19922 4315
rect 19956 4281 19962 4315
rect 19916 4243 19962 4281
rect 19916 4209 19922 4243
rect 19956 4209 19962 4243
rect 19916 4171 19962 4209
rect 19916 4137 19922 4171
rect 19956 4137 19962 4171
rect 19916 4122 19962 4137
rect 20012 5107 20058 5122
rect 20012 5073 20018 5107
rect 20052 5073 20058 5107
rect 20012 5035 20058 5073
rect 20012 5001 20018 5035
rect 20052 5001 20058 5035
rect 20012 4963 20058 5001
rect 20012 4929 20018 4963
rect 20052 4929 20058 4963
rect 20012 4891 20058 4929
rect 20012 4857 20018 4891
rect 20052 4857 20058 4891
rect 20012 4819 20058 4857
rect 20012 4785 20018 4819
rect 20052 4785 20058 4819
rect 20012 4747 20058 4785
rect 20012 4713 20018 4747
rect 20052 4713 20058 4747
rect 20012 4675 20058 4713
rect 20012 4641 20018 4675
rect 20052 4641 20058 4675
rect 20012 4603 20058 4641
rect 20012 4569 20018 4603
rect 20052 4569 20058 4603
rect 20012 4531 20058 4569
rect 20012 4497 20018 4531
rect 20052 4497 20058 4531
rect 20012 4459 20058 4497
rect 20012 4425 20018 4459
rect 20052 4425 20058 4459
rect 20012 4387 20058 4425
rect 20012 4353 20018 4387
rect 20052 4353 20058 4387
rect 20012 4315 20058 4353
rect 20012 4281 20018 4315
rect 20052 4281 20058 4315
rect 20012 4243 20058 4281
rect 20012 4209 20018 4243
rect 20052 4209 20058 4243
rect 20012 4171 20058 4209
rect 20012 4137 20018 4171
rect 20052 4137 20058 4171
rect 20012 4122 20058 4137
rect 20108 5107 20154 5122
rect 20108 5073 20114 5107
rect 20148 5073 20154 5107
rect 20108 5035 20154 5073
rect 20108 5001 20114 5035
rect 20148 5001 20154 5035
rect 20108 4963 20154 5001
rect 20108 4929 20114 4963
rect 20148 4929 20154 4963
rect 20108 4891 20154 4929
rect 20108 4857 20114 4891
rect 20148 4857 20154 4891
rect 20108 4819 20154 4857
rect 20108 4785 20114 4819
rect 20148 4785 20154 4819
rect 20108 4747 20154 4785
rect 20108 4713 20114 4747
rect 20148 4713 20154 4747
rect 20108 4675 20154 4713
rect 20108 4641 20114 4675
rect 20148 4641 20154 4675
rect 20108 4603 20154 4641
rect 20108 4569 20114 4603
rect 20148 4569 20154 4603
rect 20108 4531 20154 4569
rect 20108 4497 20114 4531
rect 20148 4497 20154 4531
rect 20108 4459 20154 4497
rect 20108 4425 20114 4459
rect 20148 4425 20154 4459
rect 20108 4387 20154 4425
rect 20108 4353 20114 4387
rect 20148 4353 20154 4387
rect 20108 4315 20154 4353
rect 20108 4281 20114 4315
rect 20148 4281 20154 4315
rect 20108 4243 20154 4281
rect 20108 4209 20114 4243
rect 20148 4209 20154 4243
rect 20108 4171 20154 4209
rect 20108 4137 20114 4171
rect 20148 4137 20154 4171
rect 20108 4122 20154 4137
rect 20332 5101 20378 5116
rect 20332 5067 20338 5101
rect 20372 5067 20378 5101
rect 20332 5029 20378 5067
rect 20332 4995 20338 5029
rect 20372 4995 20378 5029
rect 20332 4957 20378 4995
rect 20332 4923 20338 4957
rect 20372 4923 20378 4957
rect 20332 4885 20378 4923
rect 20332 4851 20338 4885
rect 20372 4851 20378 4885
rect 20332 4813 20378 4851
rect 20332 4779 20338 4813
rect 20372 4779 20378 4813
rect 20332 4741 20378 4779
rect 20332 4707 20338 4741
rect 20372 4707 20378 4741
rect 20332 4669 20378 4707
rect 20332 4635 20338 4669
rect 20372 4635 20378 4669
rect 20332 4597 20378 4635
rect 20332 4563 20338 4597
rect 20372 4563 20378 4597
rect 20332 4525 20378 4563
rect 20332 4491 20338 4525
rect 20372 4491 20378 4525
rect 20332 4453 20378 4491
rect 20332 4419 20338 4453
rect 20372 4419 20378 4453
rect 20332 4381 20378 4419
rect 20332 4347 20338 4381
rect 20372 4347 20378 4381
rect 20332 4309 20378 4347
rect 20332 4275 20338 4309
rect 20372 4275 20378 4309
rect 20332 4237 20378 4275
rect 20332 4203 20338 4237
rect 20372 4203 20378 4237
rect 20332 4165 20378 4203
rect 20332 4131 20338 4165
rect 20372 4131 20378 4165
rect 15704 4079 15750 4117
rect 20332 4116 20378 4131
rect 20428 5101 20474 5116
rect 20428 5067 20434 5101
rect 20468 5067 20474 5101
rect 20428 5029 20474 5067
rect 20428 4995 20434 5029
rect 20468 4995 20474 5029
rect 20428 4957 20474 4995
rect 20428 4923 20434 4957
rect 20468 4923 20474 4957
rect 20428 4885 20474 4923
rect 20428 4851 20434 4885
rect 20468 4851 20474 4885
rect 20428 4813 20474 4851
rect 20428 4779 20434 4813
rect 20468 4779 20474 4813
rect 20428 4741 20474 4779
rect 20428 4707 20434 4741
rect 20468 4707 20474 4741
rect 20428 4669 20474 4707
rect 20428 4635 20434 4669
rect 20468 4635 20474 4669
rect 20428 4597 20474 4635
rect 20428 4563 20434 4597
rect 20468 4563 20474 4597
rect 20428 4525 20474 4563
rect 20428 4491 20434 4525
rect 20468 4491 20474 4525
rect 20428 4453 20474 4491
rect 20428 4419 20434 4453
rect 20468 4419 20474 4453
rect 20428 4381 20474 4419
rect 20428 4347 20434 4381
rect 20468 4347 20474 4381
rect 20428 4309 20474 4347
rect 20428 4275 20434 4309
rect 20468 4275 20474 4309
rect 20428 4237 20474 4275
rect 20428 4203 20434 4237
rect 20468 4203 20474 4237
rect 20428 4165 20474 4203
rect 20428 4131 20434 4165
rect 20468 4131 20474 4165
rect 20428 4116 20474 4131
rect 20524 5101 20570 5116
rect 20524 5067 20530 5101
rect 20564 5067 20570 5101
rect 20524 5029 20570 5067
rect 20524 4995 20530 5029
rect 20564 4995 20570 5029
rect 20524 4957 20570 4995
rect 20524 4923 20530 4957
rect 20564 4923 20570 4957
rect 20524 4885 20570 4923
rect 20524 4851 20530 4885
rect 20564 4851 20570 4885
rect 20524 4813 20570 4851
rect 20524 4779 20530 4813
rect 20564 4779 20570 4813
rect 20524 4741 20570 4779
rect 20524 4707 20530 4741
rect 20564 4707 20570 4741
rect 20524 4669 20570 4707
rect 20524 4635 20530 4669
rect 20564 4635 20570 4669
rect 20524 4597 20570 4635
rect 20524 4563 20530 4597
rect 20564 4563 20570 4597
rect 20524 4525 20570 4563
rect 20524 4491 20530 4525
rect 20564 4491 20570 4525
rect 20524 4453 20570 4491
rect 20524 4419 20530 4453
rect 20564 4419 20570 4453
rect 20524 4381 20570 4419
rect 20524 4347 20530 4381
rect 20564 4347 20570 4381
rect 20524 4309 20570 4347
rect 20524 4275 20530 4309
rect 20564 4275 20570 4309
rect 20524 4237 20570 4275
rect 20524 4203 20530 4237
rect 20564 4203 20570 4237
rect 20524 4165 20570 4203
rect 20524 4131 20530 4165
rect 20564 4131 20570 4165
rect 20524 4116 20570 4131
rect 20620 5101 20666 5116
rect 20620 5067 20626 5101
rect 20660 5067 20666 5101
rect 20620 5029 20666 5067
rect 20620 4995 20626 5029
rect 20660 4995 20666 5029
rect 20620 4957 20666 4995
rect 20620 4923 20626 4957
rect 20660 4923 20666 4957
rect 20620 4885 20666 4923
rect 20620 4851 20626 4885
rect 20660 4851 20666 4885
rect 20620 4813 20666 4851
rect 20620 4779 20626 4813
rect 20660 4779 20666 4813
rect 20620 4741 20666 4779
rect 20620 4707 20626 4741
rect 20660 4707 20666 4741
rect 20620 4669 20666 4707
rect 20620 4635 20626 4669
rect 20660 4635 20666 4669
rect 20620 4597 20666 4635
rect 20620 4563 20626 4597
rect 20660 4563 20666 4597
rect 20620 4525 20666 4563
rect 20620 4491 20626 4525
rect 20660 4491 20666 4525
rect 20620 4453 20666 4491
rect 20620 4419 20626 4453
rect 20660 4419 20666 4453
rect 20620 4381 20666 4419
rect 20620 4347 20626 4381
rect 20660 4347 20666 4381
rect 20620 4309 20666 4347
rect 20620 4275 20626 4309
rect 20660 4275 20666 4309
rect 20620 4237 20666 4275
rect 20620 4203 20626 4237
rect 20660 4203 20666 4237
rect 20620 4165 20666 4203
rect 20620 4131 20626 4165
rect 20660 4131 20666 4165
rect 20620 4116 20666 4131
rect 20716 5101 20762 5116
rect 20716 5067 20722 5101
rect 20756 5067 20762 5101
rect 20716 5029 20762 5067
rect 20716 4995 20722 5029
rect 20756 4995 20762 5029
rect 20716 4957 20762 4995
rect 20716 4923 20722 4957
rect 20756 4923 20762 4957
rect 20716 4885 20762 4923
rect 20716 4851 20722 4885
rect 20756 4851 20762 4885
rect 20716 4813 20762 4851
rect 20716 4779 20722 4813
rect 20756 4779 20762 4813
rect 20716 4741 20762 4779
rect 20716 4707 20722 4741
rect 20756 4707 20762 4741
rect 20716 4669 20762 4707
rect 20716 4635 20722 4669
rect 20756 4635 20762 4669
rect 20716 4597 20762 4635
rect 20716 4563 20722 4597
rect 20756 4563 20762 4597
rect 20716 4525 20762 4563
rect 20716 4491 20722 4525
rect 20756 4491 20762 4525
rect 20716 4453 20762 4491
rect 20716 4419 20722 4453
rect 20756 4419 20762 4453
rect 20716 4381 20762 4419
rect 20716 4347 20722 4381
rect 20756 4347 20762 4381
rect 20716 4309 20762 4347
rect 20716 4275 20722 4309
rect 20756 4275 20762 4309
rect 20716 4237 20762 4275
rect 20716 4203 20722 4237
rect 20756 4203 20762 4237
rect 20716 4165 20762 4203
rect 20716 4131 20722 4165
rect 20756 4131 20762 4165
rect 20716 4116 20762 4131
rect 20812 5101 20858 5116
rect 20812 5067 20818 5101
rect 20852 5067 20858 5101
rect 20812 5029 20858 5067
rect 20812 4995 20818 5029
rect 20852 4995 20858 5029
rect 20812 4957 20858 4995
rect 20812 4923 20818 4957
rect 20852 4923 20858 4957
rect 20812 4885 20858 4923
rect 20812 4851 20818 4885
rect 20852 4851 20858 4885
rect 20812 4813 20858 4851
rect 20812 4779 20818 4813
rect 20852 4779 20858 4813
rect 20812 4741 20858 4779
rect 20812 4707 20818 4741
rect 20852 4707 20858 4741
rect 20812 4669 20858 4707
rect 20812 4635 20818 4669
rect 20852 4635 20858 4669
rect 20812 4597 20858 4635
rect 20812 4563 20818 4597
rect 20852 4563 20858 4597
rect 20812 4525 20858 4563
rect 20812 4491 20818 4525
rect 20852 4491 20858 4525
rect 20812 4453 20858 4491
rect 20812 4419 20818 4453
rect 20852 4419 20858 4453
rect 20812 4381 20858 4419
rect 20812 4347 20818 4381
rect 20852 4347 20858 4381
rect 20812 4309 20858 4347
rect 20812 4275 20818 4309
rect 20852 4275 20858 4309
rect 20812 4237 20858 4275
rect 20812 4203 20818 4237
rect 20852 4203 20858 4237
rect 20812 4165 20858 4203
rect 20812 4131 20818 4165
rect 20852 4131 20858 4165
rect 20812 4116 20858 4131
rect 20908 5101 20954 5116
rect 20908 5067 20914 5101
rect 20948 5067 20954 5101
rect 20908 5029 20954 5067
rect 20908 4995 20914 5029
rect 20948 4995 20954 5029
rect 20908 4957 20954 4995
rect 20908 4923 20914 4957
rect 20948 4923 20954 4957
rect 20908 4885 20954 4923
rect 20908 4851 20914 4885
rect 20948 4851 20954 4885
rect 20908 4813 20954 4851
rect 20908 4779 20914 4813
rect 20948 4779 20954 4813
rect 20908 4741 20954 4779
rect 20908 4707 20914 4741
rect 20948 4707 20954 4741
rect 20908 4669 20954 4707
rect 20908 4635 20914 4669
rect 20948 4635 20954 4669
rect 20908 4597 20954 4635
rect 20908 4563 20914 4597
rect 20948 4563 20954 4597
rect 20908 4525 20954 4563
rect 20908 4491 20914 4525
rect 20948 4491 20954 4525
rect 20908 4453 20954 4491
rect 20908 4419 20914 4453
rect 20948 4419 20954 4453
rect 20908 4381 20954 4419
rect 20908 4347 20914 4381
rect 20948 4347 20954 4381
rect 20908 4309 20954 4347
rect 20908 4275 20914 4309
rect 20948 4275 20954 4309
rect 20908 4237 20954 4275
rect 20908 4203 20914 4237
rect 20948 4203 20954 4237
rect 20908 4165 20954 4203
rect 20908 4131 20914 4165
rect 20948 4131 20954 4165
rect 20908 4116 20954 4131
rect 21004 5101 21050 5116
rect 21004 5067 21010 5101
rect 21044 5067 21050 5101
rect 21004 5029 21050 5067
rect 21004 4995 21010 5029
rect 21044 4995 21050 5029
rect 21004 4957 21050 4995
rect 21004 4923 21010 4957
rect 21044 4923 21050 4957
rect 21004 4885 21050 4923
rect 21004 4851 21010 4885
rect 21044 4851 21050 4885
rect 21004 4813 21050 4851
rect 21004 4779 21010 4813
rect 21044 4779 21050 4813
rect 21004 4741 21050 4779
rect 21004 4707 21010 4741
rect 21044 4707 21050 4741
rect 21004 4669 21050 4707
rect 21004 4635 21010 4669
rect 21044 4635 21050 4669
rect 21004 4597 21050 4635
rect 21004 4563 21010 4597
rect 21044 4563 21050 4597
rect 21004 4525 21050 4563
rect 21004 4491 21010 4525
rect 21044 4491 21050 4525
rect 21004 4453 21050 4491
rect 21004 4419 21010 4453
rect 21044 4419 21050 4453
rect 21004 4381 21050 4419
rect 21004 4347 21010 4381
rect 21044 4347 21050 4381
rect 21004 4309 21050 4347
rect 21004 4275 21010 4309
rect 21044 4275 21050 4309
rect 21004 4237 21050 4275
rect 21004 4203 21010 4237
rect 21044 4203 21050 4237
rect 21004 4165 21050 4203
rect 21004 4131 21010 4165
rect 21044 4131 21050 4165
rect 21004 4116 21050 4131
rect 21100 5101 21146 5116
rect 21100 5067 21106 5101
rect 21140 5067 21146 5101
rect 21100 5029 21146 5067
rect 21100 4995 21106 5029
rect 21140 4995 21146 5029
rect 21100 4957 21146 4995
rect 21100 4923 21106 4957
rect 21140 4923 21146 4957
rect 21100 4885 21146 4923
rect 21100 4851 21106 4885
rect 21140 4851 21146 4885
rect 21100 4813 21146 4851
rect 21100 4779 21106 4813
rect 21140 4779 21146 4813
rect 21100 4741 21146 4779
rect 21100 4707 21106 4741
rect 21140 4707 21146 4741
rect 21100 4669 21146 4707
rect 21100 4635 21106 4669
rect 21140 4635 21146 4669
rect 21100 4597 21146 4635
rect 21100 4563 21106 4597
rect 21140 4563 21146 4597
rect 21100 4525 21146 4563
rect 21100 4491 21106 4525
rect 21140 4491 21146 4525
rect 21100 4453 21146 4491
rect 21100 4419 21106 4453
rect 21140 4419 21146 4453
rect 21100 4381 21146 4419
rect 21100 4347 21106 4381
rect 21140 4347 21146 4381
rect 21100 4309 21146 4347
rect 21100 4275 21106 4309
rect 21140 4275 21146 4309
rect 21100 4237 21146 4275
rect 21100 4203 21106 4237
rect 21140 4203 21146 4237
rect 21100 4165 21146 4203
rect 21100 4131 21106 4165
rect 21140 4131 21146 4165
rect 21100 4116 21146 4131
rect 21196 5101 21242 5116
rect 21196 5067 21202 5101
rect 21236 5067 21242 5101
rect 21196 5029 21242 5067
rect 21196 4995 21202 5029
rect 21236 4995 21242 5029
rect 21196 4957 21242 4995
rect 21196 4923 21202 4957
rect 21236 4923 21242 4957
rect 21196 4885 21242 4923
rect 21196 4851 21202 4885
rect 21236 4851 21242 4885
rect 21196 4813 21242 4851
rect 21196 4779 21202 4813
rect 21236 4779 21242 4813
rect 21196 4741 21242 4779
rect 21196 4707 21202 4741
rect 21236 4707 21242 4741
rect 21196 4669 21242 4707
rect 21196 4635 21202 4669
rect 21236 4635 21242 4669
rect 21196 4597 21242 4635
rect 21196 4563 21202 4597
rect 21236 4563 21242 4597
rect 21196 4525 21242 4563
rect 21196 4491 21202 4525
rect 21236 4491 21242 4525
rect 21196 4453 21242 4491
rect 21196 4419 21202 4453
rect 21236 4419 21242 4453
rect 21196 4381 21242 4419
rect 21196 4347 21202 4381
rect 21236 4347 21242 4381
rect 21196 4309 21242 4347
rect 21196 4275 21202 4309
rect 21236 4275 21242 4309
rect 21196 4237 21242 4275
rect 21196 4203 21202 4237
rect 21236 4203 21242 4237
rect 21196 4165 21242 4203
rect 21196 4131 21202 4165
rect 21236 4131 21242 4165
rect 21196 4116 21242 4131
rect 21292 5101 21338 5116
rect 21292 5067 21298 5101
rect 21332 5067 21338 5101
rect 21292 5029 21338 5067
rect 21292 4995 21298 5029
rect 21332 4995 21338 5029
rect 21292 4957 21338 4995
rect 21292 4923 21298 4957
rect 21332 4923 21338 4957
rect 21292 4885 21338 4923
rect 21292 4851 21298 4885
rect 21332 4851 21338 4885
rect 21292 4813 21338 4851
rect 21292 4779 21298 4813
rect 21332 4779 21338 4813
rect 21292 4741 21338 4779
rect 21292 4707 21298 4741
rect 21332 4707 21338 4741
rect 21292 4669 21338 4707
rect 21292 4635 21298 4669
rect 21332 4635 21338 4669
rect 21292 4597 21338 4635
rect 21292 4563 21298 4597
rect 21332 4563 21338 4597
rect 21292 4525 21338 4563
rect 21292 4491 21298 4525
rect 21332 4491 21338 4525
rect 21292 4453 21338 4491
rect 21292 4419 21298 4453
rect 21332 4419 21338 4453
rect 21292 4381 21338 4419
rect 21292 4347 21298 4381
rect 21332 4347 21338 4381
rect 21292 4309 21338 4347
rect 21292 4275 21298 4309
rect 21332 4275 21338 4309
rect 21292 4237 21338 4275
rect 21292 4203 21298 4237
rect 21332 4203 21338 4237
rect 21292 4165 21338 4203
rect 21292 4131 21298 4165
rect 21332 4131 21338 4165
rect 21292 4116 21338 4131
rect 21388 5101 21434 5116
rect 21388 5067 21394 5101
rect 21428 5067 21434 5101
rect 21388 5029 21434 5067
rect 21388 4995 21394 5029
rect 21428 4995 21434 5029
rect 21388 4957 21434 4995
rect 21388 4923 21394 4957
rect 21428 4923 21434 4957
rect 21388 4885 21434 4923
rect 21388 4851 21394 4885
rect 21428 4851 21434 4885
rect 21388 4813 21434 4851
rect 21388 4779 21394 4813
rect 21428 4779 21434 4813
rect 21388 4741 21434 4779
rect 21388 4707 21394 4741
rect 21428 4707 21434 4741
rect 21388 4669 21434 4707
rect 21388 4635 21394 4669
rect 21428 4635 21434 4669
rect 21388 4597 21434 4635
rect 21388 4563 21394 4597
rect 21428 4563 21434 4597
rect 21388 4525 21434 4563
rect 21388 4491 21394 4525
rect 21428 4491 21434 4525
rect 21388 4453 21434 4491
rect 21388 4419 21394 4453
rect 21428 4419 21434 4453
rect 21388 4381 21434 4419
rect 21388 4347 21394 4381
rect 21428 4347 21434 4381
rect 21388 4309 21434 4347
rect 21388 4275 21394 4309
rect 21428 4275 21434 4309
rect 21388 4237 21434 4275
rect 21388 4203 21394 4237
rect 21428 4203 21434 4237
rect 21388 4165 21434 4203
rect 21388 4131 21394 4165
rect 21428 4131 21434 4165
rect 21388 4116 21434 4131
rect 21484 5101 21530 5116
rect 21484 5067 21490 5101
rect 21524 5067 21530 5101
rect 21484 5029 21530 5067
rect 21484 4995 21490 5029
rect 21524 4995 21530 5029
rect 21484 4957 21530 4995
rect 21484 4923 21490 4957
rect 21524 4923 21530 4957
rect 21484 4885 21530 4923
rect 21484 4851 21490 4885
rect 21524 4851 21530 4885
rect 21484 4813 21530 4851
rect 21484 4779 21490 4813
rect 21524 4779 21530 4813
rect 21484 4741 21530 4779
rect 21484 4707 21490 4741
rect 21524 4707 21530 4741
rect 21484 4669 21530 4707
rect 21484 4635 21490 4669
rect 21524 4635 21530 4669
rect 21484 4597 21530 4635
rect 21484 4563 21490 4597
rect 21524 4563 21530 4597
rect 21484 4525 21530 4563
rect 21484 4491 21490 4525
rect 21524 4491 21530 4525
rect 21484 4453 21530 4491
rect 21484 4419 21490 4453
rect 21524 4419 21530 4453
rect 21484 4381 21530 4419
rect 21484 4347 21490 4381
rect 21524 4347 21530 4381
rect 21484 4309 21530 4347
rect 21484 4275 21490 4309
rect 21524 4275 21530 4309
rect 21484 4237 21530 4275
rect 21484 4203 21490 4237
rect 21524 4203 21530 4237
rect 21484 4165 21530 4203
rect 21484 4131 21490 4165
rect 21524 4131 21530 4165
rect 21484 4116 21530 4131
rect 21580 5101 21626 5116
rect 21580 5067 21586 5101
rect 21620 5067 21626 5101
rect 21580 5029 21626 5067
rect 21580 4995 21586 5029
rect 21620 4995 21626 5029
rect 21580 4957 21626 4995
rect 21580 4923 21586 4957
rect 21620 4923 21626 4957
rect 21580 4885 21626 4923
rect 21580 4851 21586 4885
rect 21620 4851 21626 4885
rect 21580 4813 21626 4851
rect 21580 4779 21586 4813
rect 21620 4779 21626 4813
rect 21580 4741 21626 4779
rect 21580 4707 21586 4741
rect 21620 4707 21626 4741
rect 21580 4669 21626 4707
rect 21580 4635 21586 4669
rect 21620 4635 21626 4669
rect 21580 4597 21626 4635
rect 21580 4563 21586 4597
rect 21620 4563 21626 4597
rect 21580 4525 21626 4563
rect 21580 4491 21586 4525
rect 21620 4491 21626 4525
rect 21580 4453 21626 4491
rect 21580 4419 21586 4453
rect 21620 4419 21626 4453
rect 21580 4381 21626 4419
rect 21580 4347 21586 4381
rect 21620 4347 21626 4381
rect 21580 4309 21626 4347
rect 21580 4275 21586 4309
rect 21620 4275 21626 4309
rect 21580 4237 21626 4275
rect 21580 4203 21586 4237
rect 21620 4203 21626 4237
rect 21580 4165 21626 4203
rect 21580 4131 21586 4165
rect 21620 4131 21626 4165
rect 21580 4116 21626 4131
rect 21676 5101 21722 5116
rect 21676 5067 21682 5101
rect 21716 5067 21722 5101
rect 21676 5029 21722 5067
rect 21676 4995 21682 5029
rect 21716 4995 21722 5029
rect 21676 4957 21722 4995
rect 21676 4923 21682 4957
rect 21716 4923 21722 4957
rect 21676 4885 21722 4923
rect 21676 4851 21682 4885
rect 21716 4851 21722 4885
rect 21676 4813 21722 4851
rect 21676 4779 21682 4813
rect 21716 4779 21722 4813
rect 21676 4741 21722 4779
rect 21676 4707 21682 4741
rect 21716 4707 21722 4741
rect 21676 4669 21722 4707
rect 21676 4635 21682 4669
rect 21716 4635 21722 4669
rect 21676 4597 21722 4635
rect 21676 4563 21682 4597
rect 21716 4563 21722 4597
rect 21676 4525 21722 4563
rect 21676 4491 21682 4525
rect 21716 4491 21722 4525
rect 21676 4453 21722 4491
rect 21676 4419 21682 4453
rect 21716 4419 21722 4453
rect 21676 4381 21722 4419
rect 21676 4347 21682 4381
rect 21716 4347 21722 4381
rect 21676 4309 21722 4347
rect 21676 4275 21682 4309
rect 21716 4275 21722 4309
rect 21676 4237 21722 4275
rect 21676 4203 21682 4237
rect 21716 4203 21722 4237
rect 21676 4165 21722 4203
rect 21676 4131 21682 4165
rect 21716 4131 21722 4165
rect 21676 4116 21722 4131
rect 21772 5101 21818 5116
rect 21772 5067 21778 5101
rect 21812 5067 21818 5101
rect 21772 5029 21818 5067
rect 21772 4995 21778 5029
rect 21812 4995 21818 5029
rect 21772 4957 21818 4995
rect 21772 4923 21778 4957
rect 21812 4923 21818 4957
rect 21772 4885 21818 4923
rect 21772 4851 21778 4885
rect 21812 4851 21818 4885
rect 21772 4813 21818 4851
rect 21772 4779 21778 4813
rect 21812 4779 21818 4813
rect 21772 4741 21818 4779
rect 21772 4707 21778 4741
rect 21812 4707 21818 4741
rect 21772 4669 21818 4707
rect 21772 4635 21778 4669
rect 21812 4635 21818 4669
rect 21772 4597 21818 4635
rect 21772 4563 21778 4597
rect 21812 4563 21818 4597
rect 21772 4525 21818 4563
rect 21772 4491 21778 4525
rect 21812 4491 21818 4525
rect 21772 4453 21818 4491
rect 21772 4419 21778 4453
rect 21812 4419 21818 4453
rect 21772 4381 21818 4419
rect 21772 4347 21778 4381
rect 21812 4347 21818 4381
rect 21772 4309 21818 4347
rect 21772 4275 21778 4309
rect 21812 4275 21818 4309
rect 21772 4237 21818 4275
rect 21772 4203 21778 4237
rect 21812 4203 21818 4237
rect 21772 4165 21818 4203
rect 21772 4131 21778 4165
rect 21812 4131 21818 4165
rect 21772 4116 21818 4131
rect 21868 5101 21914 5116
rect 21868 5067 21874 5101
rect 21908 5067 21914 5101
rect 21868 5029 21914 5067
rect 21868 4995 21874 5029
rect 21908 4995 21914 5029
rect 21868 4957 21914 4995
rect 21868 4923 21874 4957
rect 21908 4923 21914 4957
rect 21868 4885 21914 4923
rect 21868 4851 21874 4885
rect 21908 4851 21914 4885
rect 21868 4813 21914 4851
rect 21868 4779 21874 4813
rect 21908 4779 21914 4813
rect 21868 4741 21914 4779
rect 21868 4707 21874 4741
rect 21908 4707 21914 4741
rect 21868 4669 21914 4707
rect 21868 4635 21874 4669
rect 21908 4635 21914 4669
rect 21868 4597 21914 4635
rect 21868 4563 21874 4597
rect 21908 4563 21914 4597
rect 21868 4525 21914 4563
rect 21868 4491 21874 4525
rect 21908 4491 21914 4525
rect 21868 4453 21914 4491
rect 21868 4419 21874 4453
rect 21908 4419 21914 4453
rect 21868 4381 21914 4419
rect 21868 4347 21874 4381
rect 21908 4347 21914 4381
rect 21868 4309 21914 4347
rect 21868 4275 21874 4309
rect 21908 4275 21914 4309
rect 21868 4237 21914 4275
rect 21868 4203 21874 4237
rect 21908 4203 21914 4237
rect 21868 4165 21914 4203
rect 21868 4131 21874 4165
rect 21908 4131 21914 4165
rect 21868 4116 21914 4131
rect 21964 5101 22010 5116
rect 21964 5067 21970 5101
rect 22004 5067 22010 5101
rect 21964 5029 22010 5067
rect 21964 4995 21970 5029
rect 22004 4995 22010 5029
rect 21964 4957 22010 4995
rect 21964 4923 21970 4957
rect 22004 4923 22010 4957
rect 21964 4885 22010 4923
rect 21964 4851 21970 4885
rect 22004 4851 22010 4885
rect 21964 4813 22010 4851
rect 21964 4779 21970 4813
rect 22004 4779 22010 4813
rect 21964 4741 22010 4779
rect 21964 4707 21970 4741
rect 22004 4707 22010 4741
rect 21964 4669 22010 4707
rect 21964 4635 21970 4669
rect 22004 4635 22010 4669
rect 21964 4597 22010 4635
rect 21964 4563 21970 4597
rect 22004 4563 22010 4597
rect 21964 4525 22010 4563
rect 21964 4491 21970 4525
rect 22004 4491 22010 4525
rect 21964 4453 22010 4491
rect 21964 4419 21970 4453
rect 22004 4419 22010 4453
rect 21964 4381 22010 4419
rect 21964 4347 21970 4381
rect 22004 4347 22010 4381
rect 21964 4309 22010 4347
rect 21964 4275 21970 4309
rect 22004 4275 22010 4309
rect 21964 4237 22010 4275
rect 21964 4203 21970 4237
rect 22004 4203 22010 4237
rect 21964 4165 22010 4203
rect 21964 4131 21970 4165
rect 22004 4131 22010 4165
rect 21964 4116 22010 4131
rect 22060 5101 22106 5116
rect 22060 5067 22066 5101
rect 22100 5067 22106 5101
rect 22060 5029 22106 5067
rect 22060 4995 22066 5029
rect 22100 4995 22106 5029
rect 22060 4957 22106 4995
rect 22060 4923 22066 4957
rect 22100 4923 22106 4957
rect 22060 4885 22106 4923
rect 22060 4851 22066 4885
rect 22100 4851 22106 4885
rect 22060 4813 22106 4851
rect 22060 4779 22066 4813
rect 22100 4779 22106 4813
rect 22060 4741 22106 4779
rect 22060 4707 22066 4741
rect 22100 4707 22106 4741
rect 22060 4669 22106 4707
rect 22060 4635 22066 4669
rect 22100 4635 22106 4669
rect 22060 4597 22106 4635
rect 22060 4563 22066 4597
rect 22100 4563 22106 4597
rect 22060 4525 22106 4563
rect 22060 4491 22066 4525
rect 22100 4491 22106 4525
rect 22060 4453 22106 4491
rect 22060 4419 22066 4453
rect 22100 4419 22106 4453
rect 22060 4381 22106 4419
rect 22060 4347 22066 4381
rect 22100 4347 22106 4381
rect 22060 4309 22106 4347
rect 22060 4275 22066 4309
rect 22100 4275 22106 4309
rect 22060 4237 22106 4275
rect 22060 4203 22066 4237
rect 22100 4203 22106 4237
rect 22060 4165 22106 4203
rect 22060 4131 22066 4165
rect 22100 4131 22106 4165
rect 22060 4116 22106 4131
rect 22156 5101 22202 5116
rect 22156 5067 22162 5101
rect 22196 5067 22202 5101
rect 22156 5029 22202 5067
rect 22156 4995 22162 5029
rect 22196 4995 22202 5029
rect 22156 4957 22202 4995
rect 22156 4923 22162 4957
rect 22196 4923 22202 4957
rect 22156 4885 22202 4923
rect 22156 4851 22162 4885
rect 22196 4851 22202 4885
rect 22156 4813 22202 4851
rect 22156 4779 22162 4813
rect 22196 4779 22202 4813
rect 22156 4741 22202 4779
rect 22156 4707 22162 4741
rect 22196 4707 22202 4741
rect 22156 4669 22202 4707
rect 22156 4635 22162 4669
rect 22196 4635 22202 4669
rect 22156 4597 22202 4635
rect 22156 4563 22162 4597
rect 22196 4563 22202 4597
rect 22156 4525 22202 4563
rect 22156 4491 22162 4525
rect 22196 4491 22202 4525
rect 22156 4453 22202 4491
rect 22156 4419 22162 4453
rect 22196 4419 22202 4453
rect 22156 4381 22202 4419
rect 22156 4347 22162 4381
rect 22196 4347 22202 4381
rect 22156 4309 22202 4347
rect 22156 4275 22162 4309
rect 22196 4275 22202 4309
rect 22156 4237 22202 4275
rect 22156 4203 22162 4237
rect 22196 4203 22202 4237
rect 22156 4165 22202 4203
rect 22156 4131 22162 4165
rect 22196 4131 22202 4165
rect 22156 4116 22202 4131
rect 22252 5101 22298 5116
rect 22252 5067 22258 5101
rect 22292 5067 22298 5101
rect 22252 5029 22298 5067
rect 22252 4995 22258 5029
rect 22292 4995 22298 5029
rect 22252 4957 22298 4995
rect 22252 4923 22258 4957
rect 22292 4923 22298 4957
rect 22252 4885 22298 4923
rect 22252 4851 22258 4885
rect 22292 4851 22298 4885
rect 22252 4813 22298 4851
rect 22252 4779 22258 4813
rect 22292 4779 22298 4813
rect 22252 4741 22298 4779
rect 22252 4707 22258 4741
rect 22292 4707 22298 4741
rect 22252 4669 22298 4707
rect 22252 4635 22258 4669
rect 22292 4635 22298 4669
rect 22252 4597 22298 4635
rect 22252 4563 22258 4597
rect 22292 4563 22298 4597
rect 22252 4525 22298 4563
rect 22252 4491 22258 4525
rect 22292 4491 22298 4525
rect 22252 4453 22298 4491
rect 22252 4419 22258 4453
rect 22292 4419 22298 4453
rect 22252 4381 22298 4419
rect 22252 4347 22258 4381
rect 22292 4347 22298 4381
rect 22252 4309 22298 4347
rect 22252 4275 22258 4309
rect 22292 4275 22298 4309
rect 22252 4237 22298 4275
rect 22252 4203 22258 4237
rect 22292 4203 22298 4237
rect 22252 4165 22298 4203
rect 22252 4131 22258 4165
rect 22292 4131 22298 4165
rect 22252 4116 22298 4131
rect 23264 5113 23310 5128
rect 23264 5079 23270 5113
rect 23304 5079 23310 5113
rect 23264 5041 23310 5079
rect 23264 5007 23270 5041
rect 23304 5007 23310 5041
rect 23264 4969 23310 5007
rect 23264 4935 23270 4969
rect 23304 4935 23310 4969
rect 23264 4897 23310 4935
rect 23264 4863 23270 4897
rect 23304 4863 23310 4897
rect 23264 4825 23310 4863
rect 23264 4791 23270 4825
rect 23304 4791 23310 4825
rect 23264 4753 23310 4791
rect 23264 4719 23270 4753
rect 23304 4719 23310 4753
rect 23264 4681 23310 4719
rect 23264 4647 23270 4681
rect 23304 4647 23310 4681
rect 23264 4609 23310 4647
rect 23264 4575 23270 4609
rect 23304 4575 23310 4609
rect 23264 4537 23310 4575
rect 23264 4503 23270 4537
rect 23304 4503 23310 4537
rect 23264 4465 23310 4503
rect 23264 4431 23270 4465
rect 23304 4431 23310 4465
rect 23264 4393 23310 4431
rect 23264 4359 23270 4393
rect 23304 4359 23310 4393
rect 23264 4321 23310 4359
rect 23264 4287 23270 4321
rect 23304 4287 23310 4321
rect 23264 4249 23310 4287
rect 23264 4215 23270 4249
rect 23304 4215 23310 4249
rect 23264 4177 23310 4215
rect 23264 4143 23270 4177
rect 23304 4143 23310 4177
rect 23264 4128 23310 4143
rect 23360 5113 23406 5128
rect 23360 5079 23366 5113
rect 23400 5079 23406 5113
rect 23360 5041 23406 5079
rect 23360 5007 23366 5041
rect 23400 5007 23406 5041
rect 23360 4969 23406 5007
rect 23360 4935 23366 4969
rect 23400 4935 23406 4969
rect 23360 4897 23406 4935
rect 23360 4863 23366 4897
rect 23400 4863 23406 4897
rect 23360 4825 23406 4863
rect 23360 4791 23366 4825
rect 23400 4791 23406 4825
rect 23360 4753 23406 4791
rect 23360 4719 23366 4753
rect 23400 4719 23406 4753
rect 23360 4681 23406 4719
rect 23360 4647 23366 4681
rect 23400 4647 23406 4681
rect 23360 4609 23406 4647
rect 23360 4575 23366 4609
rect 23400 4575 23406 4609
rect 23360 4537 23406 4575
rect 23360 4503 23366 4537
rect 23400 4503 23406 4537
rect 23360 4465 23406 4503
rect 23360 4431 23366 4465
rect 23400 4431 23406 4465
rect 23360 4393 23406 4431
rect 23360 4359 23366 4393
rect 23400 4359 23406 4393
rect 23360 4321 23406 4359
rect 23360 4287 23366 4321
rect 23400 4287 23406 4321
rect 23360 4249 23406 4287
rect 23360 4215 23366 4249
rect 23400 4215 23406 4249
rect 23360 4177 23406 4215
rect 23360 4143 23366 4177
rect 23400 4143 23406 4177
rect 23360 4128 23406 4143
rect 23456 5113 23502 5128
rect 23456 5079 23462 5113
rect 23496 5079 23502 5113
rect 23456 5041 23502 5079
rect 23456 5007 23462 5041
rect 23496 5007 23502 5041
rect 23456 4969 23502 5007
rect 23456 4935 23462 4969
rect 23496 4935 23502 4969
rect 23456 4897 23502 4935
rect 23456 4863 23462 4897
rect 23496 4863 23502 4897
rect 23456 4825 23502 4863
rect 23456 4791 23462 4825
rect 23496 4791 23502 4825
rect 23456 4753 23502 4791
rect 23456 4719 23462 4753
rect 23496 4719 23502 4753
rect 23456 4681 23502 4719
rect 23456 4647 23462 4681
rect 23496 4647 23502 4681
rect 23456 4609 23502 4647
rect 23456 4575 23462 4609
rect 23496 4575 23502 4609
rect 23456 4537 23502 4575
rect 23456 4503 23462 4537
rect 23496 4503 23502 4537
rect 23456 4465 23502 4503
rect 23456 4431 23462 4465
rect 23496 4431 23502 4465
rect 23456 4393 23502 4431
rect 23456 4359 23462 4393
rect 23496 4359 23502 4393
rect 23456 4321 23502 4359
rect 23456 4287 23462 4321
rect 23496 4287 23502 4321
rect 23456 4249 23502 4287
rect 23456 4215 23462 4249
rect 23496 4215 23502 4249
rect 23456 4177 23502 4215
rect 23456 4143 23462 4177
rect 23496 4143 23502 4177
rect 23456 4128 23502 4143
rect 23552 5113 23598 5128
rect 23552 5079 23558 5113
rect 23592 5079 23598 5113
rect 23552 5041 23598 5079
rect 23552 5007 23558 5041
rect 23592 5007 23598 5041
rect 23552 4969 23598 5007
rect 23552 4935 23558 4969
rect 23592 4935 23598 4969
rect 23552 4897 23598 4935
rect 23552 4863 23558 4897
rect 23592 4863 23598 4897
rect 23552 4825 23598 4863
rect 23552 4791 23558 4825
rect 23592 4791 23598 4825
rect 23552 4753 23598 4791
rect 23552 4719 23558 4753
rect 23592 4719 23598 4753
rect 23552 4681 23598 4719
rect 23552 4647 23558 4681
rect 23592 4647 23598 4681
rect 23552 4609 23598 4647
rect 23552 4575 23558 4609
rect 23592 4575 23598 4609
rect 23552 4537 23598 4575
rect 23552 4503 23558 4537
rect 23592 4503 23598 4537
rect 23552 4465 23598 4503
rect 23552 4431 23558 4465
rect 23592 4431 23598 4465
rect 23552 4393 23598 4431
rect 23552 4359 23558 4393
rect 23592 4359 23598 4393
rect 23552 4321 23598 4359
rect 23552 4287 23558 4321
rect 23592 4287 23598 4321
rect 23552 4249 23598 4287
rect 23552 4215 23558 4249
rect 23592 4215 23598 4249
rect 23552 4177 23598 4215
rect 23552 4143 23558 4177
rect 23592 4143 23598 4177
rect 23552 4128 23598 4143
rect 23648 5113 23694 5128
rect 23648 5079 23654 5113
rect 23688 5079 23694 5113
rect 23648 5041 23694 5079
rect 23648 5007 23654 5041
rect 23688 5007 23694 5041
rect 23648 4969 23694 5007
rect 23648 4935 23654 4969
rect 23688 4935 23694 4969
rect 23648 4897 23694 4935
rect 23648 4863 23654 4897
rect 23688 4863 23694 4897
rect 23648 4825 23694 4863
rect 23648 4791 23654 4825
rect 23688 4791 23694 4825
rect 23648 4753 23694 4791
rect 23648 4719 23654 4753
rect 23688 4719 23694 4753
rect 23648 4681 23694 4719
rect 23648 4647 23654 4681
rect 23688 4647 23694 4681
rect 23648 4609 23694 4647
rect 23648 4575 23654 4609
rect 23688 4575 23694 4609
rect 23648 4537 23694 4575
rect 23648 4503 23654 4537
rect 23688 4503 23694 4537
rect 23648 4465 23694 4503
rect 23648 4431 23654 4465
rect 23688 4431 23694 4465
rect 23648 4393 23694 4431
rect 23648 4359 23654 4393
rect 23688 4359 23694 4393
rect 23648 4321 23694 4359
rect 23648 4287 23654 4321
rect 23688 4287 23694 4321
rect 23648 4249 23694 4287
rect 23648 4215 23654 4249
rect 23688 4215 23694 4249
rect 23648 4177 23694 4215
rect 23648 4143 23654 4177
rect 23688 4143 23694 4177
rect 23648 4128 23694 4143
rect 23744 5113 23790 5128
rect 23744 5079 23750 5113
rect 23784 5079 23790 5113
rect 23744 5041 23790 5079
rect 23744 5007 23750 5041
rect 23784 5007 23790 5041
rect 23744 4969 23790 5007
rect 23744 4935 23750 4969
rect 23784 4935 23790 4969
rect 23744 4897 23790 4935
rect 23744 4863 23750 4897
rect 23784 4863 23790 4897
rect 23744 4825 23790 4863
rect 23744 4791 23750 4825
rect 23784 4791 23790 4825
rect 23744 4753 23790 4791
rect 23744 4719 23750 4753
rect 23784 4719 23790 4753
rect 23744 4681 23790 4719
rect 23744 4647 23750 4681
rect 23784 4647 23790 4681
rect 23744 4609 23790 4647
rect 23744 4575 23750 4609
rect 23784 4575 23790 4609
rect 23744 4537 23790 4575
rect 23744 4503 23750 4537
rect 23784 4503 23790 4537
rect 23744 4465 23790 4503
rect 23744 4431 23750 4465
rect 23784 4431 23790 4465
rect 23744 4393 23790 4431
rect 23744 4359 23750 4393
rect 23784 4359 23790 4393
rect 23744 4321 23790 4359
rect 23744 4287 23750 4321
rect 23784 4287 23790 4321
rect 23744 4249 23790 4287
rect 23744 4215 23750 4249
rect 23784 4215 23790 4249
rect 23744 4177 23790 4215
rect 23744 4143 23750 4177
rect 23784 4143 23790 4177
rect 23744 4128 23790 4143
rect 23952 5111 23998 5126
rect 23952 5077 23958 5111
rect 23992 5077 23998 5111
rect 23952 5039 23998 5077
rect 23952 5005 23958 5039
rect 23992 5005 23998 5039
rect 23952 4967 23998 5005
rect 23952 4933 23958 4967
rect 23992 4933 23998 4967
rect 23952 4895 23998 4933
rect 23952 4861 23958 4895
rect 23992 4861 23998 4895
rect 23952 4823 23998 4861
rect 23952 4789 23958 4823
rect 23992 4789 23998 4823
rect 23952 4751 23998 4789
rect 23952 4717 23958 4751
rect 23992 4717 23998 4751
rect 23952 4679 23998 4717
rect 23952 4645 23958 4679
rect 23992 4645 23998 4679
rect 23952 4607 23998 4645
rect 23952 4573 23958 4607
rect 23992 4573 23998 4607
rect 23952 4535 23998 4573
rect 23952 4501 23958 4535
rect 23992 4501 23998 4535
rect 23952 4463 23998 4501
rect 23952 4429 23958 4463
rect 23992 4429 23998 4463
rect 23952 4391 23998 4429
rect 23952 4357 23958 4391
rect 23992 4357 23998 4391
rect 23952 4319 23998 4357
rect 23952 4285 23958 4319
rect 23992 4285 23998 4319
rect 23952 4247 23998 4285
rect 23952 4213 23958 4247
rect 23992 4213 23998 4247
rect 23952 4175 23998 4213
rect 23952 4141 23958 4175
rect 23992 4141 23998 4175
rect 23952 4126 23998 4141
rect 24048 5111 24094 5126
rect 24048 5077 24054 5111
rect 24088 5077 24094 5111
rect 24048 5039 24094 5077
rect 24048 5005 24054 5039
rect 24088 5005 24094 5039
rect 24048 4967 24094 5005
rect 24048 4933 24054 4967
rect 24088 4933 24094 4967
rect 24048 4895 24094 4933
rect 24048 4861 24054 4895
rect 24088 4861 24094 4895
rect 24048 4823 24094 4861
rect 24048 4789 24054 4823
rect 24088 4789 24094 4823
rect 24048 4751 24094 4789
rect 24048 4717 24054 4751
rect 24088 4717 24094 4751
rect 24048 4679 24094 4717
rect 24048 4645 24054 4679
rect 24088 4645 24094 4679
rect 24048 4607 24094 4645
rect 24048 4573 24054 4607
rect 24088 4573 24094 4607
rect 24048 4535 24094 4573
rect 24048 4501 24054 4535
rect 24088 4501 24094 4535
rect 24048 4463 24094 4501
rect 24048 4429 24054 4463
rect 24088 4429 24094 4463
rect 24048 4391 24094 4429
rect 24048 4357 24054 4391
rect 24088 4357 24094 4391
rect 24048 4319 24094 4357
rect 24048 4285 24054 4319
rect 24088 4285 24094 4319
rect 24048 4247 24094 4285
rect 24048 4213 24054 4247
rect 24088 4213 24094 4247
rect 24048 4175 24094 4213
rect 24048 4141 24054 4175
rect 24088 4141 24094 4175
rect 24048 4126 24094 4141
rect 24144 5111 24190 5126
rect 24144 5077 24150 5111
rect 24184 5077 24190 5111
rect 24144 5039 24190 5077
rect 24144 5005 24150 5039
rect 24184 5005 24190 5039
rect 24144 4967 24190 5005
rect 24144 4933 24150 4967
rect 24184 4933 24190 4967
rect 24144 4895 24190 4933
rect 24144 4861 24150 4895
rect 24184 4861 24190 4895
rect 24144 4823 24190 4861
rect 24144 4789 24150 4823
rect 24184 4789 24190 4823
rect 24144 4751 24190 4789
rect 24144 4717 24150 4751
rect 24184 4717 24190 4751
rect 24144 4679 24190 4717
rect 24144 4645 24150 4679
rect 24184 4645 24190 4679
rect 24144 4607 24190 4645
rect 24144 4573 24150 4607
rect 24184 4573 24190 4607
rect 24144 4535 24190 4573
rect 24144 4501 24150 4535
rect 24184 4501 24190 4535
rect 24144 4463 24190 4501
rect 24144 4429 24150 4463
rect 24184 4429 24190 4463
rect 24144 4391 24190 4429
rect 24144 4357 24150 4391
rect 24184 4357 24190 4391
rect 24144 4319 24190 4357
rect 24144 4285 24150 4319
rect 24184 4285 24190 4319
rect 24144 4247 24190 4285
rect 24144 4213 24150 4247
rect 24184 4213 24190 4247
rect 24144 4175 24190 4213
rect 24144 4141 24150 4175
rect 24184 4141 24190 4175
rect 24144 4126 24190 4141
rect 24240 5111 24286 5126
rect 24240 5077 24246 5111
rect 24280 5077 24286 5111
rect 24240 5039 24286 5077
rect 24240 5005 24246 5039
rect 24280 5005 24286 5039
rect 24240 4967 24286 5005
rect 24240 4933 24246 4967
rect 24280 4933 24286 4967
rect 24240 4895 24286 4933
rect 24240 4861 24246 4895
rect 24280 4861 24286 4895
rect 24240 4823 24286 4861
rect 24240 4789 24246 4823
rect 24280 4789 24286 4823
rect 24240 4751 24286 4789
rect 24240 4717 24246 4751
rect 24280 4717 24286 4751
rect 24240 4679 24286 4717
rect 24240 4645 24246 4679
rect 24280 4645 24286 4679
rect 24240 4607 24286 4645
rect 24240 4573 24246 4607
rect 24280 4573 24286 4607
rect 24240 4535 24286 4573
rect 24240 4501 24246 4535
rect 24280 4501 24286 4535
rect 24240 4463 24286 4501
rect 24240 4429 24246 4463
rect 24280 4429 24286 4463
rect 24240 4391 24286 4429
rect 24240 4357 24246 4391
rect 24280 4357 24286 4391
rect 24240 4319 24286 4357
rect 24240 4285 24246 4319
rect 24280 4285 24286 4319
rect 24240 4247 24286 4285
rect 24240 4213 24246 4247
rect 24280 4213 24286 4247
rect 24240 4175 24286 4213
rect 24240 4141 24246 4175
rect 24280 4141 24286 4175
rect 24240 4126 24286 4141
rect 24336 5111 24382 5126
rect 24336 5077 24342 5111
rect 24376 5077 24382 5111
rect 24336 5039 24382 5077
rect 24336 5005 24342 5039
rect 24376 5005 24382 5039
rect 24336 4967 24382 5005
rect 24336 4933 24342 4967
rect 24376 4933 24382 4967
rect 24336 4895 24382 4933
rect 24336 4861 24342 4895
rect 24376 4861 24382 4895
rect 24336 4823 24382 4861
rect 24336 4789 24342 4823
rect 24376 4789 24382 4823
rect 24336 4751 24382 4789
rect 24336 4717 24342 4751
rect 24376 4717 24382 4751
rect 24336 4679 24382 4717
rect 24336 4645 24342 4679
rect 24376 4645 24382 4679
rect 24336 4607 24382 4645
rect 24336 4573 24342 4607
rect 24376 4573 24382 4607
rect 24336 4535 24382 4573
rect 24336 4501 24342 4535
rect 24376 4501 24382 4535
rect 24336 4463 24382 4501
rect 24336 4429 24342 4463
rect 24376 4429 24382 4463
rect 24336 4391 24382 4429
rect 24336 4357 24342 4391
rect 24376 4357 24382 4391
rect 24336 4319 24382 4357
rect 24336 4285 24342 4319
rect 24376 4285 24382 4319
rect 24336 4247 24382 4285
rect 24336 4213 24342 4247
rect 24376 4213 24382 4247
rect 24336 4175 24382 4213
rect 24336 4141 24342 4175
rect 24376 4141 24382 4175
rect 24336 4126 24382 4141
rect 24432 5111 24478 5126
rect 24432 5077 24438 5111
rect 24472 5077 24478 5111
rect 24432 5039 24478 5077
rect 24432 5005 24438 5039
rect 24472 5005 24478 5039
rect 24432 4967 24478 5005
rect 24432 4933 24438 4967
rect 24472 4933 24478 4967
rect 24432 4895 24478 4933
rect 24432 4861 24438 4895
rect 24472 4861 24478 4895
rect 24432 4823 24478 4861
rect 24432 4789 24438 4823
rect 24472 4789 24478 4823
rect 24432 4751 24478 4789
rect 24432 4717 24438 4751
rect 24472 4717 24478 4751
rect 24432 4679 24478 4717
rect 24432 4645 24438 4679
rect 24472 4645 24478 4679
rect 24432 4607 24478 4645
rect 24432 4573 24438 4607
rect 24472 4573 24478 4607
rect 24432 4535 24478 4573
rect 24432 4501 24438 4535
rect 24472 4501 24478 4535
rect 24432 4463 24478 4501
rect 24432 4429 24438 4463
rect 24472 4429 24478 4463
rect 24432 4391 24478 4429
rect 24432 4357 24438 4391
rect 24472 4357 24478 4391
rect 24432 4319 24478 4357
rect 24432 4285 24438 4319
rect 24472 4285 24478 4319
rect 24432 4247 24478 4285
rect 24432 4213 24438 4247
rect 24472 4213 24478 4247
rect 24432 4175 24478 4213
rect 24432 4141 24438 4175
rect 24472 4141 24478 4175
rect 24432 4126 24478 4141
rect 24528 5111 24574 5126
rect 24528 5077 24534 5111
rect 24568 5077 24574 5111
rect 24528 5039 24574 5077
rect 24528 5005 24534 5039
rect 24568 5005 24574 5039
rect 24528 4967 24574 5005
rect 24528 4933 24534 4967
rect 24568 4933 24574 4967
rect 24528 4895 24574 4933
rect 24528 4861 24534 4895
rect 24568 4861 24574 4895
rect 24528 4823 24574 4861
rect 24528 4789 24534 4823
rect 24568 4789 24574 4823
rect 24528 4751 24574 4789
rect 24528 4717 24534 4751
rect 24568 4717 24574 4751
rect 24528 4679 24574 4717
rect 24528 4645 24534 4679
rect 24568 4645 24574 4679
rect 24528 4607 24574 4645
rect 24528 4573 24534 4607
rect 24568 4573 24574 4607
rect 24528 4535 24574 4573
rect 24528 4501 24534 4535
rect 24568 4501 24574 4535
rect 24528 4463 24574 4501
rect 24528 4429 24534 4463
rect 24568 4429 24574 4463
rect 24528 4391 24574 4429
rect 24528 4357 24534 4391
rect 24568 4357 24574 4391
rect 24528 4319 24574 4357
rect 24528 4285 24534 4319
rect 24568 4285 24574 4319
rect 24528 4247 24574 4285
rect 24528 4213 24534 4247
rect 24568 4213 24574 4247
rect 24528 4175 24574 4213
rect 24528 4141 24534 4175
rect 24568 4141 24574 4175
rect 24528 4126 24574 4141
rect 24624 5111 24670 5126
rect 24624 5077 24630 5111
rect 24664 5077 24670 5111
rect 24624 5039 24670 5077
rect 24624 5005 24630 5039
rect 24664 5005 24670 5039
rect 24624 4967 24670 5005
rect 24624 4933 24630 4967
rect 24664 4933 24670 4967
rect 24624 4895 24670 4933
rect 24624 4861 24630 4895
rect 24664 4861 24670 4895
rect 24624 4823 24670 4861
rect 24624 4789 24630 4823
rect 24664 4789 24670 4823
rect 24624 4751 24670 4789
rect 24624 4717 24630 4751
rect 24664 4717 24670 4751
rect 24624 4679 24670 4717
rect 24624 4645 24630 4679
rect 24664 4645 24670 4679
rect 24624 4607 24670 4645
rect 24624 4573 24630 4607
rect 24664 4573 24670 4607
rect 24624 4535 24670 4573
rect 24624 4501 24630 4535
rect 24664 4501 24670 4535
rect 24624 4463 24670 4501
rect 24624 4429 24630 4463
rect 24664 4429 24670 4463
rect 24624 4391 24670 4429
rect 24624 4357 24630 4391
rect 24664 4357 24670 4391
rect 24624 4319 24670 4357
rect 24624 4285 24630 4319
rect 24664 4285 24670 4319
rect 24624 4247 24670 4285
rect 24624 4213 24630 4247
rect 24664 4213 24670 4247
rect 24624 4175 24670 4213
rect 24624 4141 24630 4175
rect 24664 4141 24670 4175
rect 24624 4126 24670 4141
rect 24720 5111 24766 5126
rect 24720 5077 24726 5111
rect 24760 5077 24766 5111
rect 24720 5039 24766 5077
rect 24720 5005 24726 5039
rect 24760 5005 24766 5039
rect 24720 4967 24766 5005
rect 24720 4933 24726 4967
rect 24760 4933 24766 4967
rect 24720 4895 24766 4933
rect 24720 4861 24726 4895
rect 24760 4861 24766 4895
rect 24720 4823 24766 4861
rect 24720 4789 24726 4823
rect 24760 4789 24766 4823
rect 24720 4751 24766 4789
rect 24720 4717 24726 4751
rect 24760 4717 24766 4751
rect 24720 4679 24766 4717
rect 24720 4645 24726 4679
rect 24760 4645 24766 4679
rect 24720 4607 24766 4645
rect 24720 4573 24726 4607
rect 24760 4573 24766 4607
rect 24720 4535 24766 4573
rect 24720 4501 24726 4535
rect 24760 4501 24766 4535
rect 24720 4463 24766 4501
rect 24720 4429 24726 4463
rect 24760 4429 24766 4463
rect 24720 4391 24766 4429
rect 24720 4357 24726 4391
rect 24760 4357 24766 4391
rect 24720 4319 24766 4357
rect 24720 4285 24726 4319
rect 24760 4285 24766 4319
rect 24720 4247 24766 4285
rect 24720 4213 24726 4247
rect 24760 4213 24766 4247
rect 24720 4175 24766 4213
rect 24720 4141 24726 4175
rect 24760 4141 24766 4175
rect 24720 4126 24766 4141
rect 24816 5111 24862 5126
rect 24816 5077 24822 5111
rect 24856 5077 24862 5111
rect 24816 5039 24862 5077
rect 24816 5005 24822 5039
rect 24856 5005 24862 5039
rect 24816 4967 24862 5005
rect 24816 4933 24822 4967
rect 24856 4933 24862 4967
rect 24816 4895 24862 4933
rect 24816 4861 24822 4895
rect 24856 4861 24862 4895
rect 24816 4823 24862 4861
rect 24816 4789 24822 4823
rect 24856 4789 24862 4823
rect 24816 4751 24862 4789
rect 24816 4717 24822 4751
rect 24856 4717 24862 4751
rect 24816 4679 24862 4717
rect 24816 4645 24822 4679
rect 24856 4645 24862 4679
rect 24816 4607 24862 4645
rect 24816 4573 24822 4607
rect 24856 4573 24862 4607
rect 24816 4535 24862 4573
rect 24816 4501 24822 4535
rect 24856 4501 24862 4535
rect 24816 4463 24862 4501
rect 24816 4429 24822 4463
rect 24856 4429 24862 4463
rect 24816 4391 24862 4429
rect 24816 4357 24822 4391
rect 24856 4357 24862 4391
rect 24816 4319 24862 4357
rect 24816 4285 24822 4319
rect 24856 4285 24862 4319
rect 24816 4247 24862 4285
rect 24816 4213 24822 4247
rect 24856 4213 24862 4247
rect 24816 4175 24862 4213
rect 24816 4141 24822 4175
rect 24856 4141 24862 4175
rect 24816 4126 24862 4141
rect 24912 5111 24958 5126
rect 24912 5077 24918 5111
rect 24952 5077 24958 5111
rect 24912 5039 24958 5077
rect 24912 5005 24918 5039
rect 24952 5005 24958 5039
rect 24912 4967 24958 5005
rect 24912 4933 24918 4967
rect 24952 4933 24958 4967
rect 24912 4895 24958 4933
rect 24912 4861 24918 4895
rect 24952 4861 24958 4895
rect 24912 4823 24958 4861
rect 24912 4789 24918 4823
rect 24952 4789 24958 4823
rect 24912 4751 24958 4789
rect 24912 4717 24918 4751
rect 24952 4717 24958 4751
rect 24912 4679 24958 4717
rect 24912 4645 24918 4679
rect 24952 4645 24958 4679
rect 24912 4607 24958 4645
rect 24912 4573 24918 4607
rect 24952 4573 24958 4607
rect 24912 4535 24958 4573
rect 24912 4501 24918 4535
rect 24952 4501 24958 4535
rect 24912 4463 24958 4501
rect 24912 4429 24918 4463
rect 24952 4429 24958 4463
rect 24912 4391 24958 4429
rect 24912 4357 24918 4391
rect 24952 4357 24958 4391
rect 24912 4319 24958 4357
rect 24912 4285 24918 4319
rect 24952 4285 24958 4319
rect 24912 4247 24958 4285
rect 24912 4213 24918 4247
rect 24952 4213 24958 4247
rect 24912 4175 24958 4213
rect 24912 4141 24918 4175
rect 24952 4141 24958 4175
rect 24912 4126 24958 4141
rect 25156 5105 25202 5120
rect 25156 5071 25162 5105
rect 25196 5071 25202 5105
rect 25156 5033 25202 5071
rect 25156 4999 25162 5033
rect 25196 4999 25202 5033
rect 25156 4961 25202 4999
rect 25156 4927 25162 4961
rect 25196 4927 25202 4961
rect 25156 4889 25202 4927
rect 25156 4855 25162 4889
rect 25196 4855 25202 4889
rect 25156 4817 25202 4855
rect 25156 4783 25162 4817
rect 25196 4783 25202 4817
rect 25156 4745 25202 4783
rect 25156 4711 25162 4745
rect 25196 4711 25202 4745
rect 25156 4673 25202 4711
rect 25156 4639 25162 4673
rect 25196 4639 25202 4673
rect 25156 4601 25202 4639
rect 25156 4567 25162 4601
rect 25196 4567 25202 4601
rect 25156 4529 25202 4567
rect 25156 4495 25162 4529
rect 25196 4495 25202 4529
rect 25156 4457 25202 4495
rect 25156 4423 25162 4457
rect 25196 4423 25202 4457
rect 25156 4385 25202 4423
rect 25156 4351 25162 4385
rect 25196 4351 25202 4385
rect 25156 4313 25202 4351
rect 25156 4279 25162 4313
rect 25196 4279 25202 4313
rect 25156 4241 25202 4279
rect 25156 4207 25162 4241
rect 25196 4207 25202 4241
rect 25156 4169 25202 4207
rect 25156 4135 25162 4169
rect 25196 4135 25202 4169
rect 25156 4120 25202 4135
rect 25252 5105 25298 5120
rect 25252 5071 25258 5105
rect 25292 5071 25298 5105
rect 25252 5033 25298 5071
rect 25252 4999 25258 5033
rect 25292 4999 25298 5033
rect 25252 4961 25298 4999
rect 25252 4927 25258 4961
rect 25292 4927 25298 4961
rect 25252 4889 25298 4927
rect 25252 4855 25258 4889
rect 25292 4855 25298 4889
rect 25252 4817 25298 4855
rect 25252 4783 25258 4817
rect 25292 4783 25298 4817
rect 25252 4745 25298 4783
rect 25252 4711 25258 4745
rect 25292 4711 25298 4745
rect 25252 4673 25298 4711
rect 25252 4639 25258 4673
rect 25292 4639 25298 4673
rect 25252 4601 25298 4639
rect 25252 4567 25258 4601
rect 25292 4567 25298 4601
rect 25252 4529 25298 4567
rect 25252 4495 25258 4529
rect 25292 4495 25298 4529
rect 25252 4457 25298 4495
rect 25252 4423 25258 4457
rect 25292 4423 25298 4457
rect 25252 4385 25298 4423
rect 25252 4351 25258 4385
rect 25292 4351 25298 4385
rect 25252 4313 25298 4351
rect 25252 4279 25258 4313
rect 25292 4279 25298 4313
rect 25252 4241 25298 4279
rect 25252 4207 25258 4241
rect 25292 4207 25298 4241
rect 25252 4169 25298 4207
rect 25252 4135 25258 4169
rect 25292 4135 25298 4169
rect 25252 4120 25298 4135
rect 25348 5105 25394 5120
rect 25348 5071 25354 5105
rect 25388 5071 25394 5105
rect 25348 5033 25394 5071
rect 25348 4999 25354 5033
rect 25388 4999 25394 5033
rect 25348 4961 25394 4999
rect 25348 4927 25354 4961
rect 25388 4927 25394 4961
rect 25348 4889 25394 4927
rect 25348 4855 25354 4889
rect 25388 4855 25394 4889
rect 25348 4817 25394 4855
rect 25348 4783 25354 4817
rect 25388 4783 25394 4817
rect 25348 4745 25394 4783
rect 25348 4711 25354 4745
rect 25388 4711 25394 4745
rect 25348 4673 25394 4711
rect 25348 4639 25354 4673
rect 25388 4639 25394 4673
rect 25348 4601 25394 4639
rect 25348 4567 25354 4601
rect 25388 4567 25394 4601
rect 25348 4529 25394 4567
rect 25348 4495 25354 4529
rect 25388 4495 25394 4529
rect 25348 4457 25394 4495
rect 25348 4423 25354 4457
rect 25388 4423 25394 4457
rect 25348 4385 25394 4423
rect 25348 4351 25354 4385
rect 25388 4351 25394 4385
rect 25348 4313 25394 4351
rect 25348 4279 25354 4313
rect 25388 4279 25394 4313
rect 25348 4241 25394 4279
rect 25348 4207 25354 4241
rect 25388 4207 25394 4241
rect 25348 4169 25394 4207
rect 25348 4135 25354 4169
rect 25388 4135 25394 4169
rect 25348 4120 25394 4135
rect 25444 5105 25490 5120
rect 25444 5071 25450 5105
rect 25484 5071 25490 5105
rect 25444 5033 25490 5071
rect 25444 4999 25450 5033
rect 25484 4999 25490 5033
rect 25444 4961 25490 4999
rect 25444 4927 25450 4961
rect 25484 4927 25490 4961
rect 25444 4889 25490 4927
rect 25444 4855 25450 4889
rect 25484 4855 25490 4889
rect 25444 4817 25490 4855
rect 25444 4783 25450 4817
rect 25484 4783 25490 4817
rect 25444 4745 25490 4783
rect 25444 4711 25450 4745
rect 25484 4711 25490 4745
rect 25444 4673 25490 4711
rect 25444 4639 25450 4673
rect 25484 4639 25490 4673
rect 25444 4601 25490 4639
rect 25444 4567 25450 4601
rect 25484 4567 25490 4601
rect 25444 4529 25490 4567
rect 25444 4495 25450 4529
rect 25484 4495 25490 4529
rect 25444 4457 25490 4495
rect 25444 4423 25450 4457
rect 25484 4423 25490 4457
rect 25444 4385 25490 4423
rect 25444 4351 25450 4385
rect 25484 4351 25490 4385
rect 25444 4313 25490 4351
rect 25444 4279 25450 4313
rect 25484 4279 25490 4313
rect 25444 4241 25490 4279
rect 25444 4207 25450 4241
rect 25484 4207 25490 4241
rect 25444 4169 25490 4207
rect 25444 4135 25450 4169
rect 25484 4135 25490 4169
rect 25444 4120 25490 4135
rect 25540 5105 25586 5120
rect 25540 5071 25546 5105
rect 25580 5071 25586 5105
rect 25540 5033 25586 5071
rect 25540 4999 25546 5033
rect 25580 4999 25586 5033
rect 25540 4961 25586 4999
rect 25540 4927 25546 4961
rect 25580 4927 25586 4961
rect 25540 4889 25586 4927
rect 25540 4855 25546 4889
rect 25580 4855 25586 4889
rect 25540 4817 25586 4855
rect 25540 4783 25546 4817
rect 25580 4783 25586 4817
rect 25540 4745 25586 4783
rect 25540 4711 25546 4745
rect 25580 4711 25586 4745
rect 25540 4673 25586 4711
rect 25540 4639 25546 4673
rect 25580 4639 25586 4673
rect 25540 4601 25586 4639
rect 25540 4567 25546 4601
rect 25580 4567 25586 4601
rect 25540 4529 25586 4567
rect 25540 4495 25546 4529
rect 25580 4495 25586 4529
rect 25540 4457 25586 4495
rect 25540 4423 25546 4457
rect 25580 4423 25586 4457
rect 25540 4385 25586 4423
rect 25540 4351 25546 4385
rect 25580 4351 25586 4385
rect 25540 4313 25586 4351
rect 25540 4279 25546 4313
rect 25580 4279 25586 4313
rect 25540 4241 25586 4279
rect 25540 4207 25546 4241
rect 25580 4207 25586 4241
rect 25540 4169 25586 4207
rect 25540 4135 25546 4169
rect 25580 4135 25586 4169
rect 25540 4120 25586 4135
rect 25636 5105 25682 5120
rect 25636 5071 25642 5105
rect 25676 5071 25682 5105
rect 25636 5033 25682 5071
rect 25636 4999 25642 5033
rect 25676 4999 25682 5033
rect 25636 4961 25682 4999
rect 25636 4927 25642 4961
rect 25676 4927 25682 4961
rect 25636 4889 25682 4927
rect 25636 4855 25642 4889
rect 25676 4855 25682 4889
rect 25636 4817 25682 4855
rect 25636 4783 25642 4817
rect 25676 4783 25682 4817
rect 25636 4745 25682 4783
rect 25636 4711 25642 4745
rect 25676 4711 25682 4745
rect 25636 4673 25682 4711
rect 25636 4639 25642 4673
rect 25676 4639 25682 4673
rect 25636 4601 25682 4639
rect 25636 4567 25642 4601
rect 25676 4567 25682 4601
rect 25636 4529 25682 4567
rect 25636 4495 25642 4529
rect 25676 4495 25682 4529
rect 25636 4457 25682 4495
rect 25636 4423 25642 4457
rect 25676 4423 25682 4457
rect 25636 4385 25682 4423
rect 25636 4351 25642 4385
rect 25676 4351 25682 4385
rect 25636 4313 25682 4351
rect 25636 4279 25642 4313
rect 25676 4279 25682 4313
rect 25636 4241 25682 4279
rect 25636 4207 25642 4241
rect 25676 4207 25682 4241
rect 25636 4169 25682 4207
rect 25636 4135 25642 4169
rect 25676 4135 25682 4169
rect 25636 4120 25682 4135
rect 25732 5105 25778 5120
rect 25732 5071 25738 5105
rect 25772 5071 25778 5105
rect 25732 5033 25778 5071
rect 25732 4999 25738 5033
rect 25772 4999 25778 5033
rect 25732 4961 25778 4999
rect 25732 4927 25738 4961
rect 25772 4927 25778 4961
rect 25732 4889 25778 4927
rect 25732 4855 25738 4889
rect 25772 4855 25778 4889
rect 25732 4817 25778 4855
rect 25732 4783 25738 4817
rect 25772 4783 25778 4817
rect 25732 4745 25778 4783
rect 25732 4711 25738 4745
rect 25772 4711 25778 4745
rect 25732 4673 25778 4711
rect 25732 4639 25738 4673
rect 25772 4639 25778 4673
rect 25732 4601 25778 4639
rect 25732 4567 25738 4601
rect 25772 4567 25778 4601
rect 25732 4529 25778 4567
rect 25732 4495 25738 4529
rect 25772 4495 25778 4529
rect 25732 4457 25778 4495
rect 25732 4423 25738 4457
rect 25772 4423 25778 4457
rect 25732 4385 25778 4423
rect 25732 4351 25738 4385
rect 25772 4351 25778 4385
rect 25732 4313 25778 4351
rect 25732 4279 25738 4313
rect 25772 4279 25778 4313
rect 25732 4241 25778 4279
rect 25732 4207 25738 4241
rect 25772 4207 25778 4241
rect 25732 4169 25778 4207
rect 25732 4135 25738 4169
rect 25772 4135 25778 4169
rect 25732 4120 25778 4135
rect 25828 5105 25874 5120
rect 25828 5071 25834 5105
rect 25868 5071 25874 5105
rect 25828 5033 25874 5071
rect 25828 4999 25834 5033
rect 25868 4999 25874 5033
rect 25828 4961 25874 4999
rect 25828 4927 25834 4961
rect 25868 4927 25874 4961
rect 25828 4889 25874 4927
rect 25828 4855 25834 4889
rect 25868 4855 25874 4889
rect 25828 4817 25874 4855
rect 25828 4783 25834 4817
rect 25868 4783 25874 4817
rect 25828 4745 25874 4783
rect 25828 4711 25834 4745
rect 25868 4711 25874 4745
rect 25828 4673 25874 4711
rect 25828 4639 25834 4673
rect 25868 4639 25874 4673
rect 25828 4601 25874 4639
rect 25828 4567 25834 4601
rect 25868 4567 25874 4601
rect 25828 4529 25874 4567
rect 25828 4495 25834 4529
rect 25868 4495 25874 4529
rect 25828 4457 25874 4495
rect 25828 4423 25834 4457
rect 25868 4423 25874 4457
rect 25828 4385 25874 4423
rect 25828 4351 25834 4385
rect 25868 4351 25874 4385
rect 25828 4313 25874 4351
rect 25828 4279 25834 4313
rect 25868 4279 25874 4313
rect 25828 4241 25874 4279
rect 25828 4207 25834 4241
rect 25868 4207 25874 4241
rect 25828 4169 25874 4207
rect 25828 4135 25834 4169
rect 25868 4135 25874 4169
rect 25828 4120 25874 4135
rect 25924 5105 25970 5120
rect 25924 5071 25930 5105
rect 25964 5071 25970 5105
rect 25924 5033 25970 5071
rect 25924 4999 25930 5033
rect 25964 4999 25970 5033
rect 25924 4961 25970 4999
rect 25924 4927 25930 4961
rect 25964 4927 25970 4961
rect 25924 4889 25970 4927
rect 25924 4855 25930 4889
rect 25964 4855 25970 4889
rect 25924 4817 25970 4855
rect 25924 4783 25930 4817
rect 25964 4783 25970 4817
rect 25924 4745 25970 4783
rect 25924 4711 25930 4745
rect 25964 4711 25970 4745
rect 25924 4673 25970 4711
rect 25924 4639 25930 4673
rect 25964 4639 25970 4673
rect 25924 4601 25970 4639
rect 25924 4567 25930 4601
rect 25964 4567 25970 4601
rect 25924 4529 25970 4567
rect 25924 4495 25930 4529
rect 25964 4495 25970 4529
rect 25924 4457 25970 4495
rect 25924 4423 25930 4457
rect 25964 4423 25970 4457
rect 25924 4385 25970 4423
rect 25924 4351 25930 4385
rect 25964 4351 25970 4385
rect 25924 4313 25970 4351
rect 25924 4279 25930 4313
rect 25964 4279 25970 4313
rect 25924 4241 25970 4279
rect 25924 4207 25930 4241
rect 25964 4207 25970 4241
rect 25924 4169 25970 4207
rect 25924 4135 25930 4169
rect 25964 4135 25970 4169
rect 25924 4120 25970 4135
rect 26020 5105 26066 5120
rect 26020 5071 26026 5105
rect 26060 5071 26066 5105
rect 26020 5033 26066 5071
rect 26020 4999 26026 5033
rect 26060 4999 26066 5033
rect 26020 4961 26066 4999
rect 26020 4927 26026 4961
rect 26060 4927 26066 4961
rect 26020 4889 26066 4927
rect 26020 4855 26026 4889
rect 26060 4855 26066 4889
rect 26020 4817 26066 4855
rect 26020 4783 26026 4817
rect 26060 4783 26066 4817
rect 26020 4745 26066 4783
rect 26020 4711 26026 4745
rect 26060 4711 26066 4745
rect 26020 4673 26066 4711
rect 26020 4639 26026 4673
rect 26060 4639 26066 4673
rect 26020 4601 26066 4639
rect 26020 4567 26026 4601
rect 26060 4567 26066 4601
rect 26020 4529 26066 4567
rect 26020 4495 26026 4529
rect 26060 4495 26066 4529
rect 26020 4457 26066 4495
rect 26020 4423 26026 4457
rect 26060 4423 26066 4457
rect 26020 4385 26066 4423
rect 26020 4351 26026 4385
rect 26060 4351 26066 4385
rect 26020 4313 26066 4351
rect 26020 4279 26026 4313
rect 26060 4279 26066 4313
rect 26020 4241 26066 4279
rect 26020 4207 26026 4241
rect 26060 4207 26066 4241
rect 26020 4169 26066 4207
rect 26020 4135 26026 4169
rect 26060 4135 26066 4169
rect 26020 4120 26066 4135
rect 26116 5105 26162 5120
rect 26116 5071 26122 5105
rect 26156 5071 26162 5105
rect 26116 5033 26162 5071
rect 26116 4999 26122 5033
rect 26156 4999 26162 5033
rect 26116 4961 26162 4999
rect 26116 4927 26122 4961
rect 26156 4927 26162 4961
rect 26116 4889 26162 4927
rect 26116 4855 26122 4889
rect 26156 4855 26162 4889
rect 26116 4817 26162 4855
rect 26116 4783 26122 4817
rect 26156 4783 26162 4817
rect 26116 4745 26162 4783
rect 26116 4711 26122 4745
rect 26156 4711 26162 4745
rect 26116 4673 26162 4711
rect 26116 4639 26122 4673
rect 26156 4639 26162 4673
rect 26116 4601 26162 4639
rect 26116 4567 26122 4601
rect 26156 4567 26162 4601
rect 26116 4529 26162 4567
rect 26116 4495 26122 4529
rect 26156 4495 26162 4529
rect 26116 4457 26162 4495
rect 26116 4423 26122 4457
rect 26156 4423 26162 4457
rect 26116 4385 26162 4423
rect 26116 4351 26122 4385
rect 26156 4351 26162 4385
rect 26116 4313 26162 4351
rect 26116 4279 26122 4313
rect 26156 4279 26162 4313
rect 26116 4241 26162 4279
rect 26116 4207 26122 4241
rect 26156 4207 26162 4241
rect 26116 4169 26162 4207
rect 26116 4135 26122 4169
rect 26156 4135 26162 4169
rect 26116 4120 26162 4135
rect 26212 5105 26258 5120
rect 26212 5071 26218 5105
rect 26252 5071 26258 5105
rect 26212 5033 26258 5071
rect 26212 4999 26218 5033
rect 26252 4999 26258 5033
rect 26212 4961 26258 4999
rect 26212 4927 26218 4961
rect 26252 4927 26258 4961
rect 26212 4889 26258 4927
rect 26212 4855 26218 4889
rect 26252 4855 26258 4889
rect 26212 4817 26258 4855
rect 26212 4783 26218 4817
rect 26252 4783 26258 4817
rect 26212 4745 26258 4783
rect 26212 4711 26218 4745
rect 26252 4711 26258 4745
rect 26212 4673 26258 4711
rect 26212 4639 26218 4673
rect 26252 4639 26258 4673
rect 26212 4601 26258 4639
rect 26212 4567 26218 4601
rect 26252 4567 26258 4601
rect 26212 4529 26258 4567
rect 26212 4495 26218 4529
rect 26252 4495 26258 4529
rect 26212 4457 26258 4495
rect 26212 4423 26218 4457
rect 26252 4423 26258 4457
rect 26212 4385 26258 4423
rect 26212 4351 26218 4385
rect 26252 4351 26258 4385
rect 26212 4313 26258 4351
rect 26212 4279 26218 4313
rect 26252 4279 26258 4313
rect 26212 4241 26258 4279
rect 26212 4207 26218 4241
rect 26252 4207 26258 4241
rect 26212 4169 26258 4207
rect 26212 4135 26218 4169
rect 26252 4135 26258 4169
rect 26212 4120 26258 4135
rect 26308 5105 26354 5120
rect 26308 5071 26314 5105
rect 26348 5071 26354 5105
rect 26308 5033 26354 5071
rect 26308 4999 26314 5033
rect 26348 4999 26354 5033
rect 26308 4961 26354 4999
rect 26308 4927 26314 4961
rect 26348 4927 26354 4961
rect 26308 4889 26354 4927
rect 26308 4855 26314 4889
rect 26348 4855 26354 4889
rect 26308 4817 26354 4855
rect 26308 4783 26314 4817
rect 26348 4783 26354 4817
rect 26308 4745 26354 4783
rect 26308 4711 26314 4745
rect 26348 4711 26354 4745
rect 26308 4673 26354 4711
rect 26308 4639 26314 4673
rect 26348 4639 26354 4673
rect 26308 4601 26354 4639
rect 26308 4567 26314 4601
rect 26348 4567 26354 4601
rect 26308 4529 26354 4567
rect 26308 4495 26314 4529
rect 26348 4495 26354 4529
rect 26308 4457 26354 4495
rect 26308 4423 26314 4457
rect 26348 4423 26354 4457
rect 26308 4385 26354 4423
rect 26308 4351 26314 4385
rect 26348 4351 26354 4385
rect 26308 4313 26354 4351
rect 26308 4279 26314 4313
rect 26348 4279 26354 4313
rect 26308 4241 26354 4279
rect 26308 4207 26314 4241
rect 26348 4207 26354 4241
rect 26308 4169 26354 4207
rect 26308 4135 26314 4169
rect 26348 4135 26354 4169
rect 26308 4120 26354 4135
rect 26404 5105 26450 5120
rect 26404 5071 26410 5105
rect 26444 5071 26450 5105
rect 26404 5033 26450 5071
rect 26404 4999 26410 5033
rect 26444 4999 26450 5033
rect 26404 4961 26450 4999
rect 26404 4927 26410 4961
rect 26444 4927 26450 4961
rect 26404 4889 26450 4927
rect 26404 4855 26410 4889
rect 26444 4855 26450 4889
rect 26404 4817 26450 4855
rect 26404 4783 26410 4817
rect 26444 4783 26450 4817
rect 26404 4745 26450 4783
rect 26404 4711 26410 4745
rect 26444 4711 26450 4745
rect 26404 4673 26450 4711
rect 26404 4639 26410 4673
rect 26444 4639 26450 4673
rect 26404 4601 26450 4639
rect 26404 4567 26410 4601
rect 26444 4567 26450 4601
rect 26404 4529 26450 4567
rect 26404 4495 26410 4529
rect 26444 4495 26450 4529
rect 26404 4457 26450 4495
rect 26404 4423 26410 4457
rect 26444 4423 26450 4457
rect 26404 4385 26450 4423
rect 26404 4351 26410 4385
rect 26444 4351 26450 4385
rect 26404 4313 26450 4351
rect 26404 4279 26410 4313
rect 26444 4279 26450 4313
rect 26404 4241 26450 4279
rect 26404 4207 26410 4241
rect 26444 4207 26450 4241
rect 26404 4169 26450 4207
rect 26404 4135 26410 4169
rect 26444 4135 26450 4169
rect 26404 4120 26450 4135
rect 26500 5105 26546 5120
rect 26500 5071 26506 5105
rect 26540 5071 26546 5105
rect 26500 5033 26546 5071
rect 26500 4999 26506 5033
rect 26540 4999 26546 5033
rect 26500 4961 26546 4999
rect 26500 4927 26506 4961
rect 26540 4927 26546 4961
rect 26500 4889 26546 4927
rect 26500 4855 26506 4889
rect 26540 4855 26546 4889
rect 26500 4817 26546 4855
rect 26500 4783 26506 4817
rect 26540 4783 26546 4817
rect 26500 4745 26546 4783
rect 26500 4711 26506 4745
rect 26540 4711 26546 4745
rect 26500 4673 26546 4711
rect 26500 4639 26506 4673
rect 26540 4639 26546 4673
rect 26500 4601 26546 4639
rect 26500 4567 26506 4601
rect 26540 4567 26546 4601
rect 26500 4529 26546 4567
rect 26500 4495 26506 4529
rect 26540 4495 26546 4529
rect 26500 4457 26546 4495
rect 26500 4423 26506 4457
rect 26540 4423 26546 4457
rect 26500 4385 26546 4423
rect 26500 4351 26506 4385
rect 26540 4351 26546 4385
rect 26500 4313 26546 4351
rect 26500 4279 26506 4313
rect 26540 4279 26546 4313
rect 26500 4241 26546 4279
rect 26500 4207 26506 4241
rect 26540 4207 26546 4241
rect 26500 4169 26546 4207
rect 26500 4135 26506 4169
rect 26540 4135 26546 4169
rect 26500 4120 26546 4135
rect 26596 5105 26642 5120
rect 26596 5071 26602 5105
rect 26636 5071 26642 5105
rect 26596 5033 26642 5071
rect 26596 4999 26602 5033
rect 26636 4999 26642 5033
rect 26596 4961 26642 4999
rect 26596 4927 26602 4961
rect 26636 4927 26642 4961
rect 26596 4889 26642 4927
rect 26596 4855 26602 4889
rect 26636 4855 26642 4889
rect 26596 4817 26642 4855
rect 26596 4783 26602 4817
rect 26636 4783 26642 4817
rect 26596 4745 26642 4783
rect 26596 4711 26602 4745
rect 26636 4711 26642 4745
rect 26596 4673 26642 4711
rect 26596 4639 26602 4673
rect 26636 4639 26642 4673
rect 26596 4601 26642 4639
rect 26596 4567 26602 4601
rect 26636 4567 26642 4601
rect 26596 4529 26642 4567
rect 26596 4495 26602 4529
rect 26636 4495 26642 4529
rect 26596 4457 26642 4495
rect 26596 4423 26602 4457
rect 26636 4423 26642 4457
rect 26596 4385 26642 4423
rect 26596 4351 26602 4385
rect 26636 4351 26642 4385
rect 26596 4313 26642 4351
rect 26596 4279 26602 4313
rect 26636 4279 26642 4313
rect 26596 4241 26642 4279
rect 26596 4207 26602 4241
rect 26636 4207 26642 4241
rect 26596 4169 26642 4207
rect 26596 4135 26602 4169
rect 26636 4135 26642 4169
rect 26596 4120 26642 4135
rect 26820 5099 26866 5114
rect 26820 5065 26826 5099
rect 26860 5065 26866 5099
rect 26820 5027 26866 5065
rect 26820 4993 26826 5027
rect 26860 4993 26866 5027
rect 26820 4955 26866 4993
rect 26820 4921 26826 4955
rect 26860 4921 26866 4955
rect 26820 4883 26866 4921
rect 26820 4849 26826 4883
rect 26860 4849 26866 4883
rect 26820 4811 26866 4849
rect 26820 4777 26826 4811
rect 26860 4777 26866 4811
rect 26820 4739 26866 4777
rect 26820 4705 26826 4739
rect 26860 4705 26866 4739
rect 26820 4667 26866 4705
rect 26820 4633 26826 4667
rect 26860 4633 26866 4667
rect 26820 4595 26866 4633
rect 26820 4561 26826 4595
rect 26860 4561 26866 4595
rect 26820 4523 26866 4561
rect 26820 4489 26826 4523
rect 26860 4489 26866 4523
rect 26820 4451 26866 4489
rect 26820 4417 26826 4451
rect 26860 4417 26866 4451
rect 26820 4379 26866 4417
rect 26820 4345 26826 4379
rect 26860 4345 26866 4379
rect 26820 4307 26866 4345
rect 26820 4273 26826 4307
rect 26860 4273 26866 4307
rect 26820 4235 26866 4273
rect 26820 4201 26826 4235
rect 26860 4201 26866 4235
rect 26820 4163 26866 4201
rect 26820 4129 26826 4163
rect 26860 4129 26866 4163
rect 26820 4114 26866 4129
rect 26916 5099 26962 5114
rect 26916 5065 26922 5099
rect 26956 5065 26962 5099
rect 26916 5027 26962 5065
rect 26916 4993 26922 5027
rect 26956 4993 26962 5027
rect 26916 4955 26962 4993
rect 26916 4921 26922 4955
rect 26956 4921 26962 4955
rect 26916 4883 26962 4921
rect 26916 4849 26922 4883
rect 26956 4849 26962 4883
rect 26916 4811 26962 4849
rect 26916 4777 26922 4811
rect 26956 4777 26962 4811
rect 26916 4739 26962 4777
rect 26916 4705 26922 4739
rect 26956 4705 26962 4739
rect 26916 4667 26962 4705
rect 26916 4633 26922 4667
rect 26956 4633 26962 4667
rect 26916 4595 26962 4633
rect 26916 4561 26922 4595
rect 26956 4561 26962 4595
rect 26916 4523 26962 4561
rect 26916 4489 26922 4523
rect 26956 4489 26962 4523
rect 26916 4451 26962 4489
rect 26916 4417 26922 4451
rect 26956 4417 26962 4451
rect 26916 4379 26962 4417
rect 26916 4345 26922 4379
rect 26956 4345 26962 4379
rect 26916 4307 26962 4345
rect 26916 4273 26922 4307
rect 26956 4273 26962 4307
rect 26916 4235 26962 4273
rect 26916 4201 26922 4235
rect 26956 4201 26962 4235
rect 26916 4163 26962 4201
rect 26916 4129 26922 4163
rect 26956 4129 26962 4163
rect 26916 4114 26962 4129
rect 27012 5099 27058 5114
rect 27012 5065 27018 5099
rect 27052 5065 27058 5099
rect 27012 5027 27058 5065
rect 27012 4993 27018 5027
rect 27052 4993 27058 5027
rect 27012 4955 27058 4993
rect 27012 4921 27018 4955
rect 27052 4921 27058 4955
rect 27012 4883 27058 4921
rect 27012 4849 27018 4883
rect 27052 4849 27058 4883
rect 27012 4811 27058 4849
rect 27012 4777 27018 4811
rect 27052 4777 27058 4811
rect 27012 4739 27058 4777
rect 27012 4705 27018 4739
rect 27052 4705 27058 4739
rect 27012 4667 27058 4705
rect 27012 4633 27018 4667
rect 27052 4633 27058 4667
rect 27012 4595 27058 4633
rect 27012 4561 27018 4595
rect 27052 4561 27058 4595
rect 27012 4523 27058 4561
rect 27012 4489 27018 4523
rect 27052 4489 27058 4523
rect 27012 4451 27058 4489
rect 27012 4417 27018 4451
rect 27052 4417 27058 4451
rect 27012 4379 27058 4417
rect 27012 4345 27018 4379
rect 27052 4345 27058 4379
rect 27012 4307 27058 4345
rect 27012 4273 27018 4307
rect 27052 4273 27058 4307
rect 27012 4235 27058 4273
rect 27012 4201 27018 4235
rect 27052 4201 27058 4235
rect 27012 4163 27058 4201
rect 27012 4129 27018 4163
rect 27052 4129 27058 4163
rect 27012 4114 27058 4129
rect 27108 5099 27154 5114
rect 27108 5065 27114 5099
rect 27148 5065 27154 5099
rect 27108 5027 27154 5065
rect 27108 4993 27114 5027
rect 27148 4993 27154 5027
rect 27108 4955 27154 4993
rect 27108 4921 27114 4955
rect 27148 4921 27154 4955
rect 27108 4883 27154 4921
rect 27108 4849 27114 4883
rect 27148 4849 27154 4883
rect 27108 4811 27154 4849
rect 27108 4777 27114 4811
rect 27148 4777 27154 4811
rect 27108 4739 27154 4777
rect 27108 4705 27114 4739
rect 27148 4705 27154 4739
rect 27108 4667 27154 4705
rect 27108 4633 27114 4667
rect 27148 4633 27154 4667
rect 27108 4595 27154 4633
rect 27108 4561 27114 4595
rect 27148 4561 27154 4595
rect 27108 4523 27154 4561
rect 27108 4489 27114 4523
rect 27148 4489 27154 4523
rect 27108 4451 27154 4489
rect 27108 4417 27114 4451
rect 27148 4417 27154 4451
rect 27108 4379 27154 4417
rect 27108 4345 27114 4379
rect 27148 4345 27154 4379
rect 27108 4307 27154 4345
rect 27108 4273 27114 4307
rect 27148 4273 27154 4307
rect 27108 4235 27154 4273
rect 27108 4201 27114 4235
rect 27148 4201 27154 4235
rect 27108 4163 27154 4201
rect 27108 4129 27114 4163
rect 27148 4129 27154 4163
rect 27108 4114 27154 4129
rect 27204 5099 27250 5114
rect 27204 5065 27210 5099
rect 27244 5065 27250 5099
rect 27204 5027 27250 5065
rect 27204 4993 27210 5027
rect 27244 4993 27250 5027
rect 27204 4955 27250 4993
rect 27204 4921 27210 4955
rect 27244 4921 27250 4955
rect 27204 4883 27250 4921
rect 27204 4849 27210 4883
rect 27244 4849 27250 4883
rect 27204 4811 27250 4849
rect 27204 4777 27210 4811
rect 27244 4777 27250 4811
rect 27204 4739 27250 4777
rect 27204 4705 27210 4739
rect 27244 4705 27250 4739
rect 27204 4667 27250 4705
rect 27204 4633 27210 4667
rect 27244 4633 27250 4667
rect 27204 4595 27250 4633
rect 27204 4561 27210 4595
rect 27244 4561 27250 4595
rect 27204 4523 27250 4561
rect 27204 4489 27210 4523
rect 27244 4489 27250 4523
rect 27204 4451 27250 4489
rect 27204 4417 27210 4451
rect 27244 4417 27250 4451
rect 27204 4379 27250 4417
rect 27204 4345 27210 4379
rect 27244 4345 27250 4379
rect 27204 4307 27250 4345
rect 27204 4273 27210 4307
rect 27244 4273 27250 4307
rect 27204 4235 27250 4273
rect 27204 4201 27210 4235
rect 27244 4201 27250 4235
rect 27204 4163 27250 4201
rect 27204 4129 27210 4163
rect 27244 4129 27250 4163
rect 27204 4114 27250 4129
rect 27300 5099 27346 5114
rect 27300 5065 27306 5099
rect 27340 5065 27346 5099
rect 27300 5027 27346 5065
rect 27300 4993 27306 5027
rect 27340 4993 27346 5027
rect 27300 4955 27346 4993
rect 27300 4921 27306 4955
rect 27340 4921 27346 4955
rect 27300 4883 27346 4921
rect 27300 4849 27306 4883
rect 27340 4849 27346 4883
rect 27300 4811 27346 4849
rect 27300 4777 27306 4811
rect 27340 4777 27346 4811
rect 27300 4739 27346 4777
rect 27300 4705 27306 4739
rect 27340 4705 27346 4739
rect 27300 4667 27346 4705
rect 27300 4633 27306 4667
rect 27340 4633 27346 4667
rect 27300 4595 27346 4633
rect 27300 4561 27306 4595
rect 27340 4561 27346 4595
rect 27300 4523 27346 4561
rect 27300 4489 27306 4523
rect 27340 4489 27346 4523
rect 27300 4451 27346 4489
rect 27300 4417 27306 4451
rect 27340 4417 27346 4451
rect 27300 4379 27346 4417
rect 27300 4345 27306 4379
rect 27340 4345 27346 4379
rect 27300 4307 27346 4345
rect 27300 4273 27306 4307
rect 27340 4273 27346 4307
rect 27300 4235 27346 4273
rect 27300 4201 27306 4235
rect 27340 4201 27346 4235
rect 27300 4163 27346 4201
rect 27300 4129 27306 4163
rect 27340 4129 27346 4163
rect 27300 4114 27346 4129
rect 27396 5099 27442 5114
rect 27396 5065 27402 5099
rect 27436 5065 27442 5099
rect 27396 5027 27442 5065
rect 27396 4993 27402 5027
rect 27436 4993 27442 5027
rect 27396 4955 27442 4993
rect 27396 4921 27402 4955
rect 27436 4921 27442 4955
rect 27396 4883 27442 4921
rect 27396 4849 27402 4883
rect 27436 4849 27442 4883
rect 27396 4811 27442 4849
rect 27396 4777 27402 4811
rect 27436 4777 27442 4811
rect 27396 4739 27442 4777
rect 27396 4705 27402 4739
rect 27436 4705 27442 4739
rect 27396 4667 27442 4705
rect 27396 4633 27402 4667
rect 27436 4633 27442 4667
rect 27396 4595 27442 4633
rect 27396 4561 27402 4595
rect 27436 4561 27442 4595
rect 27396 4523 27442 4561
rect 27396 4489 27402 4523
rect 27436 4489 27442 4523
rect 27396 4451 27442 4489
rect 27396 4417 27402 4451
rect 27436 4417 27442 4451
rect 27396 4379 27442 4417
rect 27396 4345 27402 4379
rect 27436 4345 27442 4379
rect 27396 4307 27442 4345
rect 27396 4273 27402 4307
rect 27436 4273 27442 4307
rect 27396 4235 27442 4273
rect 27396 4201 27402 4235
rect 27436 4201 27442 4235
rect 27396 4163 27442 4201
rect 27396 4129 27402 4163
rect 27436 4129 27442 4163
rect 27396 4114 27442 4129
rect 27492 5099 27538 5114
rect 27492 5065 27498 5099
rect 27532 5065 27538 5099
rect 27492 5027 27538 5065
rect 27492 4993 27498 5027
rect 27532 4993 27538 5027
rect 27492 4955 27538 4993
rect 27492 4921 27498 4955
rect 27532 4921 27538 4955
rect 27492 4883 27538 4921
rect 27492 4849 27498 4883
rect 27532 4849 27538 4883
rect 27492 4811 27538 4849
rect 27492 4777 27498 4811
rect 27532 4777 27538 4811
rect 27492 4739 27538 4777
rect 27492 4705 27498 4739
rect 27532 4705 27538 4739
rect 27492 4667 27538 4705
rect 27492 4633 27498 4667
rect 27532 4633 27538 4667
rect 27492 4595 27538 4633
rect 27492 4561 27498 4595
rect 27532 4561 27538 4595
rect 27492 4523 27538 4561
rect 27492 4489 27498 4523
rect 27532 4489 27538 4523
rect 27492 4451 27538 4489
rect 27492 4417 27498 4451
rect 27532 4417 27538 4451
rect 27492 4379 27538 4417
rect 27492 4345 27498 4379
rect 27532 4345 27538 4379
rect 27492 4307 27538 4345
rect 27492 4273 27498 4307
rect 27532 4273 27538 4307
rect 27492 4235 27538 4273
rect 27492 4201 27498 4235
rect 27532 4201 27538 4235
rect 27492 4163 27538 4201
rect 27492 4129 27498 4163
rect 27532 4129 27538 4163
rect 27492 4114 27538 4129
rect 27588 5099 27634 5114
rect 27588 5065 27594 5099
rect 27628 5065 27634 5099
rect 27588 5027 27634 5065
rect 27588 4993 27594 5027
rect 27628 4993 27634 5027
rect 27588 4955 27634 4993
rect 27588 4921 27594 4955
rect 27628 4921 27634 4955
rect 27588 4883 27634 4921
rect 27588 4849 27594 4883
rect 27628 4849 27634 4883
rect 27588 4811 27634 4849
rect 27588 4777 27594 4811
rect 27628 4777 27634 4811
rect 27588 4739 27634 4777
rect 27588 4705 27594 4739
rect 27628 4705 27634 4739
rect 27588 4667 27634 4705
rect 27588 4633 27594 4667
rect 27628 4633 27634 4667
rect 27588 4595 27634 4633
rect 27588 4561 27594 4595
rect 27628 4561 27634 4595
rect 27588 4523 27634 4561
rect 27588 4489 27594 4523
rect 27628 4489 27634 4523
rect 27588 4451 27634 4489
rect 27588 4417 27594 4451
rect 27628 4417 27634 4451
rect 27588 4379 27634 4417
rect 27588 4345 27594 4379
rect 27628 4345 27634 4379
rect 27588 4307 27634 4345
rect 27588 4273 27594 4307
rect 27628 4273 27634 4307
rect 27588 4235 27634 4273
rect 27588 4201 27594 4235
rect 27628 4201 27634 4235
rect 27588 4163 27634 4201
rect 27588 4129 27594 4163
rect 27628 4129 27634 4163
rect 27588 4114 27634 4129
rect 27684 5099 27730 5114
rect 27684 5065 27690 5099
rect 27724 5065 27730 5099
rect 27684 5027 27730 5065
rect 27684 4993 27690 5027
rect 27724 4993 27730 5027
rect 27684 4955 27730 4993
rect 27684 4921 27690 4955
rect 27724 4921 27730 4955
rect 27684 4883 27730 4921
rect 27684 4849 27690 4883
rect 27724 4849 27730 4883
rect 27684 4811 27730 4849
rect 27684 4777 27690 4811
rect 27724 4777 27730 4811
rect 27684 4739 27730 4777
rect 27684 4705 27690 4739
rect 27724 4705 27730 4739
rect 27684 4667 27730 4705
rect 27684 4633 27690 4667
rect 27724 4633 27730 4667
rect 27684 4595 27730 4633
rect 27684 4561 27690 4595
rect 27724 4561 27730 4595
rect 27684 4523 27730 4561
rect 27684 4489 27690 4523
rect 27724 4489 27730 4523
rect 27684 4451 27730 4489
rect 27684 4417 27690 4451
rect 27724 4417 27730 4451
rect 27684 4379 27730 4417
rect 27684 4345 27690 4379
rect 27724 4345 27730 4379
rect 27684 4307 27730 4345
rect 27684 4273 27690 4307
rect 27724 4273 27730 4307
rect 27684 4235 27730 4273
rect 27684 4201 27690 4235
rect 27724 4201 27730 4235
rect 27684 4163 27730 4201
rect 27684 4129 27690 4163
rect 27724 4129 27730 4163
rect 27684 4114 27730 4129
rect 27780 5099 27826 5114
rect 27780 5065 27786 5099
rect 27820 5065 27826 5099
rect 27780 5027 27826 5065
rect 27780 4993 27786 5027
rect 27820 4993 27826 5027
rect 27780 4955 27826 4993
rect 27780 4921 27786 4955
rect 27820 4921 27826 4955
rect 27780 4883 27826 4921
rect 27780 4849 27786 4883
rect 27820 4849 27826 4883
rect 27780 4811 27826 4849
rect 27780 4777 27786 4811
rect 27820 4777 27826 4811
rect 27780 4739 27826 4777
rect 27780 4705 27786 4739
rect 27820 4705 27826 4739
rect 27780 4667 27826 4705
rect 27780 4633 27786 4667
rect 27820 4633 27826 4667
rect 27780 4595 27826 4633
rect 27780 4561 27786 4595
rect 27820 4561 27826 4595
rect 27780 4523 27826 4561
rect 27780 4489 27786 4523
rect 27820 4489 27826 4523
rect 27780 4451 27826 4489
rect 27780 4417 27786 4451
rect 27820 4417 27826 4451
rect 27780 4379 27826 4417
rect 27780 4345 27786 4379
rect 27820 4345 27826 4379
rect 27780 4307 27826 4345
rect 27780 4273 27786 4307
rect 27820 4273 27826 4307
rect 27780 4235 27826 4273
rect 27780 4201 27786 4235
rect 27820 4201 27826 4235
rect 27780 4163 27826 4201
rect 27780 4129 27786 4163
rect 27820 4129 27826 4163
rect 27780 4114 27826 4129
rect 27876 5099 27922 5114
rect 27876 5065 27882 5099
rect 27916 5065 27922 5099
rect 27876 5027 27922 5065
rect 27876 4993 27882 5027
rect 27916 4993 27922 5027
rect 27876 4955 27922 4993
rect 27876 4921 27882 4955
rect 27916 4921 27922 4955
rect 27876 4883 27922 4921
rect 27876 4849 27882 4883
rect 27916 4849 27922 4883
rect 27876 4811 27922 4849
rect 27876 4777 27882 4811
rect 27916 4777 27922 4811
rect 27876 4739 27922 4777
rect 27876 4705 27882 4739
rect 27916 4705 27922 4739
rect 27876 4667 27922 4705
rect 27876 4633 27882 4667
rect 27916 4633 27922 4667
rect 27876 4595 27922 4633
rect 27876 4561 27882 4595
rect 27916 4561 27922 4595
rect 27876 4523 27922 4561
rect 27876 4489 27882 4523
rect 27916 4489 27922 4523
rect 27876 4451 27922 4489
rect 27876 4417 27882 4451
rect 27916 4417 27922 4451
rect 27876 4379 27922 4417
rect 27876 4345 27882 4379
rect 27916 4345 27922 4379
rect 27876 4307 27922 4345
rect 27876 4273 27882 4307
rect 27916 4273 27922 4307
rect 27876 4235 27922 4273
rect 27876 4201 27882 4235
rect 27916 4201 27922 4235
rect 27876 4163 27922 4201
rect 27876 4129 27882 4163
rect 27916 4129 27922 4163
rect 27876 4114 27922 4129
rect 27972 5099 28018 5114
rect 27972 5065 27978 5099
rect 28012 5065 28018 5099
rect 27972 5027 28018 5065
rect 27972 4993 27978 5027
rect 28012 4993 28018 5027
rect 27972 4955 28018 4993
rect 27972 4921 27978 4955
rect 28012 4921 28018 4955
rect 27972 4883 28018 4921
rect 27972 4849 27978 4883
rect 28012 4849 28018 4883
rect 27972 4811 28018 4849
rect 27972 4777 27978 4811
rect 28012 4777 28018 4811
rect 27972 4739 28018 4777
rect 27972 4705 27978 4739
rect 28012 4705 28018 4739
rect 27972 4667 28018 4705
rect 27972 4633 27978 4667
rect 28012 4633 28018 4667
rect 27972 4595 28018 4633
rect 27972 4561 27978 4595
rect 28012 4561 28018 4595
rect 27972 4523 28018 4561
rect 27972 4489 27978 4523
rect 28012 4489 28018 4523
rect 27972 4451 28018 4489
rect 27972 4417 27978 4451
rect 28012 4417 28018 4451
rect 27972 4379 28018 4417
rect 27972 4345 27978 4379
rect 28012 4345 28018 4379
rect 27972 4307 28018 4345
rect 27972 4273 27978 4307
rect 28012 4273 28018 4307
rect 27972 4235 28018 4273
rect 27972 4201 27978 4235
rect 28012 4201 28018 4235
rect 27972 4163 28018 4201
rect 27972 4129 27978 4163
rect 28012 4129 28018 4163
rect 27972 4114 28018 4129
rect 28068 5099 28114 5114
rect 28068 5065 28074 5099
rect 28108 5065 28114 5099
rect 28068 5027 28114 5065
rect 28068 4993 28074 5027
rect 28108 4993 28114 5027
rect 28068 4955 28114 4993
rect 28068 4921 28074 4955
rect 28108 4921 28114 4955
rect 28068 4883 28114 4921
rect 28068 4849 28074 4883
rect 28108 4849 28114 4883
rect 28068 4811 28114 4849
rect 28068 4777 28074 4811
rect 28108 4777 28114 4811
rect 28068 4739 28114 4777
rect 28068 4705 28074 4739
rect 28108 4705 28114 4739
rect 28068 4667 28114 4705
rect 28068 4633 28074 4667
rect 28108 4633 28114 4667
rect 28068 4595 28114 4633
rect 28068 4561 28074 4595
rect 28108 4561 28114 4595
rect 28068 4523 28114 4561
rect 28068 4489 28074 4523
rect 28108 4489 28114 4523
rect 28068 4451 28114 4489
rect 28068 4417 28074 4451
rect 28108 4417 28114 4451
rect 28068 4379 28114 4417
rect 28068 4345 28074 4379
rect 28108 4345 28114 4379
rect 28068 4307 28114 4345
rect 28068 4273 28074 4307
rect 28108 4273 28114 4307
rect 28068 4235 28114 4273
rect 28068 4201 28074 4235
rect 28108 4201 28114 4235
rect 28068 4163 28114 4201
rect 28068 4129 28074 4163
rect 28108 4129 28114 4163
rect 28068 4114 28114 4129
rect 28164 5099 28210 5114
rect 28164 5065 28170 5099
rect 28204 5065 28210 5099
rect 28164 5027 28210 5065
rect 28164 4993 28170 5027
rect 28204 4993 28210 5027
rect 28164 4955 28210 4993
rect 28164 4921 28170 4955
rect 28204 4921 28210 4955
rect 28164 4883 28210 4921
rect 28164 4849 28170 4883
rect 28204 4849 28210 4883
rect 28164 4811 28210 4849
rect 28164 4777 28170 4811
rect 28204 4777 28210 4811
rect 28164 4739 28210 4777
rect 28164 4705 28170 4739
rect 28204 4705 28210 4739
rect 28164 4667 28210 4705
rect 28164 4633 28170 4667
rect 28204 4633 28210 4667
rect 28164 4595 28210 4633
rect 28164 4561 28170 4595
rect 28204 4561 28210 4595
rect 28164 4523 28210 4561
rect 28164 4489 28170 4523
rect 28204 4489 28210 4523
rect 28164 4451 28210 4489
rect 28164 4417 28170 4451
rect 28204 4417 28210 4451
rect 28164 4379 28210 4417
rect 28164 4345 28170 4379
rect 28204 4345 28210 4379
rect 28164 4307 28210 4345
rect 28164 4273 28170 4307
rect 28204 4273 28210 4307
rect 28164 4235 28210 4273
rect 28164 4201 28170 4235
rect 28204 4201 28210 4235
rect 28164 4163 28210 4201
rect 28164 4129 28170 4163
rect 28204 4129 28210 4163
rect 28164 4114 28210 4129
rect 28260 5099 28306 5114
rect 28260 5065 28266 5099
rect 28300 5065 28306 5099
rect 28260 5027 28306 5065
rect 28260 4993 28266 5027
rect 28300 4993 28306 5027
rect 28260 4955 28306 4993
rect 28260 4921 28266 4955
rect 28300 4921 28306 4955
rect 28260 4883 28306 4921
rect 28260 4849 28266 4883
rect 28300 4849 28306 4883
rect 28260 4811 28306 4849
rect 28260 4777 28266 4811
rect 28300 4777 28306 4811
rect 28260 4739 28306 4777
rect 28260 4705 28266 4739
rect 28300 4705 28306 4739
rect 28260 4667 28306 4705
rect 28260 4633 28266 4667
rect 28300 4633 28306 4667
rect 28260 4595 28306 4633
rect 28260 4561 28266 4595
rect 28300 4561 28306 4595
rect 28260 4523 28306 4561
rect 28260 4489 28266 4523
rect 28300 4489 28306 4523
rect 28260 4451 28306 4489
rect 28260 4417 28266 4451
rect 28300 4417 28306 4451
rect 28260 4379 28306 4417
rect 28260 4345 28266 4379
rect 28300 4345 28306 4379
rect 28260 4307 28306 4345
rect 28260 4273 28266 4307
rect 28300 4273 28306 4307
rect 28260 4235 28306 4273
rect 28260 4201 28266 4235
rect 28300 4201 28306 4235
rect 28260 4163 28306 4201
rect 28260 4129 28266 4163
rect 28300 4129 28306 4163
rect 28260 4114 28306 4129
rect 28356 5099 28402 5114
rect 28356 5065 28362 5099
rect 28396 5065 28402 5099
rect 28356 5027 28402 5065
rect 28356 4993 28362 5027
rect 28396 4993 28402 5027
rect 28356 4955 28402 4993
rect 28356 4921 28362 4955
rect 28396 4921 28402 4955
rect 28356 4883 28402 4921
rect 28356 4849 28362 4883
rect 28396 4849 28402 4883
rect 28356 4811 28402 4849
rect 28356 4777 28362 4811
rect 28396 4777 28402 4811
rect 28356 4739 28402 4777
rect 28356 4705 28362 4739
rect 28396 4705 28402 4739
rect 28356 4667 28402 4705
rect 28356 4633 28362 4667
rect 28396 4633 28402 4667
rect 28356 4595 28402 4633
rect 28356 4561 28362 4595
rect 28396 4561 28402 4595
rect 28356 4523 28402 4561
rect 28356 4489 28362 4523
rect 28396 4489 28402 4523
rect 28356 4451 28402 4489
rect 28356 4417 28362 4451
rect 28396 4417 28402 4451
rect 28356 4379 28402 4417
rect 28356 4345 28362 4379
rect 28396 4345 28402 4379
rect 28356 4307 28402 4345
rect 28356 4273 28362 4307
rect 28396 4273 28402 4307
rect 28356 4235 28402 4273
rect 28356 4201 28362 4235
rect 28396 4201 28402 4235
rect 28356 4163 28402 4201
rect 28356 4129 28362 4163
rect 28396 4129 28402 4163
rect 28356 4114 28402 4129
rect 28452 5099 28498 5114
rect 28452 5065 28458 5099
rect 28492 5065 28498 5099
rect 28452 5027 28498 5065
rect 28452 4993 28458 5027
rect 28492 4993 28498 5027
rect 28452 4955 28498 4993
rect 28452 4921 28458 4955
rect 28492 4921 28498 4955
rect 28452 4883 28498 4921
rect 28452 4849 28458 4883
rect 28492 4849 28498 4883
rect 28452 4811 28498 4849
rect 28452 4777 28458 4811
rect 28492 4777 28498 4811
rect 28452 4739 28498 4777
rect 28452 4705 28458 4739
rect 28492 4705 28498 4739
rect 28452 4667 28498 4705
rect 28452 4633 28458 4667
rect 28492 4633 28498 4667
rect 28452 4595 28498 4633
rect 28452 4561 28458 4595
rect 28492 4561 28498 4595
rect 28452 4523 28498 4561
rect 28452 4489 28458 4523
rect 28492 4489 28498 4523
rect 28452 4451 28498 4489
rect 28452 4417 28458 4451
rect 28492 4417 28498 4451
rect 28452 4379 28498 4417
rect 28452 4345 28458 4379
rect 28492 4345 28498 4379
rect 28452 4307 28498 4345
rect 28452 4273 28458 4307
rect 28492 4273 28498 4307
rect 28452 4235 28498 4273
rect 28452 4201 28458 4235
rect 28492 4201 28498 4235
rect 28452 4163 28498 4201
rect 28452 4129 28458 4163
rect 28492 4129 28498 4163
rect 28452 4114 28498 4129
rect 28548 5099 28594 5114
rect 28548 5065 28554 5099
rect 28588 5065 28594 5099
rect 28548 5027 28594 5065
rect 28548 4993 28554 5027
rect 28588 4993 28594 5027
rect 28548 4955 28594 4993
rect 28548 4921 28554 4955
rect 28588 4921 28594 4955
rect 28548 4883 28594 4921
rect 28548 4849 28554 4883
rect 28588 4849 28594 4883
rect 28548 4811 28594 4849
rect 28548 4777 28554 4811
rect 28588 4777 28594 4811
rect 28548 4739 28594 4777
rect 28548 4705 28554 4739
rect 28588 4705 28594 4739
rect 28548 4667 28594 4705
rect 28548 4633 28554 4667
rect 28588 4633 28594 4667
rect 28548 4595 28594 4633
rect 28548 4561 28554 4595
rect 28588 4561 28594 4595
rect 28548 4523 28594 4561
rect 28548 4489 28554 4523
rect 28588 4489 28594 4523
rect 28548 4451 28594 4489
rect 28548 4417 28554 4451
rect 28588 4417 28594 4451
rect 28548 4379 28594 4417
rect 28548 4345 28554 4379
rect 28588 4345 28594 4379
rect 28548 4307 28594 4345
rect 28548 4273 28554 4307
rect 28588 4273 28594 4307
rect 28548 4235 28594 4273
rect 28548 4201 28554 4235
rect 28588 4201 28594 4235
rect 28548 4163 28594 4201
rect 28548 4129 28554 4163
rect 28588 4129 28594 4163
rect 28548 4114 28594 4129
rect 28644 5099 28690 5114
rect 28644 5065 28650 5099
rect 28684 5065 28690 5099
rect 28644 5027 28690 5065
rect 28644 4993 28650 5027
rect 28684 4993 28690 5027
rect 28644 4955 28690 4993
rect 28644 4921 28650 4955
rect 28684 4921 28690 4955
rect 28644 4883 28690 4921
rect 28644 4849 28650 4883
rect 28684 4849 28690 4883
rect 28644 4811 28690 4849
rect 28644 4777 28650 4811
rect 28684 4777 28690 4811
rect 28644 4739 28690 4777
rect 28644 4705 28650 4739
rect 28684 4705 28690 4739
rect 28644 4667 28690 4705
rect 28644 4633 28650 4667
rect 28684 4633 28690 4667
rect 28644 4595 28690 4633
rect 28644 4561 28650 4595
rect 28684 4561 28690 4595
rect 28644 4523 28690 4561
rect 28644 4489 28650 4523
rect 28684 4489 28690 4523
rect 28644 4451 28690 4489
rect 28644 4417 28650 4451
rect 28684 4417 28690 4451
rect 28644 4379 28690 4417
rect 28644 4345 28650 4379
rect 28684 4345 28690 4379
rect 28644 4307 28690 4345
rect 28644 4273 28650 4307
rect 28684 4273 28690 4307
rect 28644 4235 28690 4273
rect 28644 4201 28650 4235
rect 28684 4201 28690 4235
rect 28644 4163 28690 4201
rect 28644 4129 28650 4163
rect 28684 4129 28690 4163
rect 28644 4114 28690 4129
rect 28740 5099 28786 5114
rect 28740 5065 28746 5099
rect 28780 5065 28786 5099
rect 28740 5027 28786 5065
rect 28740 4993 28746 5027
rect 28780 4993 28786 5027
rect 28740 4955 28786 4993
rect 28740 4921 28746 4955
rect 28780 4921 28786 4955
rect 28740 4883 28786 4921
rect 28740 4849 28746 4883
rect 28780 4849 28786 4883
rect 28740 4811 28786 4849
rect 28740 4777 28746 4811
rect 28780 4777 28786 4811
rect 28740 4739 28786 4777
rect 28740 4705 28746 4739
rect 28780 4705 28786 4739
rect 28740 4667 28786 4705
rect 28740 4633 28746 4667
rect 28780 4633 28786 4667
rect 28740 4595 28786 4633
rect 28740 4561 28746 4595
rect 28780 4561 28786 4595
rect 28740 4523 28786 4561
rect 28740 4489 28746 4523
rect 28780 4489 28786 4523
rect 28740 4451 28786 4489
rect 28740 4417 28746 4451
rect 28780 4417 28786 4451
rect 28740 4379 28786 4417
rect 28740 4345 28746 4379
rect 28780 4345 28786 4379
rect 28740 4307 28786 4345
rect 28740 4273 28746 4307
rect 28780 4273 28786 4307
rect 28740 4235 28786 4273
rect 28740 4201 28746 4235
rect 28780 4201 28786 4235
rect 28740 4163 28786 4201
rect 28740 4129 28746 4163
rect 28780 4129 28786 4163
rect 28740 4114 28786 4129
rect 15704 4045 15710 4079
rect 15744 4045 15750 4079
rect 15704 4007 15750 4045
rect 15704 3973 15710 4007
rect 15744 3973 15750 4007
rect 15704 3926 15750 3973
rect 16796 3943 16894 3970
rect 14092 3900 14138 3915
rect 16796 3909 16830 3943
rect 16864 3909 16894 3943
rect 16796 3846 16894 3909
rect 16456 3820 16894 3846
rect 17498 3961 17578 3992
rect 17498 3927 17518 3961
rect 17552 3927 17578 3961
rect 17498 3840 17578 3927
rect 18688 3955 18788 3986
rect 18688 3921 18722 3955
rect 18756 3921 18788 3955
rect 18688 3850 18788 3921
rect 1842 3790 2168 3792
rect 1566 3783 1624 3788
rect 1760 3787 2168 3790
rect 1566 3777 1626 3783
rect 1566 3743 1580 3777
rect 1614 3743 1626 3777
rect 1760 3777 2101 3787
rect 1566 3737 1626 3743
rect 1662 3754 1724 3770
rect 1566 3730 1624 3737
rect 1662 3720 1676 3754
rect 1710 3720 1724 3754
rect 1760 3743 1772 3777
rect 1806 3743 2101 3777
rect 1760 3735 2101 3743
rect 2153 3735 2168 3787
rect 11054 3774 11160 3780
rect 1760 3732 2168 3735
rect 1842 3730 2168 3732
rect 4522 3767 4580 3772
rect 4714 3769 5000 3774
rect 4522 3761 4582 3767
rect 1662 3472 1724 3720
rect 4522 3727 4536 3761
rect 4570 3727 4582 3761
rect 4714 3761 4933 3769
rect 4522 3721 4582 3727
rect 4618 3738 4680 3754
rect 4522 3714 4580 3721
rect 4618 3704 4632 3738
rect 4666 3704 4680 3738
rect 4714 3727 4728 3761
rect 4762 3727 4933 3761
rect 4714 3717 4933 3727
rect 4985 3717 5000 3769
rect 4714 3712 5000 3717
rect 5598 3761 7614 3774
rect 5598 3727 7566 3761
rect 7600 3727 7614 3761
rect 7744 3761 8364 3774
rect 5598 3712 7614 3727
rect 7648 3738 7710 3754
rect 4618 3662 4680 3704
rect 4592 3568 4602 3662
rect 4696 3568 4706 3662
rect 1632 3358 1642 3472
rect 1744 3358 1754 3472
rect -1126 3290 -1110 3324
rect -1076 3290 -1020 3324
rect -1126 3276 -1020 3290
rect -2244 2544 -1864 2624
rect -1692 3221 -1646 3236
rect -1692 3187 -1686 3221
rect -1652 3187 -1646 3221
rect -1692 3149 -1646 3187
rect -1692 3115 -1686 3149
rect -1652 3115 -1646 3149
rect -1692 3077 -1646 3115
rect -1692 3043 -1686 3077
rect -1652 3043 -1646 3077
rect -1692 3005 -1646 3043
rect -1692 2971 -1686 3005
rect -1652 2971 -1646 3005
rect -1692 2933 -1646 2971
rect -1692 2899 -1686 2933
rect -1652 2899 -1646 2933
rect -1692 2861 -1646 2899
rect -1692 2827 -1686 2861
rect -1652 2827 -1646 2861
rect -1692 2789 -1646 2827
rect -1692 2755 -1686 2789
rect -1652 2755 -1646 2789
rect -1692 2717 -1646 2755
rect -1692 2683 -1686 2717
rect -1652 2683 -1646 2717
rect -1692 2645 -1646 2683
rect -1692 2611 -1686 2645
rect -1652 2611 -1646 2645
rect -1692 2573 -1646 2611
rect -2244 2506 -2234 2544
rect -1692 2539 -1686 2573
rect -1652 2539 -1646 2573
rect -4724 2461 -4718 2495
rect -4684 2461 -4678 2495
rect -4724 2423 -4678 2461
rect -4724 2389 -4718 2423
rect -4684 2389 -4678 2423
rect -4724 2351 -4678 2389
rect -4724 2317 -4718 2351
rect -4684 2317 -4678 2351
rect -4724 2279 -4678 2317
rect -4724 2245 -4718 2279
rect -4684 2245 -4678 2279
rect -4724 2207 -4678 2245
rect -1692 2501 -1646 2539
rect -1692 2467 -1686 2501
rect -1652 2467 -1646 2501
rect -1692 2429 -1646 2467
rect -1692 2395 -1686 2429
rect -1652 2395 -1646 2429
rect -1692 2357 -1646 2395
rect -1692 2323 -1686 2357
rect -1652 2323 -1646 2357
rect -1692 2285 -1646 2323
rect -1692 2251 -1686 2285
rect -1652 2251 -1646 2285
rect -1692 2236 -1646 2251
rect -1596 3221 -1550 3236
rect -1596 3187 -1590 3221
rect -1556 3187 -1550 3221
rect -1596 3149 -1550 3187
rect -1596 3115 -1590 3149
rect -1556 3115 -1550 3149
rect -1596 3077 -1550 3115
rect -1596 3043 -1590 3077
rect -1556 3043 -1550 3077
rect -1596 3005 -1550 3043
rect -1596 2971 -1590 3005
rect -1556 2971 -1550 3005
rect -1596 2933 -1550 2971
rect -1596 2899 -1590 2933
rect -1556 2899 -1550 2933
rect -1596 2861 -1550 2899
rect -1596 2827 -1590 2861
rect -1556 2827 -1550 2861
rect -1596 2789 -1550 2827
rect -1596 2755 -1590 2789
rect -1556 2755 -1550 2789
rect -1596 2717 -1550 2755
rect -1596 2683 -1590 2717
rect -1556 2683 -1550 2717
rect -1596 2645 -1550 2683
rect -1596 2611 -1590 2645
rect -1556 2611 -1550 2645
rect -1596 2573 -1550 2611
rect -1596 2539 -1590 2573
rect -1556 2539 -1550 2573
rect -1596 2501 -1550 2539
rect -1596 2467 -1590 2501
rect -1556 2467 -1550 2501
rect -1596 2429 -1550 2467
rect -1596 2395 -1590 2429
rect -1556 2395 -1550 2429
rect -1596 2357 -1550 2395
rect -1596 2323 -1590 2357
rect -1556 2323 -1550 2357
rect -1596 2285 -1550 2323
rect -1596 2251 -1590 2285
rect -1556 2251 -1550 2285
rect -1596 2236 -1550 2251
rect -1500 3221 -1454 3236
rect -1500 3187 -1494 3221
rect -1460 3187 -1454 3221
rect -1500 3149 -1454 3187
rect -1500 3115 -1494 3149
rect -1460 3115 -1454 3149
rect -1500 3077 -1454 3115
rect -1500 3043 -1494 3077
rect -1460 3043 -1454 3077
rect -1500 3005 -1454 3043
rect -1500 2971 -1494 3005
rect -1460 2971 -1454 3005
rect -1500 2933 -1454 2971
rect -1500 2899 -1494 2933
rect -1460 2899 -1454 2933
rect -1500 2861 -1454 2899
rect -1500 2827 -1494 2861
rect -1460 2827 -1454 2861
rect -1500 2789 -1454 2827
rect -1500 2755 -1494 2789
rect -1460 2755 -1454 2789
rect -1500 2717 -1454 2755
rect -1500 2683 -1494 2717
rect -1460 2683 -1454 2717
rect -1500 2645 -1454 2683
rect -1500 2611 -1494 2645
rect -1460 2611 -1454 2645
rect -1500 2573 -1454 2611
rect -1500 2539 -1494 2573
rect -1460 2539 -1454 2573
rect -1500 2501 -1454 2539
rect -1500 2467 -1494 2501
rect -1460 2467 -1454 2501
rect -1500 2429 -1454 2467
rect -1500 2395 -1494 2429
rect -1460 2395 -1454 2429
rect -1500 2357 -1454 2395
rect -1500 2323 -1494 2357
rect -1460 2323 -1454 2357
rect -1500 2285 -1454 2323
rect -1500 2251 -1494 2285
rect -1460 2251 -1454 2285
rect -1500 2236 -1454 2251
rect -1404 3221 -1358 3236
rect -1404 3187 -1398 3221
rect -1364 3187 -1358 3221
rect -1404 3149 -1358 3187
rect -1404 3115 -1398 3149
rect -1364 3115 -1358 3149
rect -1404 3077 -1358 3115
rect -1404 3043 -1398 3077
rect -1364 3043 -1358 3077
rect -1404 3005 -1358 3043
rect -1404 2971 -1398 3005
rect -1364 2971 -1358 3005
rect -1404 2933 -1358 2971
rect -1404 2899 -1398 2933
rect -1364 2899 -1358 2933
rect -1404 2861 -1358 2899
rect -1404 2827 -1398 2861
rect -1364 2827 -1358 2861
rect -1404 2789 -1358 2827
rect -1404 2755 -1398 2789
rect -1364 2755 -1358 2789
rect -1404 2717 -1358 2755
rect -1404 2683 -1398 2717
rect -1364 2683 -1358 2717
rect -1404 2645 -1358 2683
rect -1404 2611 -1398 2645
rect -1364 2611 -1358 2645
rect -1404 2573 -1358 2611
rect -1404 2539 -1398 2573
rect -1364 2539 -1358 2573
rect -1404 2501 -1358 2539
rect -1404 2467 -1398 2501
rect -1364 2467 -1358 2501
rect -1404 2429 -1358 2467
rect -1404 2395 -1398 2429
rect -1364 2395 -1358 2429
rect -1404 2357 -1358 2395
rect -1404 2323 -1398 2357
rect -1364 2323 -1358 2357
rect -1404 2285 -1358 2323
rect -1404 2251 -1398 2285
rect -1364 2251 -1358 2285
rect -1404 2236 -1358 2251
rect -1308 3221 -1262 3236
rect -1308 3187 -1302 3221
rect -1268 3187 -1262 3221
rect -1308 3149 -1262 3187
rect -1308 3115 -1302 3149
rect -1268 3115 -1262 3149
rect -1308 3077 -1262 3115
rect -1308 3043 -1302 3077
rect -1268 3043 -1262 3077
rect -1308 3005 -1262 3043
rect -1308 2971 -1302 3005
rect -1268 2971 -1262 3005
rect -1308 2933 -1262 2971
rect -1308 2899 -1302 2933
rect -1268 2899 -1262 2933
rect -1308 2861 -1262 2899
rect -1308 2827 -1302 2861
rect -1268 2827 -1262 2861
rect -1308 2789 -1262 2827
rect -1308 2755 -1302 2789
rect -1268 2755 -1262 2789
rect -1308 2717 -1262 2755
rect -1308 2683 -1302 2717
rect -1268 2683 -1262 2717
rect -1308 2645 -1262 2683
rect -1308 2611 -1302 2645
rect -1268 2611 -1262 2645
rect -1308 2573 -1262 2611
rect -1308 2539 -1302 2573
rect -1268 2539 -1262 2573
rect -1308 2501 -1262 2539
rect -1308 2467 -1302 2501
rect -1268 2467 -1262 2501
rect -1308 2429 -1262 2467
rect -1308 2395 -1302 2429
rect -1268 2395 -1262 2429
rect -1308 2357 -1262 2395
rect -1308 2323 -1302 2357
rect -1268 2323 -1262 2357
rect -1308 2285 -1262 2323
rect -1308 2251 -1302 2285
rect -1268 2251 -1262 2285
rect -1308 2236 -1262 2251
rect -1212 3221 -1166 3236
rect -1212 3187 -1206 3221
rect -1172 3187 -1166 3221
rect -1212 3149 -1166 3187
rect -1212 3115 -1206 3149
rect -1172 3115 -1166 3149
rect -1212 3077 -1166 3115
rect -1212 3043 -1206 3077
rect -1172 3043 -1166 3077
rect -1212 3005 -1166 3043
rect -1212 2971 -1206 3005
rect -1172 2971 -1166 3005
rect -1212 2933 -1166 2971
rect -1212 2899 -1206 2933
rect -1172 2899 -1166 2933
rect -1212 2861 -1166 2899
rect -1212 2827 -1206 2861
rect -1172 2827 -1166 2861
rect -1212 2789 -1166 2827
rect -1212 2755 -1206 2789
rect -1172 2755 -1166 2789
rect -1212 2717 -1166 2755
rect -1212 2683 -1206 2717
rect -1172 2683 -1166 2717
rect -1212 2645 -1166 2683
rect -1212 2611 -1206 2645
rect -1172 2611 -1166 2645
rect -1212 2573 -1166 2611
rect -1212 2539 -1206 2573
rect -1172 2539 -1166 2573
rect -1212 2501 -1166 2539
rect -1212 2467 -1206 2501
rect -1172 2467 -1166 2501
rect -1212 2429 -1166 2467
rect -1212 2395 -1206 2429
rect -1172 2395 -1166 2429
rect -1212 2357 -1166 2395
rect -1212 2323 -1206 2357
rect -1172 2323 -1166 2357
rect -1212 2285 -1166 2323
rect -1212 2251 -1206 2285
rect -1172 2251 -1166 2285
rect -1212 2236 -1166 2251
rect -1116 3221 -1070 3236
rect -1116 3187 -1110 3221
rect -1076 3187 -1070 3221
rect -1116 3149 -1070 3187
rect -1116 3115 -1110 3149
rect -1076 3115 -1070 3149
rect -1116 3077 -1070 3115
rect -1116 3043 -1110 3077
rect -1076 3043 -1070 3077
rect -1116 3005 -1070 3043
rect -1116 2971 -1110 3005
rect -1076 2971 -1070 3005
rect -1116 2933 -1070 2971
rect -1116 2899 -1110 2933
rect -1076 2899 -1070 2933
rect -1116 2861 -1070 2899
rect -1116 2827 -1110 2861
rect -1076 2827 -1070 2861
rect -1116 2789 -1070 2827
rect -1116 2755 -1110 2789
rect -1076 2755 -1070 2789
rect -1116 2717 -1070 2755
rect -1116 2683 -1110 2717
rect -1076 2683 -1070 2717
rect -1116 2645 -1070 2683
rect -1116 2611 -1110 2645
rect -1076 2611 -1070 2645
rect -1116 2573 -1070 2611
rect -1116 2539 -1110 2573
rect -1076 2539 -1070 2573
rect -1116 2501 -1070 2539
rect -1116 2467 -1110 2501
rect -1076 2467 -1070 2501
rect -1116 2429 -1070 2467
rect -1116 2395 -1110 2429
rect -1076 2395 -1070 2429
rect -1116 2357 -1070 2395
rect -1116 2323 -1110 2357
rect -1076 2323 -1070 2357
rect -1116 2285 -1070 2323
rect -1116 2251 -1110 2285
rect -1076 2251 -1070 2285
rect -1116 2236 -1070 2251
rect -1020 3221 -974 3236
rect -1020 3187 -1014 3221
rect -980 3187 -974 3221
rect -1020 3149 -974 3187
rect -1020 3115 -1014 3149
rect -980 3115 -974 3149
rect -1020 3077 -974 3115
rect -1020 3043 -1014 3077
rect -980 3043 -974 3077
rect -1020 3005 -974 3043
rect -1020 2971 -1014 3005
rect -980 2971 -974 3005
rect -1020 2933 -974 2971
rect -1020 2899 -1014 2933
rect -980 2899 -974 2933
rect -1020 2861 -974 2899
rect -1020 2827 -1014 2861
rect -980 2827 -974 2861
rect -1020 2789 -974 2827
rect -1020 2755 -1014 2789
rect -980 2755 -974 2789
rect -1020 2717 -974 2755
rect -1020 2683 -1014 2717
rect -980 2683 -974 2717
rect -1020 2645 -974 2683
rect -1020 2611 -1014 2645
rect -980 2611 -974 2645
rect -1020 2573 -974 2611
rect -1020 2539 -1014 2573
rect -980 2539 -974 2573
rect -1020 2501 -974 2539
rect -1020 2467 -1014 2501
rect -980 2467 -974 2501
rect -1020 2429 -974 2467
rect -1020 2395 -1014 2429
rect -980 2395 -974 2429
rect -1020 2357 -974 2395
rect -1020 2323 -1014 2357
rect -980 2323 -974 2357
rect -1020 2285 -974 2323
rect -1020 2251 -1014 2285
rect -980 2251 -974 2285
rect -1020 2236 -974 2251
rect -924 3221 -878 3236
rect -924 3187 -918 3221
rect -884 3187 -878 3221
rect -924 3149 -878 3187
rect -924 3115 -918 3149
rect -884 3115 -878 3149
rect -924 3077 -878 3115
rect -924 3043 -918 3077
rect -884 3043 -878 3077
rect -924 3005 -878 3043
rect 1662 3086 1724 3358
rect 3658 3305 3720 3320
rect 3658 3253 3663 3305
rect 3715 3253 3720 3305
rect 3658 3086 3720 3253
rect 1662 3024 4244 3086
rect -924 2971 -918 3005
rect -884 2971 -878 3005
rect -924 2933 -878 2971
rect 1394 3013 1626 3018
rect 1394 2961 1409 3013
rect 1461 3002 1626 3013
rect 1461 2968 1578 3002
rect 1612 2968 1626 3002
rect 1461 2961 1626 2968
rect 1394 2956 1626 2961
rect 1662 2994 1724 3024
rect 1662 2960 1674 2994
rect 1708 2960 1724 2994
rect 1662 2948 1724 2960
rect -924 2899 -918 2933
rect -884 2899 -878 2933
rect -924 2861 -878 2899
rect -924 2827 -918 2861
rect -884 2827 -878 2861
rect -924 2789 -878 2827
rect -924 2755 -918 2789
rect -884 2755 -878 2789
rect -924 2717 -878 2755
rect -924 2683 -918 2717
rect -884 2683 -878 2717
rect -924 2645 -878 2683
rect -924 2611 -918 2645
rect -884 2611 -878 2645
rect -924 2573 -878 2611
rect -924 2539 -918 2573
rect -884 2539 -878 2573
rect -924 2501 -878 2539
rect -924 2467 -918 2501
rect -884 2467 -878 2501
rect -924 2429 -878 2467
rect -924 2395 -918 2429
rect -884 2395 -878 2429
rect -924 2357 -878 2395
rect -924 2323 -918 2357
rect -884 2323 -878 2357
rect -924 2285 -878 2323
rect -924 2251 -918 2285
rect -884 2251 -878 2285
rect -924 2236 -878 2251
rect 1476 2815 1522 2830
rect 1476 2781 1482 2815
rect 1516 2781 1522 2815
rect 1476 2743 1522 2781
rect 1476 2709 1482 2743
rect 1516 2709 1522 2743
rect 1476 2671 1522 2709
rect 1476 2637 1482 2671
rect 1516 2637 1522 2671
rect 1476 2599 1522 2637
rect 1476 2565 1482 2599
rect 1516 2565 1522 2599
rect 1476 2527 1522 2565
rect 1476 2493 1482 2527
rect 1516 2493 1522 2527
rect 1476 2455 1522 2493
rect 1476 2421 1482 2455
rect 1516 2421 1522 2455
rect 1476 2383 1522 2421
rect 1476 2349 1482 2383
rect 1516 2349 1522 2383
rect 1476 2311 1522 2349
rect 1476 2277 1482 2311
rect 1516 2277 1522 2311
rect 1476 2239 1522 2277
rect -4724 2173 -4718 2207
rect -4684 2173 -4678 2207
rect 1476 2205 1482 2239
rect 1516 2205 1522 2239
rect -4724 2135 -4678 2173
rect -4724 2101 -4718 2135
rect -4684 2101 -4678 2135
rect -4724 2063 -4678 2101
rect -4724 2029 -4718 2063
rect -4684 2029 -4678 2063
rect -4724 1991 -4678 2029
rect -4724 1957 -4718 1991
rect -4684 1957 -4678 1991
rect -4724 1919 -4678 1957
rect -4724 1885 -4718 1919
rect -4684 1885 -4678 1919
rect -4724 1870 -4678 1885
rect -1110 2172 -1048 2190
rect -1110 2138 -1097 2172
rect -1063 2138 -1048 2172
rect -9442 1675 -9066 1678
rect -9442 1495 -9408 1675
rect -9100 1495 -9066 1675
rect -9442 1492 -9066 1495
rect -7442 1675 -7066 1678
rect -7442 1495 -7408 1675
rect -7100 1495 -7066 1675
rect -7442 1492 -7066 1495
rect -5444 1675 -5066 1678
rect -5444 1495 -5409 1675
rect -5101 1495 -5066 1675
rect -5444 1492 -5066 1495
rect -1110 1298 -1048 2138
rect 1476 2167 1522 2205
rect 1476 2133 1482 2167
rect 1516 2133 1522 2167
rect 1476 2095 1522 2133
rect 1476 2061 1482 2095
rect 1516 2061 1522 2095
rect 1476 2023 1522 2061
rect 1476 1989 1482 2023
rect 1516 1989 1522 2023
rect 1476 1951 1522 1989
rect 1476 1917 1482 1951
rect 1516 1917 1522 1951
rect 1476 1879 1522 1917
rect 1476 1845 1482 1879
rect 1516 1845 1522 1879
rect 1476 1830 1522 1845
rect 1572 2815 1618 2830
rect 1572 2781 1578 2815
rect 1612 2781 1618 2815
rect 1572 2743 1618 2781
rect 1572 2709 1578 2743
rect 1612 2709 1618 2743
rect 1572 2671 1618 2709
rect 1572 2637 1578 2671
rect 1612 2637 1618 2671
rect 1572 2599 1618 2637
rect 1572 2565 1578 2599
rect 1612 2565 1618 2599
rect 1572 2527 1618 2565
rect 1572 2493 1578 2527
rect 1612 2493 1618 2527
rect 1572 2455 1618 2493
rect 1572 2421 1578 2455
rect 1612 2421 1618 2455
rect 1572 2383 1618 2421
rect 1572 2349 1578 2383
rect 1612 2349 1618 2383
rect 1572 2311 1618 2349
rect 1572 2277 1578 2311
rect 1612 2277 1618 2311
rect 1572 2239 1618 2277
rect 1572 2205 1578 2239
rect 1612 2205 1618 2239
rect 1572 2167 1618 2205
rect 1572 2133 1578 2167
rect 1612 2133 1618 2167
rect 1572 2095 1618 2133
rect 1572 2061 1578 2095
rect 1612 2061 1618 2095
rect 1572 2023 1618 2061
rect 1572 1989 1578 2023
rect 1612 1989 1618 2023
rect 1572 1951 1618 1989
rect 1572 1917 1578 1951
rect 1612 1917 1618 1951
rect 1572 1879 1618 1917
rect 1572 1845 1578 1879
rect 1612 1845 1618 1879
rect 1572 1830 1618 1845
rect 1668 2815 1714 2830
rect 1668 2781 1674 2815
rect 1708 2781 1714 2815
rect 1668 2743 1714 2781
rect 1668 2709 1674 2743
rect 1708 2709 1714 2743
rect 1668 2671 1714 2709
rect 1668 2637 1674 2671
rect 1708 2637 1714 2671
rect 1668 2599 1714 2637
rect 1668 2565 1674 2599
rect 1708 2565 1714 2599
rect 1668 2527 1714 2565
rect 1668 2493 1674 2527
rect 1708 2493 1714 2527
rect 1668 2455 1714 2493
rect 1668 2421 1674 2455
rect 1708 2421 1714 2455
rect 1668 2383 1714 2421
rect 1668 2349 1674 2383
rect 1708 2349 1714 2383
rect 1668 2311 1714 2349
rect 1668 2277 1674 2311
rect 1708 2277 1714 2311
rect 1668 2239 1714 2277
rect 1668 2205 1674 2239
rect 1708 2205 1714 2239
rect 1668 2167 1714 2205
rect 1668 2133 1674 2167
rect 1708 2133 1714 2167
rect 1668 2095 1714 2133
rect 1668 2061 1674 2095
rect 1708 2061 1714 2095
rect 1668 2023 1714 2061
rect 1668 1989 1674 2023
rect 1708 1989 1714 2023
rect 1668 1951 1714 1989
rect 1668 1917 1674 1951
rect 1708 1917 1714 1951
rect 1668 1879 1714 1917
rect 1668 1845 1674 1879
rect 1708 1845 1714 1879
rect 1668 1830 1714 1845
rect 1764 2815 1810 2830
rect 1764 2781 1770 2815
rect 1804 2781 1810 2815
rect 1764 2743 1810 2781
rect 1764 2709 1770 2743
rect 1804 2709 1810 2743
rect 1764 2671 1810 2709
rect 1764 2637 1770 2671
rect 1804 2637 1810 2671
rect 1764 2599 1810 2637
rect 1764 2565 1770 2599
rect 1804 2565 1810 2599
rect 1764 2527 1810 2565
rect 1764 2493 1770 2527
rect 1804 2493 1810 2527
rect 1764 2455 1810 2493
rect 1764 2421 1770 2455
rect 1804 2421 1810 2455
rect 1764 2383 1810 2421
rect 1764 2349 1770 2383
rect 1804 2349 1810 2383
rect 1764 2311 1810 2349
rect 1764 2277 1770 2311
rect 1804 2277 1810 2311
rect 1764 2239 1810 2277
rect 1764 2205 1770 2239
rect 1804 2205 1810 2239
rect 1764 2167 1810 2205
rect 1764 2133 1770 2167
rect 1804 2133 1810 2167
rect 1764 2095 1810 2133
rect 1764 2061 1770 2095
rect 1804 2061 1810 2095
rect 1764 2023 1810 2061
rect 1764 1989 1770 2023
rect 1804 1989 1810 2023
rect 1764 1951 1810 1989
rect 1764 1917 1770 1951
rect 1804 1917 1810 1951
rect 1764 1879 1810 1917
rect 1764 1845 1770 1879
rect 1804 1845 1810 1879
rect 1764 1830 1810 1845
rect 1860 2815 1906 2830
rect 1860 2781 1866 2815
rect 1900 2781 1906 2815
rect 1860 2743 1906 2781
rect 1860 2709 1866 2743
rect 1900 2709 1906 2743
rect 1860 2671 1906 2709
rect 1860 2637 1866 2671
rect 1900 2637 1906 2671
rect 1860 2599 1906 2637
rect 1860 2565 1866 2599
rect 1900 2565 1906 2599
rect 1860 2527 1906 2565
rect 1860 2493 1866 2527
rect 1900 2493 1906 2527
rect 1860 2455 1906 2493
rect 1860 2421 1866 2455
rect 1900 2421 1906 2455
rect 1860 2383 1906 2421
rect 1860 2349 1866 2383
rect 1900 2349 1906 2383
rect 1860 2311 1906 2349
rect 1860 2277 1866 2311
rect 1900 2277 1906 2311
rect 2232 2360 2294 3024
rect 4182 3000 4244 3024
rect 4618 3068 4680 3568
rect 5600 3215 5662 3712
rect 7648 3704 7662 3738
rect 7696 3704 7710 3738
rect 7744 3727 7758 3761
rect 7792 3727 8364 3761
rect 7744 3712 8364 3727
rect 10008 3767 10698 3772
rect 10008 3715 10023 3767
rect 10075 3765 10698 3767
rect 10830 3769 11160 3774
rect 10075 3759 10700 3765
rect 10075 3725 10654 3759
rect 10688 3725 10700 3759
rect 10830 3759 11081 3769
rect 10075 3719 10700 3725
rect 10736 3736 10798 3752
rect 10075 3715 10698 3719
rect 7648 3532 7710 3704
rect 7122 3479 7710 3532
rect 7122 3427 7127 3479
rect 7179 3470 7710 3479
rect 7179 3427 7184 3470
rect 7122 3412 7184 3427
rect 5600 3163 5605 3215
rect 5657 3163 5662 3215
rect 5600 3148 5662 3163
rect 7284 3158 7346 3170
rect 7276 3151 7384 3158
rect 7276 3099 7304 3151
rect 7356 3099 7384 3151
rect 7276 3092 7384 3099
rect 4618 3006 7200 3068
rect 4182 2992 4560 3000
rect 4182 2986 4580 2992
rect 4182 2952 4534 2986
rect 4568 2952 4580 2986
rect 4182 2946 4580 2952
rect 4618 2978 4680 3006
rect 4182 2938 4560 2946
rect 4618 2944 4630 2978
rect 4664 2944 4680 2978
rect 4618 2932 4680 2944
rect 4432 2799 4478 2814
rect 4432 2765 4438 2799
rect 4472 2765 4478 2799
rect 4432 2727 4478 2765
rect 4432 2693 4438 2727
rect 4472 2693 4478 2727
rect 4432 2655 4478 2693
rect 2550 2592 2642 2622
rect 2550 2540 2570 2592
rect 2622 2540 2642 2592
rect 2550 2428 2642 2540
rect 2550 2394 2579 2428
rect 2613 2394 2642 2428
rect 2550 2388 2642 2394
rect 4432 2621 4438 2655
rect 4472 2621 4478 2655
rect 4432 2583 4478 2621
rect 4432 2549 4438 2583
rect 4472 2549 4478 2583
rect 4432 2511 4478 2549
rect 4432 2477 4438 2511
rect 4472 2477 4478 2511
rect 4432 2439 4478 2477
rect 4432 2405 4438 2439
rect 4472 2405 4478 2439
rect 4432 2367 4478 2405
rect 2232 2350 2438 2360
rect 2232 2316 2392 2350
rect 2426 2316 2438 2350
rect 2232 2298 2438 2316
rect 4432 2333 4438 2367
rect 4472 2333 4478 2367
rect 1860 2239 1906 2277
rect 4432 2295 4478 2333
rect 1860 2205 1866 2239
rect 1900 2205 1906 2239
rect 1860 2167 1906 2205
rect 1860 2133 1866 2167
rect 1900 2133 1906 2167
rect 1860 2095 1906 2133
rect 1860 2061 1866 2095
rect 1900 2061 1906 2095
rect 2494 2229 2540 2276
rect 2494 2195 2500 2229
rect 2534 2195 2540 2229
rect 2494 2157 2540 2195
rect 2494 2123 2500 2157
rect 2534 2123 2540 2157
rect 2494 2076 2540 2123
rect 2652 2229 2698 2276
rect 2652 2195 2658 2229
rect 2692 2195 2698 2229
rect 2652 2157 2698 2195
rect 2652 2123 2658 2157
rect 2692 2123 2698 2157
rect 2652 2076 2698 2123
rect 4432 2261 4438 2295
rect 4472 2261 4478 2295
rect 4432 2223 4478 2261
rect 4432 2189 4438 2223
rect 4472 2189 4478 2223
rect 4432 2151 4478 2189
rect 4432 2117 4438 2151
rect 4472 2117 4478 2151
rect 4432 2079 4478 2117
rect 1860 2023 1906 2061
rect 1860 1989 1866 2023
rect 1900 1989 1906 2023
rect 1860 1951 1906 1989
rect 1860 1917 1866 1951
rect 1900 1917 1906 1951
rect 1860 1879 1906 1917
rect 1860 1845 1866 1879
rect 1900 1845 1906 1879
rect 1860 1830 1906 1845
rect 4432 2045 4438 2079
rect 4472 2045 4478 2079
rect 4432 2007 4478 2045
rect 4432 1973 4438 2007
rect 4472 1973 4478 2007
rect 4432 1935 4478 1973
rect 4432 1901 4438 1935
rect 4472 1901 4478 1935
rect 4432 1863 4478 1901
rect 4432 1829 4438 1863
rect 4472 1829 4478 1863
rect 4432 1814 4478 1829
rect 4528 2799 4574 2814
rect 4528 2765 4534 2799
rect 4568 2765 4574 2799
rect 4528 2727 4574 2765
rect 4528 2693 4534 2727
rect 4568 2693 4574 2727
rect 4528 2655 4574 2693
rect 4528 2621 4534 2655
rect 4568 2621 4574 2655
rect 4528 2583 4574 2621
rect 4528 2549 4534 2583
rect 4568 2549 4574 2583
rect 4528 2511 4574 2549
rect 4528 2477 4534 2511
rect 4568 2477 4574 2511
rect 4528 2439 4574 2477
rect 4528 2405 4534 2439
rect 4568 2405 4574 2439
rect 4528 2367 4574 2405
rect 4528 2333 4534 2367
rect 4568 2333 4574 2367
rect 4528 2295 4574 2333
rect 4528 2261 4534 2295
rect 4568 2261 4574 2295
rect 4528 2223 4574 2261
rect 4528 2189 4534 2223
rect 4568 2189 4574 2223
rect 4528 2151 4574 2189
rect 4528 2117 4534 2151
rect 4568 2117 4574 2151
rect 4528 2079 4574 2117
rect 4528 2045 4534 2079
rect 4568 2045 4574 2079
rect 4528 2007 4574 2045
rect 4528 1973 4534 2007
rect 4568 1973 4574 2007
rect 4528 1935 4574 1973
rect 4528 1901 4534 1935
rect 4568 1901 4574 1935
rect 4528 1863 4574 1901
rect 4528 1829 4534 1863
rect 4568 1829 4574 1863
rect 4528 1814 4574 1829
rect 4624 2799 4670 2814
rect 4624 2765 4630 2799
rect 4664 2765 4670 2799
rect 4624 2727 4670 2765
rect 4624 2693 4630 2727
rect 4664 2693 4670 2727
rect 4624 2655 4670 2693
rect 4624 2621 4630 2655
rect 4664 2621 4670 2655
rect 4624 2583 4670 2621
rect 4624 2549 4630 2583
rect 4664 2549 4670 2583
rect 4624 2511 4670 2549
rect 4624 2477 4630 2511
rect 4664 2477 4670 2511
rect 4624 2439 4670 2477
rect 4624 2405 4630 2439
rect 4664 2405 4670 2439
rect 4624 2367 4670 2405
rect 4624 2333 4630 2367
rect 4664 2333 4670 2367
rect 4624 2295 4670 2333
rect 4624 2261 4630 2295
rect 4664 2261 4670 2295
rect 4624 2223 4670 2261
rect 4624 2189 4630 2223
rect 4664 2189 4670 2223
rect 4624 2151 4670 2189
rect 4624 2117 4630 2151
rect 4664 2117 4670 2151
rect 4624 2079 4670 2117
rect 4624 2045 4630 2079
rect 4664 2045 4670 2079
rect 4624 2007 4670 2045
rect 4624 1973 4630 2007
rect 4664 1973 4670 2007
rect 4624 1935 4670 1973
rect 4624 1901 4630 1935
rect 4664 1901 4670 1935
rect 4624 1863 4670 1901
rect 4624 1829 4630 1863
rect 4664 1829 4670 1863
rect 4624 1814 4670 1829
rect 4720 2799 4766 2814
rect 4720 2765 4726 2799
rect 4760 2765 4766 2799
rect 4720 2727 4766 2765
rect 4720 2693 4726 2727
rect 4760 2693 4766 2727
rect 4720 2655 4766 2693
rect 4720 2621 4726 2655
rect 4760 2621 4766 2655
rect 4720 2583 4766 2621
rect 4720 2549 4726 2583
rect 4760 2549 4766 2583
rect 4720 2511 4766 2549
rect 4720 2477 4726 2511
rect 4760 2477 4766 2511
rect 4720 2439 4766 2477
rect 4720 2405 4726 2439
rect 4760 2405 4766 2439
rect 4720 2367 4766 2405
rect 4720 2333 4726 2367
rect 4760 2333 4766 2367
rect 4720 2295 4766 2333
rect 4720 2261 4726 2295
rect 4760 2261 4766 2295
rect 4720 2223 4766 2261
rect 4720 2189 4726 2223
rect 4760 2189 4766 2223
rect 4720 2151 4766 2189
rect 4720 2117 4726 2151
rect 4760 2117 4766 2151
rect 4720 2079 4766 2117
rect 4720 2045 4726 2079
rect 4760 2045 4766 2079
rect 4720 2007 4766 2045
rect 4720 1973 4726 2007
rect 4760 1973 4766 2007
rect 4720 1935 4766 1973
rect 4720 1901 4726 1935
rect 4760 1901 4766 1935
rect 4720 1863 4766 1901
rect 4720 1829 4726 1863
rect 4760 1829 4766 1863
rect 4720 1814 4766 1829
rect 4816 2799 4862 2814
rect 4816 2765 4822 2799
rect 4856 2765 4862 2799
rect 4816 2727 4862 2765
rect 4816 2693 4822 2727
rect 4856 2693 4862 2727
rect 4816 2655 4862 2693
rect 4816 2621 4822 2655
rect 4856 2621 4862 2655
rect 4816 2583 4862 2621
rect 4816 2549 4822 2583
rect 4856 2549 4862 2583
rect 4816 2511 4862 2549
rect 4816 2477 4822 2511
rect 4856 2477 4862 2511
rect 4816 2439 4862 2477
rect 4816 2405 4822 2439
rect 4856 2405 4862 2439
rect 4816 2367 4862 2405
rect 4816 2333 4822 2367
rect 4856 2333 4862 2367
rect 4816 2295 4862 2333
rect 5132 2360 5194 3006
rect 7138 3000 7200 3006
rect 7284 3000 7346 3092
rect 7648 3048 7710 3470
rect 8298 3408 8360 3712
rect 10008 3710 10698 3715
rect 10736 3702 10750 3736
rect 10784 3702 10798 3736
rect 10830 3725 10846 3759
rect 10880 3725 11081 3759
rect 10830 3717 11081 3725
rect 11133 3717 11160 3769
rect 15332 3779 15614 3794
rect 10830 3710 11160 3717
rect 11054 3706 11160 3710
rect 13560 3739 13854 3748
rect 13560 3733 13856 3739
rect 8672 3660 8762 3676
rect 8672 3608 8691 3660
rect 8743 3652 8762 3660
rect 10736 3652 10798 3702
rect 8743 3608 10798 3652
rect 8672 3596 10798 3608
rect 8672 3592 8762 3596
rect 10404 3471 10466 3486
rect 10404 3419 10409 3471
rect 10461 3419 10466 3471
rect 10404 3408 10466 3419
rect 8298 3406 10466 3408
rect 8298 3354 8772 3406
rect 8824 3354 10466 3406
rect 8298 3350 10466 3354
rect 8298 3346 10464 3350
rect 7138 2992 7608 3000
rect 7648 2998 10260 3048
rect 10736 3046 10798 3596
rect 13560 3699 13810 3733
rect 13844 3699 13856 3733
rect 13988 3733 14642 3750
rect 13560 3693 13856 3699
rect 13892 3710 13954 3726
rect 13560 3684 13854 3693
rect 13076 3471 13138 3486
rect 13560 3474 13628 3684
rect 13892 3676 13906 3710
rect 13940 3676 13954 3710
rect 13988 3699 14002 3733
rect 14036 3699 14642 3733
rect 13988 3684 14642 3699
rect 13892 3490 13954 3676
rect 13076 3419 13081 3471
rect 13133 3419 13138 3471
rect 13076 3300 13138 3419
rect 13426 3464 13628 3474
rect 13426 3412 13441 3464
rect 13493 3412 13628 3464
rect 13882 3481 13972 3490
rect 13882 3429 13901 3481
rect 13953 3429 13972 3481
rect 13882 3420 13972 3429
rect 13426 3410 13628 3412
rect 13892 3300 13954 3420
rect 13076 3238 13954 3300
rect 13892 3174 13954 3238
rect 13892 3112 14296 3174
rect 7138 2986 7610 2992
rect 7138 2952 7564 2986
rect 7598 2952 7610 2986
rect 7138 2946 7610 2952
rect 7648 2986 10698 2998
rect 7648 2978 7710 2986
rect 7138 2938 7608 2946
rect 7648 2944 7660 2978
rect 7694 2944 7710 2978
rect 7648 2932 7710 2944
rect 7462 2799 7508 2814
rect 7462 2765 7468 2799
rect 7502 2765 7508 2799
rect 7462 2727 7508 2765
rect 7462 2693 7468 2727
rect 7502 2693 7508 2727
rect 7462 2655 7508 2693
rect 5550 2592 5642 2622
rect 5550 2540 5570 2592
rect 5622 2540 5642 2592
rect 5550 2428 5642 2540
rect 5550 2394 5579 2428
rect 5613 2394 5642 2428
rect 5550 2388 5642 2394
rect 7462 2621 7468 2655
rect 7502 2621 7508 2655
rect 7462 2583 7508 2621
rect 7462 2549 7468 2583
rect 7502 2549 7508 2583
rect 7462 2511 7508 2549
rect 7462 2477 7468 2511
rect 7502 2477 7508 2511
rect 7462 2439 7508 2477
rect 7462 2405 7468 2439
rect 7502 2405 7508 2439
rect 7462 2367 7508 2405
rect 5132 2350 5438 2360
rect 5132 2316 5392 2350
rect 5426 2316 5438 2350
rect 5132 2298 5438 2316
rect 7462 2333 7468 2367
rect 7502 2333 7508 2367
rect 4816 2261 4822 2295
rect 4856 2261 4862 2295
rect 7462 2295 7508 2333
rect 4816 2223 4862 2261
rect 4816 2189 4822 2223
rect 4856 2189 4862 2223
rect 4816 2151 4862 2189
rect 4816 2117 4822 2151
rect 4856 2117 4862 2151
rect 4816 2079 4862 2117
rect 4816 2045 4822 2079
rect 4856 2045 4862 2079
rect 5494 2229 5540 2276
rect 5494 2195 5500 2229
rect 5534 2195 5540 2229
rect 5494 2157 5540 2195
rect 5494 2123 5500 2157
rect 5534 2123 5540 2157
rect 5494 2076 5540 2123
rect 5652 2229 5698 2276
rect 5652 2195 5658 2229
rect 5692 2195 5698 2229
rect 5652 2157 5698 2195
rect 5652 2123 5658 2157
rect 5692 2123 5698 2157
rect 5652 2076 5698 2123
rect 7462 2261 7468 2295
rect 7502 2261 7508 2295
rect 7462 2223 7508 2261
rect 7462 2189 7468 2223
rect 7502 2189 7508 2223
rect 7462 2151 7508 2189
rect 7462 2117 7468 2151
rect 7502 2117 7508 2151
rect 7462 2079 7508 2117
rect 4816 2007 4862 2045
rect 4816 1973 4822 2007
rect 4856 1973 4862 2007
rect 4816 1935 4862 1973
rect 4816 1901 4822 1935
rect 4856 1901 4862 1935
rect 4816 1863 4862 1901
rect 4816 1829 4822 1863
rect 4856 1829 4862 1863
rect 4816 1814 4862 1829
rect 7462 2045 7468 2079
rect 7502 2045 7508 2079
rect 7462 2007 7508 2045
rect 7462 1973 7468 2007
rect 7502 1973 7508 2007
rect 7462 1935 7508 1973
rect 7462 1901 7468 1935
rect 7502 1901 7508 1935
rect 7462 1863 7508 1901
rect 7462 1829 7468 1863
rect 7502 1829 7508 1863
rect 7462 1814 7508 1829
rect 7558 2799 7604 2814
rect 7558 2765 7564 2799
rect 7598 2765 7604 2799
rect 7558 2727 7604 2765
rect 7558 2693 7564 2727
rect 7598 2693 7604 2727
rect 7558 2655 7604 2693
rect 7558 2621 7564 2655
rect 7598 2621 7604 2655
rect 7558 2583 7604 2621
rect 7558 2549 7564 2583
rect 7598 2549 7604 2583
rect 7558 2511 7604 2549
rect 7558 2477 7564 2511
rect 7598 2477 7604 2511
rect 7558 2439 7604 2477
rect 7558 2405 7564 2439
rect 7598 2405 7604 2439
rect 7558 2367 7604 2405
rect 7558 2333 7564 2367
rect 7598 2333 7604 2367
rect 7558 2295 7604 2333
rect 7558 2261 7564 2295
rect 7598 2261 7604 2295
rect 7558 2223 7604 2261
rect 7558 2189 7564 2223
rect 7598 2189 7604 2223
rect 7558 2151 7604 2189
rect 7558 2117 7564 2151
rect 7598 2117 7604 2151
rect 7558 2079 7604 2117
rect 7558 2045 7564 2079
rect 7598 2045 7604 2079
rect 7558 2007 7604 2045
rect 7558 1973 7564 2007
rect 7598 1973 7604 2007
rect 7558 1935 7604 1973
rect 7558 1901 7564 1935
rect 7598 1901 7604 1935
rect 7558 1863 7604 1901
rect 7558 1829 7564 1863
rect 7598 1829 7604 1863
rect 7558 1814 7604 1829
rect 7654 2799 7700 2814
rect 7654 2765 7660 2799
rect 7694 2765 7700 2799
rect 7654 2727 7700 2765
rect 7654 2693 7660 2727
rect 7694 2693 7700 2727
rect 7654 2655 7700 2693
rect 7654 2621 7660 2655
rect 7694 2621 7700 2655
rect 7654 2583 7700 2621
rect 7654 2549 7660 2583
rect 7694 2549 7700 2583
rect 7654 2511 7700 2549
rect 7654 2477 7660 2511
rect 7694 2477 7700 2511
rect 7654 2439 7700 2477
rect 7654 2405 7660 2439
rect 7694 2405 7700 2439
rect 7654 2367 7700 2405
rect 7654 2333 7660 2367
rect 7694 2333 7700 2367
rect 7654 2295 7700 2333
rect 7654 2261 7660 2295
rect 7694 2261 7700 2295
rect 7654 2223 7700 2261
rect 7654 2189 7660 2223
rect 7694 2189 7700 2223
rect 7654 2151 7700 2189
rect 7654 2117 7660 2151
rect 7694 2117 7700 2151
rect 7654 2079 7700 2117
rect 7654 2045 7660 2079
rect 7694 2045 7700 2079
rect 7654 2007 7700 2045
rect 7654 1973 7660 2007
rect 7694 1973 7700 2007
rect 7654 1935 7700 1973
rect 7654 1901 7660 1935
rect 7694 1901 7700 1935
rect 7654 1863 7700 1901
rect 7654 1829 7660 1863
rect 7694 1829 7700 1863
rect 7654 1814 7700 1829
rect 7750 2799 7796 2814
rect 7750 2765 7756 2799
rect 7790 2765 7796 2799
rect 7750 2727 7796 2765
rect 7750 2693 7756 2727
rect 7790 2693 7796 2727
rect 7750 2655 7796 2693
rect 7750 2621 7756 2655
rect 7790 2621 7796 2655
rect 7750 2583 7796 2621
rect 7750 2549 7756 2583
rect 7790 2549 7796 2583
rect 7750 2511 7796 2549
rect 7750 2477 7756 2511
rect 7790 2477 7796 2511
rect 7750 2439 7796 2477
rect 7750 2405 7756 2439
rect 7790 2405 7796 2439
rect 7750 2367 7796 2405
rect 7750 2333 7756 2367
rect 7790 2333 7796 2367
rect 7750 2295 7796 2333
rect 7750 2261 7756 2295
rect 7790 2261 7796 2295
rect 7750 2223 7796 2261
rect 7750 2189 7756 2223
rect 7790 2189 7796 2223
rect 7750 2151 7796 2189
rect 7750 2117 7756 2151
rect 7790 2117 7796 2151
rect 7750 2079 7796 2117
rect 7750 2045 7756 2079
rect 7790 2045 7796 2079
rect 7750 2007 7796 2045
rect 7750 1973 7756 2007
rect 7790 1973 7796 2007
rect 7750 1935 7796 1973
rect 7750 1901 7756 1935
rect 7790 1901 7796 1935
rect 7750 1863 7796 1901
rect 7750 1829 7756 1863
rect 7790 1829 7796 1863
rect 7750 1814 7796 1829
rect 7846 2799 7892 2814
rect 7846 2765 7852 2799
rect 7886 2765 7892 2799
rect 7846 2727 7892 2765
rect 7846 2693 7852 2727
rect 7886 2693 7892 2727
rect 7846 2655 7892 2693
rect 7846 2621 7852 2655
rect 7886 2621 7892 2655
rect 7846 2583 7892 2621
rect 7846 2549 7852 2583
rect 7886 2549 7892 2583
rect 7846 2511 7892 2549
rect 7846 2477 7852 2511
rect 7886 2477 7892 2511
rect 7846 2439 7892 2477
rect 7846 2405 7852 2439
rect 7886 2405 7892 2439
rect 7846 2367 7892 2405
rect 7846 2333 7852 2367
rect 7886 2333 7892 2367
rect 7846 2295 7892 2333
rect 8232 2360 8294 2986
rect 10196 2984 10698 2986
rect 10196 2950 10652 2984
rect 10686 2950 10698 2984
rect 10196 2936 10698 2950
rect 10736 2984 13522 3046
rect 10736 2976 10798 2984
rect 10736 2942 10748 2976
rect 10782 2942 10798 2976
rect 10736 2930 10798 2942
rect 10550 2797 10596 2812
rect 10550 2763 10556 2797
rect 10590 2763 10596 2797
rect 10550 2725 10596 2763
rect 10550 2691 10556 2725
rect 10590 2691 10596 2725
rect 10550 2653 10596 2691
rect 8550 2597 8644 2628
rect 8550 2545 8571 2597
rect 8623 2545 8644 2597
rect 8550 2514 8644 2545
rect 10550 2619 10556 2653
rect 10590 2619 10596 2653
rect 10550 2581 10596 2619
rect 10550 2547 10556 2581
rect 10590 2547 10596 2581
rect 8550 2428 8642 2514
rect 8550 2394 8579 2428
rect 8613 2394 8642 2428
rect 8550 2388 8642 2394
rect 10550 2509 10596 2547
rect 10550 2475 10556 2509
rect 10590 2475 10596 2509
rect 10550 2437 10596 2475
rect 10550 2403 10556 2437
rect 10590 2403 10596 2437
rect 10550 2365 10596 2403
rect 8232 2350 8440 2360
rect 8232 2316 8392 2350
rect 8426 2316 8440 2350
rect 8232 2298 8440 2316
rect 10550 2331 10556 2365
rect 10590 2331 10596 2365
rect 7846 2261 7852 2295
rect 7886 2261 7892 2295
rect 10550 2293 10596 2331
rect 7846 2223 7892 2261
rect 7846 2189 7852 2223
rect 7886 2189 7892 2223
rect 7846 2151 7892 2189
rect 7846 2117 7852 2151
rect 7886 2117 7892 2151
rect 7846 2079 7892 2117
rect 7846 2045 7852 2079
rect 7886 2045 7892 2079
rect 8494 2229 8540 2276
rect 8494 2195 8500 2229
rect 8534 2195 8540 2229
rect 8494 2157 8540 2195
rect 8494 2123 8500 2157
rect 8534 2123 8540 2157
rect 8494 2076 8540 2123
rect 8652 2229 8698 2276
rect 8652 2195 8658 2229
rect 8692 2195 8698 2229
rect 8652 2157 8698 2195
rect 8652 2123 8658 2157
rect 8692 2123 8698 2157
rect 8652 2076 8698 2123
rect 10550 2259 10556 2293
rect 10590 2259 10596 2293
rect 10550 2221 10596 2259
rect 10550 2187 10556 2221
rect 10590 2187 10596 2221
rect 10550 2149 10596 2187
rect 10550 2115 10556 2149
rect 10590 2115 10596 2149
rect 10550 2077 10596 2115
rect 7846 2007 7892 2045
rect 7846 1973 7852 2007
rect 7886 1973 7892 2007
rect 7846 1935 7892 1973
rect 7846 1901 7852 1935
rect 7886 1901 7892 1935
rect 7846 1863 7892 1901
rect 7846 1829 7852 1863
rect 7886 1829 7892 1863
rect 7846 1814 7892 1829
rect 10550 2043 10556 2077
rect 10590 2043 10596 2077
rect 10550 2005 10596 2043
rect 10550 1971 10556 2005
rect 10590 1971 10596 2005
rect 10550 1933 10596 1971
rect 10550 1899 10556 1933
rect 10590 1899 10596 1933
rect 10550 1861 10596 1899
rect 10550 1827 10556 1861
rect 10590 1827 10596 1861
rect 10550 1812 10596 1827
rect 10646 2797 10692 2812
rect 10646 2763 10652 2797
rect 10686 2763 10692 2797
rect 10646 2725 10692 2763
rect 10646 2691 10652 2725
rect 10686 2691 10692 2725
rect 10646 2653 10692 2691
rect 10646 2619 10652 2653
rect 10686 2619 10692 2653
rect 10646 2581 10692 2619
rect 10646 2547 10652 2581
rect 10686 2547 10692 2581
rect 10646 2509 10692 2547
rect 10646 2475 10652 2509
rect 10686 2475 10692 2509
rect 10646 2437 10692 2475
rect 10646 2403 10652 2437
rect 10686 2403 10692 2437
rect 10646 2365 10692 2403
rect 10646 2331 10652 2365
rect 10686 2331 10692 2365
rect 10646 2293 10692 2331
rect 10646 2259 10652 2293
rect 10686 2259 10692 2293
rect 10646 2221 10692 2259
rect 10646 2187 10652 2221
rect 10686 2187 10692 2221
rect 10646 2149 10692 2187
rect 10646 2115 10652 2149
rect 10686 2115 10692 2149
rect 10646 2077 10692 2115
rect 10646 2043 10652 2077
rect 10686 2043 10692 2077
rect 10646 2005 10692 2043
rect 10646 1971 10652 2005
rect 10686 1971 10692 2005
rect 10646 1933 10692 1971
rect 10646 1899 10652 1933
rect 10686 1899 10692 1933
rect 10646 1861 10692 1899
rect 10646 1827 10652 1861
rect 10686 1827 10692 1861
rect 10646 1812 10692 1827
rect 10742 2797 10788 2812
rect 10742 2763 10748 2797
rect 10782 2763 10788 2797
rect 10742 2725 10788 2763
rect 10742 2691 10748 2725
rect 10782 2691 10788 2725
rect 10742 2653 10788 2691
rect 10742 2619 10748 2653
rect 10782 2619 10788 2653
rect 10742 2581 10788 2619
rect 10742 2547 10748 2581
rect 10782 2547 10788 2581
rect 10742 2509 10788 2547
rect 10742 2475 10748 2509
rect 10782 2475 10788 2509
rect 10742 2437 10788 2475
rect 10742 2403 10748 2437
rect 10782 2403 10788 2437
rect 10742 2365 10788 2403
rect 10742 2331 10748 2365
rect 10782 2331 10788 2365
rect 10742 2293 10788 2331
rect 10742 2259 10748 2293
rect 10782 2259 10788 2293
rect 10742 2221 10788 2259
rect 10742 2187 10748 2221
rect 10782 2187 10788 2221
rect 10742 2149 10788 2187
rect 10742 2115 10748 2149
rect 10782 2115 10788 2149
rect 10742 2077 10788 2115
rect 10742 2043 10748 2077
rect 10782 2043 10788 2077
rect 10742 2005 10788 2043
rect 10742 1971 10748 2005
rect 10782 1971 10788 2005
rect 10742 1933 10788 1971
rect 10742 1899 10748 1933
rect 10782 1899 10788 1933
rect 10742 1861 10788 1899
rect 10742 1827 10748 1861
rect 10782 1827 10788 1861
rect 10742 1812 10788 1827
rect 10838 2797 10884 2812
rect 10838 2763 10844 2797
rect 10878 2763 10884 2797
rect 10838 2725 10884 2763
rect 10838 2691 10844 2725
rect 10878 2691 10884 2725
rect 10838 2653 10884 2691
rect 10838 2619 10844 2653
rect 10878 2619 10884 2653
rect 10838 2581 10884 2619
rect 10838 2547 10844 2581
rect 10878 2547 10884 2581
rect 10838 2509 10884 2547
rect 10838 2475 10844 2509
rect 10878 2475 10884 2509
rect 10838 2437 10884 2475
rect 10838 2403 10844 2437
rect 10878 2403 10884 2437
rect 10838 2365 10884 2403
rect 10838 2331 10844 2365
rect 10878 2331 10884 2365
rect 10838 2293 10884 2331
rect 10838 2259 10844 2293
rect 10878 2259 10884 2293
rect 10838 2221 10884 2259
rect 10838 2187 10844 2221
rect 10878 2187 10884 2221
rect 10838 2149 10884 2187
rect 10838 2115 10844 2149
rect 10878 2115 10884 2149
rect 10838 2077 10884 2115
rect 10838 2043 10844 2077
rect 10878 2043 10884 2077
rect 10838 2005 10884 2043
rect 10838 1971 10844 2005
rect 10878 1971 10884 2005
rect 10838 1933 10884 1971
rect 10838 1899 10844 1933
rect 10878 1899 10884 1933
rect 10838 1861 10884 1899
rect 10838 1827 10844 1861
rect 10878 1827 10884 1861
rect 10838 1812 10884 1827
rect 10934 2797 10980 2812
rect 10934 2763 10940 2797
rect 10974 2763 10980 2797
rect 10934 2725 10980 2763
rect 10934 2691 10940 2725
rect 10974 2691 10980 2725
rect 10934 2653 10980 2691
rect 10934 2619 10940 2653
rect 10974 2619 10980 2653
rect 10934 2581 10980 2619
rect 10934 2547 10940 2581
rect 10974 2547 10980 2581
rect 10934 2509 10980 2547
rect 10934 2475 10940 2509
rect 10974 2475 10980 2509
rect 10934 2437 10980 2475
rect 10934 2403 10940 2437
rect 10974 2403 10980 2437
rect 10934 2365 10980 2403
rect 10934 2331 10940 2365
rect 10974 2331 10980 2365
rect 10934 2293 10980 2331
rect 11232 2360 11294 2984
rect 13460 2972 13522 2984
rect 13460 2967 13856 2972
rect 13460 2915 13578 2967
rect 13630 2958 13856 2967
rect 13630 2924 13808 2958
rect 13842 2924 13856 2958
rect 13630 2915 13856 2924
rect 13460 2910 13856 2915
rect 13892 2950 13954 3112
rect 13892 2916 13904 2950
rect 13938 2916 13954 2950
rect 13892 2904 13954 2916
rect 13706 2771 13752 2786
rect 13706 2737 13712 2771
rect 13746 2737 13752 2771
rect 13706 2699 13752 2737
rect 13706 2665 13712 2699
rect 13746 2665 13752 2699
rect 13706 2627 13752 2665
rect 11550 2568 11642 2598
rect 11550 2516 11570 2568
rect 11622 2516 11642 2568
rect 11550 2428 11642 2516
rect 11550 2394 11579 2428
rect 11613 2394 11642 2428
rect 11550 2388 11642 2394
rect 13706 2593 13712 2627
rect 13746 2593 13752 2627
rect 13706 2555 13752 2593
rect 13706 2521 13712 2555
rect 13746 2521 13752 2555
rect 13706 2483 13752 2521
rect 13706 2449 13712 2483
rect 13746 2449 13752 2483
rect 13706 2411 13752 2449
rect 13706 2377 13712 2411
rect 13746 2377 13752 2411
rect 11232 2350 11440 2360
rect 11232 2316 11392 2350
rect 11426 2316 11440 2350
rect 11232 2298 11440 2316
rect 13706 2339 13752 2377
rect 13706 2305 13712 2339
rect 13746 2305 13752 2339
rect 10934 2259 10940 2293
rect 10974 2259 10980 2293
rect 10934 2221 10980 2259
rect 10934 2187 10940 2221
rect 10974 2187 10980 2221
rect 10934 2149 10980 2187
rect 10934 2115 10940 2149
rect 10974 2115 10980 2149
rect 10934 2077 10980 2115
rect 10934 2043 10940 2077
rect 10974 2043 10980 2077
rect 11494 2229 11540 2276
rect 11494 2195 11500 2229
rect 11534 2195 11540 2229
rect 11494 2157 11540 2195
rect 11494 2123 11500 2157
rect 11534 2123 11540 2157
rect 11494 2076 11540 2123
rect 11652 2229 11698 2276
rect 11652 2195 11658 2229
rect 11692 2195 11698 2229
rect 11652 2157 11698 2195
rect 11652 2123 11658 2157
rect 11692 2123 11698 2157
rect 11652 2076 11698 2123
rect 13706 2267 13752 2305
rect 13706 2233 13712 2267
rect 13746 2233 13752 2267
rect 13706 2195 13752 2233
rect 13706 2161 13712 2195
rect 13746 2161 13752 2195
rect 13706 2123 13752 2161
rect 13706 2089 13712 2123
rect 13746 2089 13752 2123
rect 10934 2005 10980 2043
rect 10934 1971 10940 2005
rect 10974 1971 10980 2005
rect 10934 1933 10980 1971
rect 10934 1899 10940 1933
rect 10974 1899 10980 1933
rect 10934 1861 10980 1899
rect 10934 1827 10940 1861
rect 10974 1827 10980 1861
rect 10934 1812 10980 1827
rect 13706 2051 13752 2089
rect 13706 2017 13712 2051
rect 13746 2017 13752 2051
rect 13706 1979 13752 2017
rect 13706 1945 13712 1979
rect 13746 1945 13752 1979
rect 13706 1907 13752 1945
rect 13706 1873 13712 1907
rect 13746 1873 13752 1907
rect 13706 1835 13752 1873
rect 13706 1801 13712 1835
rect 13746 1801 13752 1835
rect 13706 1786 13752 1801
rect 13802 2771 13848 2786
rect 13802 2737 13808 2771
rect 13842 2737 13848 2771
rect 13802 2699 13848 2737
rect 13802 2665 13808 2699
rect 13842 2665 13848 2699
rect 13802 2627 13848 2665
rect 13802 2593 13808 2627
rect 13842 2593 13848 2627
rect 13802 2555 13848 2593
rect 13802 2521 13808 2555
rect 13842 2521 13848 2555
rect 13802 2483 13848 2521
rect 13802 2449 13808 2483
rect 13842 2449 13848 2483
rect 13802 2411 13848 2449
rect 13802 2377 13808 2411
rect 13842 2377 13848 2411
rect 13802 2339 13848 2377
rect 13802 2305 13808 2339
rect 13842 2305 13848 2339
rect 13802 2267 13848 2305
rect 13802 2233 13808 2267
rect 13842 2233 13848 2267
rect 13802 2195 13848 2233
rect 13802 2161 13808 2195
rect 13842 2161 13848 2195
rect 13802 2123 13848 2161
rect 13802 2089 13808 2123
rect 13842 2089 13848 2123
rect 13802 2051 13848 2089
rect 13802 2017 13808 2051
rect 13842 2017 13848 2051
rect 13802 1979 13848 2017
rect 13802 1945 13808 1979
rect 13842 1945 13848 1979
rect 13802 1907 13848 1945
rect 13802 1873 13808 1907
rect 13842 1873 13848 1907
rect 13802 1835 13848 1873
rect 13802 1801 13808 1835
rect 13842 1801 13848 1835
rect 13802 1786 13848 1801
rect 13898 2771 13944 2786
rect 13898 2737 13904 2771
rect 13938 2737 13944 2771
rect 13898 2699 13944 2737
rect 13898 2665 13904 2699
rect 13938 2665 13944 2699
rect 13898 2627 13944 2665
rect 13898 2593 13904 2627
rect 13938 2593 13944 2627
rect 13898 2555 13944 2593
rect 13898 2521 13904 2555
rect 13938 2521 13944 2555
rect 13898 2483 13944 2521
rect 13898 2449 13904 2483
rect 13938 2449 13944 2483
rect 13898 2411 13944 2449
rect 13898 2377 13904 2411
rect 13938 2377 13944 2411
rect 13898 2339 13944 2377
rect 13898 2305 13904 2339
rect 13938 2305 13944 2339
rect 13898 2267 13944 2305
rect 13898 2233 13904 2267
rect 13938 2233 13944 2267
rect 13898 2195 13944 2233
rect 13898 2161 13904 2195
rect 13938 2161 13944 2195
rect 13898 2123 13944 2161
rect 13898 2089 13904 2123
rect 13938 2089 13944 2123
rect 13898 2051 13944 2089
rect 13898 2017 13904 2051
rect 13938 2017 13944 2051
rect 13898 1979 13944 2017
rect 13898 1945 13904 1979
rect 13938 1945 13944 1979
rect 13898 1907 13944 1945
rect 13898 1873 13904 1907
rect 13938 1873 13944 1907
rect 13898 1835 13944 1873
rect 13898 1801 13904 1835
rect 13938 1801 13944 1835
rect 13898 1786 13944 1801
rect 13994 2771 14040 2786
rect 13994 2737 14000 2771
rect 14034 2737 14040 2771
rect 13994 2699 14040 2737
rect 13994 2665 14000 2699
rect 14034 2665 14040 2699
rect 13994 2627 14040 2665
rect 13994 2593 14000 2627
rect 14034 2593 14040 2627
rect 13994 2555 14040 2593
rect 13994 2521 14000 2555
rect 14034 2521 14040 2555
rect 13994 2483 14040 2521
rect 13994 2449 14000 2483
rect 14034 2449 14040 2483
rect 13994 2411 14040 2449
rect 13994 2377 14000 2411
rect 14034 2377 14040 2411
rect 13994 2339 14040 2377
rect 13994 2305 14000 2339
rect 14034 2305 14040 2339
rect 13994 2267 14040 2305
rect 13994 2233 14000 2267
rect 14034 2233 14040 2267
rect 13994 2195 14040 2233
rect 13994 2161 14000 2195
rect 14034 2161 14040 2195
rect 13994 2123 14040 2161
rect 13994 2089 14000 2123
rect 14034 2089 14040 2123
rect 13994 2051 14040 2089
rect 13994 2017 14000 2051
rect 14034 2017 14040 2051
rect 13994 1979 14040 2017
rect 13994 1945 14000 1979
rect 14034 1945 14040 1979
rect 13994 1907 14040 1945
rect 13994 1873 14000 1907
rect 14034 1873 14040 1907
rect 13994 1835 14040 1873
rect 13994 1801 14000 1835
rect 14034 1801 14040 1835
rect 13994 1786 14040 1801
rect 14090 2771 14136 2786
rect 14090 2737 14096 2771
rect 14130 2737 14136 2771
rect 14090 2699 14136 2737
rect 14090 2665 14096 2699
rect 14130 2665 14136 2699
rect 14090 2627 14136 2665
rect 14090 2593 14096 2627
rect 14130 2593 14136 2627
rect 14090 2555 14136 2593
rect 14090 2521 14096 2555
rect 14130 2521 14136 2555
rect 14090 2483 14136 2521
rect 14090 2449 14096 2483
rect 14130 2449 14136 2483
rect 14090 2411 14136 2449
rect 14090 2377 14096 2411
rect 14130 2377 14136 2411
rect 14090 2339 14136 2377
rect 14090 2305 14096 2339
rect 14130 2305 14136 2339
rect 14090 2267 14136 2305
rect 14232 2360 14294 3112
rect 14550 2428 14642 3684
rect 14550 2394 14579 2428
rect 14613 2394 14642 2428
rect 14550 2388 14642 2394
rect 15332 3745 15566 3779
rect 15600 3745 15614 3779
rect 15332 3732 15614 3745
rect 15698 3760 15760 3772
rect 14232 2350 14442 2360
rect 14232 2316 14392 2350
rect 14426 2316 14442 2350
rect 14232 2298 14442 2316
rect 14090 2233 14096 2267
rect 14130 2233 14136 2267
rect 14090 2195 14136 2233
rect 14090 2161 14096 2195
rect 14130 2161 14136 2195
rect 14090 2123 14136 2161
rect 14090 2089 14096 2123
rect 14130 2089 14136 2123
rect 14090 2051 14136 2089
rect 14494 2229 14540 2276
rect 14494 2195 14500 2229
rect 14534 2195 14540 2229
rect 14494 2157 14540 2195
rect 14494 2123 14500 2157
rect 14534 2123 14540 2157
rect 14494 2076 14540 2123
rect 14652 2229 14698 2276
rect 14652 2195 14658 2229
rect 14692 2195 14698 2229
rect 14652 2157 14698 2195
rect 14652 2123 14658 2157
rect 14692 2123 14698 2157
rect 14652 2076 14698 2123
rect 14090 2017 14096 2051
rect 14130 2017 14136 2051
rect 14090 1979 14136 2017
rect 14090 1945 14096 1979
rect 14130 1945 14136 1979
rect 15332 1948 15394 3732
rect 15698 3726 15710 3760
rect 15744 3726 15760 3760
rect 16456 3768 16487 3820
rect 16539 3768 16894 3820
rect 16946 3821 17578 3840
rect 16946 3787 16974 3821
rect 17008 3787 17578 3821
rect 16946 3770 17578 3787
rect 16456 3742 16894 3768
rect 14090 1907 14136 1945
rect 14090 1873 14096 1907
rect 14130 1873 14136 1907
rect 14090 1835 14136 1873
rect 15314 1856 15324 1948
rect 15408 1856 15418 1948
rect 14090 1801 14096 1835
rect 14130 1801 14136 1835
rect 14090 1786 14136 1801
rect 1566 1696 1624 1708
rect 1566 1662 1578 1696
rect 1612 1662 1624 1696
rect 1566 1626 1624 1662
rect 4522 1680 4580 1692
rect 4522 1646 4534 1680
rect 4568 1646 4580 1680
rect 706 1546 2456 1626
rect 4522 1614 4580 1646
rect 7552 1680 7610 1692
rect 7552 1646 7564 1680
rect 7598 1646 7610 1680
rect 3674 1612 5408 1614
rect 706 1458 798 1546
rect 706 1424 734 1458
rect 768 1424 798 1458
rect 706 1404 798 1424
rect 2382 1452 2456 1546
rect 2382 1418 2400 1452
rect 2434 1418 2456 1452
rect 2382 1404 2456 1418
rect 3672 1530 5408 1612
rect 7552 1610 7610 1646
rect 10640 1678 10698 1690
rect 10640 1644 10652 1678
rect 10686 1644 10698 1678
rect 10640 1612 10698 1644
rect 13796 1652 13854 1664
rect 13796 1618 13808 1652
rect 13842 1618 13854 1652
rect 3672 1442 3746 1530
rect 3672 1408 3690 1442
rect 3724 1408 3746 1442
rect 3672 1390 3746 1408
rect 5332 1436 5408 1530
rect 5332 1402 5356 1436
rect 5390 1402 5408 1436
rect 5332 1388 5408 1402
rect 6700 1524 8436 1610
rect 6700 1442 6776 1524
rect 6700 1408 6720 1442
rect 6754 1408 6776 1442
rect 6700 1384 6776 1408
rect 8360 1436 8436 1524
rect 8360 1402 8386 1436
rect 8420 1402 8436 1436
rect 8360 1378 8436 1402
rect 9788 1526 11530 1612
rect 13796 1592 13854 1618
rect 9788 1440 9864 1526
rect 9788 1406 9808 1440
rect 9842 1406 9864 1440
rect 9788 1380 9864 1406
rect 11452 1434 11530 1526
rect 11452 1400 11474 1434
rect 11508 1400 11530 1434
rect 11452 1388 11530 1400
rect 12940 1510 14684 1592
rect 12940 1414 13018 1510
rect 12940 1380 12964 1414
rect 12998 1380 13018 1414
rect 12940 1354 13018 1380
rect 14608 1408 14684 1510
rect 14608 1374 14630 1408
rect 14664 1374 14684 1408
rect 14608 1358 14684 1374
rect 15332 1380 15394 1856
rect 15452 1670 15548 1692
rect 15452 1618 15471 1670
rect 15523 1618 15548 1670
rect 15452 1596 15548 1618
rect 15452 1492 15514 1596
rect 15452 1458 15466 1492
rect 15500 1458 15514 1492
rect 15452 1444 15514 1458
rect 15332 1370 15468 1380
rect -1110 1264 -1095 1298
rect -1061 1264 -1048 1298
rect -1110 1256 -1048 1264
rect -916 1298 -420 1354
rect 15332 1336 15422 1370
rect 15456 1336 15468 1370
rect 15332 1328 15468 1336
rect 15332 1326 15394 1328
rect -916 1264 -899 1298
rect -865 1264 -420 1298
rect -916 1238 -420 1264
rect -1692 1051 -1646 1066
rect -1692 1017 -1686 1051
rect -1652 1017 -1646 1051
rect -1692 979 -1646 1017
rect -1692 945 -1686 979
rect -1652 945 -1646 979
rect -1692 907 -1646 945
rect -1692 873 -1686 907
rect -1652 873 -1646 907
rect -1692 835 -1646 873
rect -1692 801 -1686 835
rect -1652 801 -1646 835
rect -1692 763 -1646 801
rect -1692 729 -1686 763
rect -1652 729 -1646 763
rect -1692 691 -1646 729
rect -1692 657 -1686 691
rect -1652 657 -1646 691
rect -1692 619 -1646 657
rect -1692 585 -1686 619
rect -1652 585 -1646 619
rect -1692 547 -1646 585
rect -1692 513 -1686 547
rect -1652 513 -1646 547
rect -1692 475 -1646 513
rect -1692 441 -1686 475
rect -1652 441 -1646 475
rect -1692 403 -1646 441
rect -1692 369 -1686 403
rect -1652 369 -1646 403
rect -1692 331 -1646 369
rect -1692 297 -1686 331
rect -1652 297 -1646 331
rect -1692 259 -1646 297
rect -1692 225 -1686 259
rect -1652 225 -1646 259
rect -1692 187 -1646 225
rect -1692 153 -1686 187
rect -1652 153 -1646 187
rect -1692 115 -1646 153
rect -1692 81 -1686 115
rect -1652 81 -1646 115
rect -1692 66 -1646 81
rect -1594 1051 -1548 1066
rect -1594 1017 -1588 1051
rect -1554 1017 -1548 1051
rect -1594 979 -1548 1017
rect -1594 945 -1588 979
rect -1554 945 -1548 979
rect -1594 907 -1548 945
rect -1594 873 -1588 907
rect -1554 873 -1548 907
rect -1594 835 -1548 873
rect -1594 801 -1588 835
rect -1554 801 -1548 835
rect -1594 763 -1548 801
rect -1594 729 -1588 763
rect -1554 729 -1548 763
rect -1594 691 -1548 729
rect -1594 657 -1588 691
rect -1554 657 -1548 691
rect -1594 619 -1548 657
rect -1594 585 -1588 619
rect -1554 585 -1548 619
rect -1594 547 -1548 585
rect -1594 513 -1588 547
rect -1554 513 -1548 547
rect -1594 475 -1548 513
rect -1594 441 -1588 475
rect -1554 441 -1548 475
rect -1594 403 -1548 441
rect -1594 369 -1588 403
rect -1554 369 -1548 403
rect -1594 331 -1548 369
rect -1594 297 -1588 331
rect -1554 297 -1548 331
rect -1594 259 -1548 297
rect -1594 225 -1588 259
rect -1554 225 -1548 259
rect -1594 187 -1548 225
rect -1594 153 -1588 187
rect -1554 153 -1548 187
rect -1594 115 -1548 153
rect -1594 81 -1588 115
rect -1554 81 -1548 115
rect -1594 66 -1548 81
rect -1496 1051 -1450 1066
rect -1496 1017 -1490 1051
rect -1456 1017 -1450 1051
rect -1496 979 -1450 1017
rect -1496 945 -1490 979
rect -1456 945 -1450 979
rect -1496 907 -1450 945
rect -1496 873 -1490 907
rect -1456 873 -1450 907
rect -1496 835 -1450 873
rect -1496 801 -1490 835
rect -1456 801 -1450 835
rect -1496 763 -1450 801
rect -1496 729 -1490 763
rect -1456 729 -1450 763
rect -1496 691 -1450 729
rect -1496 657 -1490 691
rect -1456 657 -1450 691
rect -1496 619 -1450 657
rect -1496 585 -1490 619
rect -1456 585 -1450 619
rect -1496 547 -1450 585
rect -1496 513 -1490 547
rect -1456 513 -1450 547
rect -1496 475 -1450 513
rect -1496 441 -1490 475
rect -1456 441 -1450 475
rect -1496 403 -1450 441
rect -1496 369 -1490 403
rect -1456 369 -1450 403
rect -1496 331 -1450 369
rect -1496 297 -1490 331
rect -1456 297 -1450 331
rect -1496 259 -1450 297
rect -1496 225 -1490 259
rect -1456 225 -1450 259
rect -1496 187 -1450 225
rect -1496 153 -1490 187
rect -1456 153 -1450 187
rect -1496 115 -1450 153
rect -1496 81 -1490 115
rect -1456 81 -1450 115
rect -1496 66 -1450 81
rect -1398 1051 -1352 1066
rect -1398 1017 -1392 1051
rect -1358 1017 -1352 1051
rect -1398 979 -1352 1017
rect -1398 945 -1392 979
rect -1358 945 -1352 979
rect -1398 907 -1352 945
rect -1398 873 -1392 907
rect -1358 873 -1352 907
rect -1398 835 -1352 873
rect -1398 801 -1392 835
rect -1358 801 -1352 835
rect -1398 763 -1352 801
rect -1398 729 -1392 763
rect -1358 729 -1352 763
rect -1398 691 -1352 729
rect -1398 657 -1392 691
rect -1358 657 -1352 691
rect -1398 619 -1352 657
rect -1398 585 -1392 619
rect -1358 585 -1352 619
rect -1398 547 -1352 585
rect -1398 513 -1392 547
rect -1358 513 -1352 547
rect -1398 475 -1352 513
rect -1398 441 -1392 475
rect -1358 441 -1352 475
rect -1398 403 -1352 441
rect -1398 369 -1392 403
rect -1358 369 -1352 403
rect -1398 331 -1352 369
rect -1398 297 -1392 331
rect -1358 297 -1352 331
rect -1398 259 -1352 297
rect -1398 225 -1392 259
rect -1358 225 -1352 259
rect -1398 187 -1352 225
rect -1398 153 -1392 187
rect -1358 153 -1352 187
rect -1398 115 -1352 153
rect -1398 81 -1392 115
rect -1358 81 -1352 115
rect -1398 66 -1352 81
rect -1300 1051 -1254 1066
rect -1300 1017 -1294 1051
rect -1260 1017 -1254 1051
rect -1300 979 -1254 1017
rect -1300 945 -1294 979
rect -1260 945 -1254 979
rect -1300 907 -1254 945
rect -1300 873 -1294 907
rect -1260 873 -1254 907
rect -1300 835 -1254 873
rect -1300 801 -1294 835
rect -1260 801 -1254 835
rect -1300 763 -1254 801
rect -1300 729 -1294 763
rect -1260 729 -1254 763
rect -1300 691 -1254 729
rect -1300 657 -1294 691
rect -1260 657 -1254 691
rect -1300 619 -1254 657
rect -1300 585 -1294 619
rect -1260 585 -1254 619
rect -1300 547 -1254 585
rect -1300 513 -1294 547
rect -1260 513 -1254 547
rect -1300 475 -1254 513
rect -1300 441 -1294 475
rect -1260 441 -1254 475
rect -1300 403 -1254 441
rect -1300 369 -1294 403
rect -1260 369 -1254 403
rect -1300 331 -1254 369
rect -1300 297 -1294 331
rect -1260 297 -1254 331
rect -1300 259 -1254 297
rect -1300 225 -1294 259
rect -1260 225 -1254 259
rect -1300 187 -1254 225
rect -1300 153 -1294 187
rect -1260 153 -1254 187
rect -1300 115 -1254 153
rect -1300 81 -1294 115
rect -1260 81 -1254 115
rect -1300 66 -1254 81
rect -1202 1051 -1156 1066
rect -1202 1017 -1196 1051
rect -1162 1017 -1156 1051
rect -1202 979 -1156 1017
rect -1202 945 -1196 979
rect -1162 945 -1156 979
rect -1202 907 -1156 945
rect -1202 873 -1196 907
rect -1162 873 -1156 907
rect -1202 835 -1156 873
rect -1202 801 -1196 835
rect -1162 801 -1156 835
rect -1202 763 -1156 801
rect -1202 729 -1196 763
rect -1162 729 -1156 763
rect -1202 691 -1156 729
rect -1202 657 -1196 691
rect -1162 657 -1156 691
rect -1202 619 -1156 657
rect -1202 585 -1196 619
rect -1162 585 -1156 619
rect -1202 547 -1156 585
rect -1202 513 -1196 547
rect -1162 513 -1156 547
rect -1202 475 -1156 513
rect -1202 441 -1196 475
rect -1162 441 -1156 475
rect -1202 403 -1156 441
rect -1202 369 -1196 403
rect -1162 369 -1156 403
rect -1202 331 -1156 369
rect -1202 297 -1196 331
rect -1162 297 -1156 331
rect -1202 259 -1156 297
rect -1202 225 -1196 259
rect -1162 225 -1156 259
rect -1202 187 -1156 225
rect -1202 153 -1196 187
rect -1162 153 -1156 187
rect -1202 115 -1156 153
rect -1202 81 -1196 115
rect -1162 81 -1156 115
rect -1202 66 -1156 81
rect -1104 1051 -1058 1066
rect -1104 1017 -1098 1051
rect -1064 1017 -1058 1051
rect -1104 979 -1058 1017
rect -1104 945 -1098 979
rect -1064 945 -1058 979
rect -1104 907 -1058 945
rect -1104 873 -1098 907
rect -1064 873 -1058 907
rect -1104 835 -1058 873
rect -1104 801 -1098 835
rect -1064 801 -1058 835
rect -1104 763 -1058 801
rect -1104 729 -1098 763
rect -1064 729 -1058 763
rect -1104 691 -1058 729
rect -1104 657 -1098 691
rect -1064 657 -1058 691
rect -1104 619 -1058 657
rect -1104 585 -1098 619
rect -1064 585 -1058 619
rect -1104 547 -1058 585
rect -1104 513 -1098 547
rect -1064 513 -1058 547
rect -1104 475 -1058 513
rect -1104 441 -1098 475
rect -1064 441 -1058 475
rect -1104 403 -1058 441
rect -1104 369 -1098 403
rect -1064 369 -1058 403
rect -1104 331 -1058 369
rect -1104 297 -1098 331
rect -1064 297 -1058 331
rect -1104 259 -1058 297
rect -1104 225 -1098 259
rect -1064 225 -1058 259
rect -1104 187 -1058 225
rect -1104 153 -1098 187
rect -1064 153 -1058 187
rect -1104 115 -1058 153
rect -1104 81 -1098 115
rect -1064 81 -1058 115
rect -1104 66 -1058 81
rect -1006 1051 -960 1066
rect -1006 1017 -1000 1051
rect -966 1017 -960 1051
rect -1006 979 -960 1017
rect -1006 945 -1000 979
rect -966 945 -960 979
rect -1006 907 -960 945
rect -1006 873 -1000 907
rect -966 873 -960 907
rect -1006 835 -960 873
rect -1006 801 -1000 835
rect -966 801 -960 835
rect -1006 763 -960 801
rect -1006 729 -1000 763
rect -966 729 -960 763
rect -1006 691 -960 729
rect -1006 657 -1000 691
rect -966 657 -960 691
rect -1006 619 -960 657
rect -1006 585 -1000 619
rect -966 585 -960 619
rect -1006 547 -960 585
rect -1006 513 -1000 547
rect -966 513 -960 547
rect -1006 475 -960 513
rect -1006 441 -1000 475
rect -966 441 -960 475
rect -1006 403 -960 441
rect -1006 369 -1000 403
rect -966 369 -960 403
rect -1006 331 -960 369
rect -1006 297 -1000 331
rect -966 297 -960 331
rect -1006 259 -960 297
rect -1006 225 -1000 259
rect -966 225 -960 259
rect -1006 187 -960 225
rect -1006 153 -1000 187
rect -966 153 -960 187
rect -1006 115 -960 153
rect -1006 81 -1000 115
rect -966 81 -960 115
rect -1006 66 -960 81
rect -908 1051 -862 1066
rect -908 1017 -902 1051
rect -868 1017 -862 1051
rect -908 979 -862 1017
rect -908 945 -902 979
rect -868 945 -862 979
rect -908 907 -862 945
rect -908 873 -902 907
rect -868 873 -862 907
rect -908 835 -862 873
rect -908 801 -902 835
rect -868 801 -862 835
rect -908 763 -862 801
rect -908 729 -902 763
rect -868 729 -862 763
rect -908 691 -862 729
rect -908 657 -902 691
rect -868 657 -862 691
rect -908 619 -862 657
rect -908 585 -902 619
rect -868 585 -862 619
rect -908 547 -862 585
rect -908 513 -902 547
rect -868 513 -862 547
rect -908 475 -862 513
rect -908 441 -902 475
rect -868 441 -862 475
rect -908 403 -862 441
rect -908 369 -902 403
rect -868 369 -862 403
rect -908 331 -862 369
rect -908 297 -902 331
rect -868 297 -862 331
rect -908 259 -862 297
rect -908 225 -902 259
rect -868 225 -862 259
rect -908 187 -862 225
rect -908 153 -902 187
rect -868 153 -862 187
rect -908 115 -862 153
rect -908 81 -902 115
rect -868 81 -862 115
rect -908 66 -862 81
rect -560 -126 -420 1238
rect 152 1253 198 1268
rect 152 1219 158 1253
rect 192 1219 198 1253
rect 152 1181 198 1219
rect 152 1147 158 1181
rect 192 1147 198 1181
rect 152 1109 198 1147
rect 152 1075 158 1109
rect 192 1075 198 1109
rect 152 1037 198 1075
rect 152 1003 158 1037
rect 192 1003 198 1037
rect 152 965 198 1003
rect 152 931 158 965
rect 192 931 198 965
rect 152 893 198 931
rect 152 859 158 893
rect 192 859 198 893
rect 152 821 198 859
rect 152 787 158 821
rect 192 787 198 821
rect 152 749 198 787
rect 152 715 158 749
rect 192 715 198 749
rect 152 677 198 715
rect 152 643 158 677
rect 192 643 198 677
rect 152 605 198 643
rect 152 571 158 605
rect 192 571 198 605
rect 152 533 198 571
rect 152 499 158 533
rect 192 499 198 533
rect 152 461 198 499
rect 152 427 158 461
rect 192 427 198 461
rect 152 389 198 427
rect 152 355 158 389
rect 192 355 198 389
rect 152 317 198 355
rect 152 283 158 317
rect 192 283 198 317
rect 152 268 198 283
rect 248 1253 294 1268
rect 248 1219 254 1253
rect 288 1219 294 1253
rect 248 1181 294 1219
rect 248 1147 254 1181
rect 288 1147 294 1181
rect 248 1109 294 1147
rect 248 1075 254 1109
rect 288 1075 294 1109
rect 248 1037 294 1075
rect 248 1003 254 1037
rect 288 1003 294 1037
rect 248 965 294 1003
rect 248 931 254 965
rect 288 931 294 965
rect 248 893 294 931
rect 248 859 254 893
rect 288 859 294 893
rect 248 821 294 859
rect 248 787 254 821
rect 288 787 294 821
rect 248 749 294 787
rect 248 715 254 749
rect 288 715 294 749
rect 248 677 294 715
rect 248 643 254 677
rect 288 643 294 677
rect 248 605 294 643
rect 248 571 254 605
rect 288 571 294 605
rect 248 533 294 571
rect 248 499 254 533
rect 288 499 294 533
rect 248 461 294 499
rect 248 427 254 461
rect 288 427 294 461
rect 248 389 294 427
rect 248 355 254 389
rect 288 355 294 389
rect 248 317 294 355
rect 248 283 254 317
rect 288 283 294 317
rect 248 268 294 283
rect 344 1253 390 1268
rect 344 1219 350 1253
rect 384 1219 390 1253
rect 344 1181 390 1219
rect 344 1147 350 1181
rect 384 1147 390 1181
rect 344 1109 390 1147
rect 344 1075 350 1109
rect 384 1075 390 1109
rect 344 1037 390 1075
rect 344 1003 350 1037
rect 384 1003 390 1037
rect 344 965 390 1003
rect 344 931 350 965
rect 384 931 390 965
rect 344 893 390 931
rect 344 859 350 893
rect 384 859 390 893
rect 344 821 390 859
rect 344 787 350 821
rect 384 787 390 821
rect 344 749 390 787
rect 344 715 350 749
rect 384 715 390 749
rect 344 677 390 715
rect 344 643 350 677
rect 384 643 390 677
rect 344 605 390 643
rect 344 571 350 605
rect 384 571 390 605
rect 344 533 390 571
rect 344 499 350 533
rect 384 499 390 533
rect 344 461 390 499
rect 344 427 350 461
rect 384 427 390 461
rect 344 389 390 427
rect 344 355 350 389
rect 384 355 390 389
rect 344 317 390 355
rect 344 283 350 317
rect 384 283 390 317
rect 344 268 390 283
rect 440 1253 486 1268
rect 440 1219 446 1253
rect 480 1219 486 1253
rect 440 1181 486 1219
rect 440 1147 446 1181
rect 480 1147 486 1181
rect 440 1109 486 1147
rect 440 1075 446 1109
rect 480 1075 486 1109
rect 440 1037 486 1075
rect 440 1003 446 1037
rect 480 1003 486 1037
rect 440 965 486 1003
rect 440 931 446 965
rect 480 931 486 965
rect 440 893 486 931
rect 440 859 446 893
rect 480 859 486 893
rect 440 821 486 859
rect 440 787 446 821
rect 480 787 486 821
rect 440 749 486 787
rect 440 715 446 749
rect 480 715 486 749
rect 440 677 486 715
rect 440 643 446 677
rect 480 643 486 677
rect 440 605 486 643
rect 440 571 446 605
rect 480 571 486 605
rect 440 533 486 571
rect 440 499 446 533
rect 480 499 486 533
rect 440 461 486 499
rect 440 427 446 461
rect 480 427 486 461
rect 440 389 486 427
rect 440 355 446 389
rect 480 355 486 389
rect 440 317 486 355
rect 440 283 446 317
rect 480 283 486 317
rect 440 268 486 283
rect 536 1253 582 1268
rect 536 1219 542 1253
rect 576 1219 582 1253
rect 536 1181 582 1219
rect 536 1147 542 1181
rect 576 1147 582 1181
rect 536 1109 582 1147
rect 536 1075 542 1109
rect 576 1075 582 1109
rect 536 1037 582 1075
rect 536 1003 542 1037
rect 576 1003 582 1037
rect 536 965 582 1003
rect 536 931 542 965
rect 576 931 582 965
rect 536 893 582 931
rect 536 859 542 893
rect 576 859 582 893
rect 536 821 582 859
rect 536 787 542 821
rect 576 787 582 821
rect 536 749 582 787
rect 536 715 542 749
rect 576 715 582 749
rect 536 677 582 715
rect 536 643 542 677
rect 576 643 582 677
rect 536 605 582 643
rect 536 571 542 605
rect 576 571 582 605
rect 536 533 582 571
rect 536 499 542 533
rect 576 499 582 533
rect 536 461 582 499
rect 536 427 542 461
rect 576 427 582 461
rect 536 389 582 427
rect 536 355 542 389
rect 576 355 582 389
rect 536 317 582 355
rect 536 283 542 317
rect 576 283 582 317
rect 536 268 582 283
rect 632 1253 678 1268
rect 632 1219 638 1253
rect 672 1219 678 1253
rect 632 1181 678 1219
rect 632 1147 638 1181
rect 672 1147 678 1181
rect 632 1109 678 1147
rect 632 1075 638 1109
rect 672 1075 678 1109
rect 632 1037 678 1075
rect 632 1003 638 1037
rect 672 1003 678 1037
rect 632 965 678 1003
rect 632 931 638 965
rect 672 931 678 965
rect 632 893 678 931
rect 632 859 638 893
rect 672 859 678 893
rect 632 821 678 859
rect 632 787 638 821
rect 672 787 678 821
rect 632 749 678 787
rect 632 715 638 749
rect 672 715 678 749
rect 632 677 678 715
rect 632 643 638 677
rect 672 643 678 677
rect 632 605 678 643
rect 632 571 638 605
rect 672 571 678 605
rect 632 533 678 571
rect 632 499 638 533
rect 672 499 678 533
rect 632 461 678 499
rect 632 427 638 461
rect 672 427 678 461
rect 632 389 678 427
rect 632 355 638 389
rect 672 355 678 389
rect 632 317 678 355
rect 632 283 638 317
rect 672 283 678 317
rect 632 268 678 283
rect 728 1253 774 1268
rect 728 1219 734 1253
rect 768 1219 774 1253
rect 728 1181 774 1219
rect 728 1147 734 1181
rect 768 1147 774 1181
rect 728 1109 774 1147
rect 728 1075 734 1109
rect 768 1075 774 1109
rect 728 1037 774 1075
rect 728 1003 734 1037
rect 768 1003 774 1037
rect 728 965 774 1003
rect 728 931 734 965
rect 768 931 774 965
rect 728 893 774 931
rect 728 859 734 893
rect 768 859 774 893
rect 728 821 774 859
rect 728 787 734 821
rect 768 787 774 821
rect 728 749 774 787
rect 728 715 734 749
rect 768 715 774 749
rect 728 677 774 715
rect 728 643 734 677
rect 768 643 774 677
rect 728 605 774 643
rect 728 571 734 605
rect 768 571 774 605
rect 728 533 774 571
rect 728 499 734 533
rect 768 499 774 533
rect 728 461 774 499
rect 728 427 734 461
rect 768 427 774 461
rect 728 389 774 427
rect 728 355 734 389
rect 768 355 774 389
rect 728 317 774 355
rect 728 283 734 317
rect 768 283 774 317
rect 728 268 774 283
rect 824 1253 870 1268
rect 824 1219 830 1253
rect 864 1219 870 1253
rect 824 1181 870 1219
rect 824 1147 830 1181
rect 864 1147 870 1181
rect 824 1109 870 1147
rect 824 1075 830 1109
rect 864 1075 870 1109
rect 824 1037 870 1075
rect 824 1003 830 1037
rect 864 1003 870 1037
rect 824 965 870 1003
rect 824 931 830 965
rect 864 931 870 965
rect 824 893 870 931
rect 824 859 830 893
rect 864 859 870 893
rect 824 821 870 859
rect 824 787 830 821
rect 864 787 870 821
rect 824 749 870 787
rect 824 715 830 749
rect 864 715 870 749
rect 824 677 870 715
rect 824 643 830 677
rect 864 643 870 677
rect 824 605 870 643
rect 824 571 830 605
rect 864 571 870 605
rect 824 533 870 571
rect 824 499 830 533
rect 864 499 870 533
rect 824 461 870 499
rect 824 427 830 461
rect 864 427 870 461
rect 824 389 870 427
rect 824 355 830 389
rect 864 355 870 389
rect 824 317 870 355
rect 824 283 830 317
rect 864 283 870 317
rect 824 268 870 283
rect 920 1253 966 1268
rect 920 1219 926 1253
rect 960 1219 966 1253
rect 920 1181 966 1219
rect 920 1147 926 1181
rect 960 1147 966 1181
rect 920 1109 966 1147
rect 920 1075 926 1109
rect 960 1075 966 1109
rect 920 1037 966 1075
rect 920 1003 926 1037
rect 960 1003 966 1037
rect 920 965 966 1003
rect 920 931 926 965
rect 960 931 966 965
rect 920 893 966 931
rect 920 859 926 893
rect 960 859 966 893
rect 920 821 966 859
rect 920 787 926 821
rect 960 787 966 821
rect 920 749 966 787
rect 920 715 926 749
rect 960 715 966 749
rect 920 677 966 715
rect 920 643 926 677
rect 960 643 966 677
rect 920 605 966 643
rect 920 571 926 605
rect 960 571 966 605
rect 920 533 966 571
rect 920 499 926 533
rect 960 499 966 533
rect 920 461 966 499
rect 920 427 926 461
rect 960 427 966 461
rect 920 389 966 427
rect 920 355 926 389
rect 960 355 966 389
rect 920 317 966 355
rect 920 283 926 317
rect 960 283 966 317
rect 920 268 966 283
rect 1016 1253 1062 1268
rect 1016 1219 1022 1253
rect 1056 1219 1062 1253
rect 1016 1181 1062 1219
rect 1016 1147 1022 1181
rect 1056 1147 1062 1181
rect 1016 1109 1062 1147
rect 1016 1075 1022 1109
rect 1056 1075 1062 1109
rect 1016 1037 1062 1075
rect 1016 1003 1022 1037
rect 1056 1003 1062 1037
rect 1016 965 1062 1003
rect 1016 931 1022 965
rect 1056 931 1062 965
rect 1016 893 1062 931
rect 1016 859 1022 893
rect 1056 859 1062 893
rect 1016 821 1062 859
rect 1016 787 1022 821
rect 1056 787 1062 821
rect 1016 749 1062 787
rect 1016 715 1022 749
rect 1056 715 1062 749
rect 1016 677 1062 715
rect 1016 643 1022 677
rect 1056 643 1062 677
rect 1016 605 1062 643
rect 1016 571 1022 605
rect 1056 571 1062 605
rect 1016 533 1062 571
rect 1016 499 1022 533
rect 1056 499 1062 533
rect 1016 461 1062 499
rect 1016 427 1022 461
rect 1056 427 1062 461
rect 1016 389 1062 427
rect 1016 355 1022 389
rect 1056 355 1062 389
rect 1016 317 1062 355
rect 1016 283 1022 317
rect 1056 283 1062 317
rect 1016 268 1062 283
rect 1112 1253 1158 1268
rect 1112 1219 1118 1253
rect 1152 1219 1158 1253
rect 1112 1181 1158 1219
rect 1112 1147 1118 1181
rect 1152 1147 1158 1181
rect 1112 1109 1158 1147
rect 1112 1075 1118 1109
rect 1152 1075 1158 1109
rect 1112 1037 1158 1075
rect 1112 1003 1118 1037
rect 1152 1003 1158 1037
rect 1112 965 1158 1003
rect 1112 931 1118 965
rect 1152 931 1158 965
rect 1112 893 1158 931
rect 1112 859 1118 893
rect 1152 859 1158 893
rect 1112 821 1158 859
rect 1112 787 1118 821
rect 1152 787 1158 821
rect 1112 749 1158 787
rect 1112 715 1118 749
rect 1152 715 1158 749
rect 1112 677 1158 715
rect 1112 643 1118 677
rect 1152 643 1158 677
rect 1112 605 1158 643
rect 1112 571 1118 605
rect 1152 571 1158 605
rect 1112 533 1158 571
rect 1112 499 1118 533
rect 1152 499 1158 533
rect 1112 461 1158 499
rect 1112 427 1118 461
rect 1152 427 1158 461
rect 1112 389 1158 427
rect 1112 355 1118 389
rect 1152 355 1158 389
rect 1112 317 1158 355
rect 1112 283 1118 317
rect 1152 283 1158 317
rect 1112 268 1158 283
rect 1208 1253 1254 1268
rect 1208 1219 1214 1253
rect 1248 1219 1254 1253
rect 1208 1181 1254 1219
rect 1208 1147 1214 1181
rect 1248 1147 1254 1181
rect 1208 1109 1254 1147
rect 1208 1075 1214 1109
rect 1248 1075 1254 1109
rect 1208 1037 1254 1075
rect 1208 1003 1214 1037
rect 1248 1003 1254 1037
rect 1208 965 1254 1003
rect 1208 931 1214 965
rect 1248 931 1254 965
rect 1208 893 1254 931
rect 1208 859 1214 893
rect 1248 859 1254 893
rect 1208 821 1254 859
rect 1208 787 1214 821
rect 1248 787 1254 821
rect 1208 749 1254 787
rect 1208 715 1214 749
rect 1248 715 1254 749
rect 1208 677 1254 715
rect 1208 643 1214 677
rect 1248 643 1254 677
rect 1208 605 1254 643
rect 1208 571 1214 605
rect 1248 571 1254 605
rect 1208 533 1254 571
rect 1208 499 1214 533
rect 1248 499 1254 533
rect 1208 461 1254 499
rect 1208 427 1214 461
rect 1248 427 1254 461
rect 1208 389 1254 427
rect 1208 355 1214 389
rect 1248 355 1254 389
rect 1208 317 1254 355
rect 1208 283 1214 317
rect 1248 283 1254 317
rect 1208 268 1254 283
rect 1304 1253 1350 1268
rect 1304 1219 1310 1253
rect 1344 1219 1350 1253
rect 1304 1181 1350 1219
rect 1304 1147 1310 1181
rect 1344 1147 1350 1181
rect 1304 1109 1350 1147
rect 1304 1075 1310 1109
rect 1344 1075 1350 1109
rect 1304 1037 1350 1075
rect 1304 1003 1310 1037
rect 1344 1003 1350 1037
rect 1304 965 1350 1003
rect 1304 931 1310 965
rect 1344 931 1350 965
rect 1304 893 1350 931
rect 1304 859 1310 893
rect 1344 859 1350 893
rect 1304 821 1350 859
rect 1304 787 1310 821
rect 1344 787 1350 821
rect 1304 749 1350 787
rect 1304 715 1310 749
rect 1344 715 1350 749
rect 1304 677 1350 715
rect 1304 643 1310 677
rect 1344 643 1350 677
rect 1304 605 1350 643
rect 1304 571 1310 605
rect 1344 571 1350 605
rect 1304 533 1350 571
rect 1304 499 1310 533
rect 1344 499 1350 533
rect 1304 461 1350 499
rect 1304 427 1310 461
rect 1344 427 1350 461
rect 1304 389 1350 427
rect 1304 355 1310 389
rect 1344 355 1350 389
rect 1304 317 1350 355
rect 1304 283 1310 317
rect 1344 283 1350 317
rect 1304 268 1350 283
rect 1920 1253 1966 1268
rect 1920 1219 1926 1253
rect 1960 1219 1966 1253
rect 1920 1181 1966 1219
rect 1920 1147 1926 1181
rect 1960 1147 1966 1181
rect 1920 1109 1966 1147
rect 1920 1075 1926 1109
rect 1960 1075 1966 1109
rect 1920 1037 1966 1075
rect 1920 1003 1926 1037
rect 1960 1003 1966 1037
rect 1920 965 1966 1003
rect 1920 931 1926 965
rect 1960 931 1966 965
rect 1920 893 1966 931
rect 1920 859 1926 893
rect 1960 859 1966 893
rect 1920 821 1966 859
rect 1920 787 1926 821
rect 1960 787 1966 821
rect 1920 749 1966 787
rect 1920 715 1926 749
rect 1960 715 1966 749
rect 1920 677 1966 715
rect 1920 643 1926 677
rect 1960 643 1966 677
rect 1920 605 1966 643
rect 1920 571 1926 605
rect 1960 571 1966 605
rect 1920 533 1966 571
rect 1920 499 1926 533
rect 1960 499 1966 533
rect 1920 461 1966 499
rect 1920 427 1926 461
rect 1960 427 1966 461
rect 1920 389 1966 427
rect 1920 355 1926 389
rect 1960 355 1966 389
rect 1920 317 1966 355
rect 1920 283 1926 317
rect 1960 283 1966 317
rect 1920 268 1966 283
rect 2016 1253 2062 1268
rect 2016 1219 2022 1253
rect 2056 1219 2062 1253
rect 2016 1181 2062 1219
rect 2016 1147 2022 1181
rect 2056 1147 2062 1181
rect 2016 1109 2062 1147
rect 2016 1075 2022 1109
rect 2056 1075 2062 1109
rect 2016 1037 2062 1075
rect 2016 1003 2022 1037
rect 2056 1003 2062 1037
rect 2016 965 2062 1003
rect 2016 931 2022 965
rect 2056 931 2062 965
rect 2016 893 2062 931
rect 2016 859 2022 893
rect 2056 859 2062 893
rect 2016 821 2062 859
rect 2016 787 2022 821
rect 2056 787 2062 821
rect 2016 749 2062 787
rect 2016 715 2022 749
rect 2056 715 2062 749
rect 2016 677 2062 715
rect 2016 643 2022 677
rect 2056 643 2062 677
rect 2016 605 2062 643
rect 2016 571 2022 605
rect 2056 571 2062 605
rect 2016 533 2062 571
rect 2016 499 2022 533
rect 2056 499 2062 533
rect 2016 461 2062 499
rect 2016 427 2022 461
rect 2056 427 2062 461
rect 2016 389 2062 427
rect 2016 355 2022 389
rect 2056 355 2062 389
rect 2016 317 2062 355
rect 2016 283 2022 317
rect 2056 283 2062 317
rect 2016 268 2062 283
rect 2112 1253 2158 1268
rect 2112 1219 2118 1253
rect 2152 1219 2158 1253
rect 2112 1181 2158 1219
rect 2112 1147 2118 1181
rect 2152 1147 2158 1181
rect 2112 1109 2158 1147
rect 2112 1075 2118 1109
rect 2152 1075 2158 1109
rect 2112 1037 2158 1075
rect 2112 1003 2118 1037
rect 2152 1003 2158 1037
rect 2112 965 2158 1003
rect 2112 931 2118 965
rect 2152 931 2158 965
rect 2112 893 2158 931
rect 2112 859 2118 893
rect 2152 859 2158 893
rect 2112 821 2158 859
rect 2112 787 2118 821
rect 2152 787 2158 821
rect 2112 749 2158 787
rect 2112 715 2118 749
rect 2152 715 2158 749
rect 2112 677 2158 715
rect 2112 643 2118 677
rect 2152 643 2158 677
rect 2112 605 2158 643
rect 2112 571 2118 605
rect 2152 571 2158 605
rect 2112 533 2158 571
rect 2112 499 2118 533
rect 2152 499 2158 533
rect 2112 461 2158 499
rect 2112 427 2118 461
rect 2152 427 2158 461
rect 2112 389 2158 427
rect 2112 355 2118 389
rect 2152 355 2158 389
rect 2112 317 2158 355
rect 2112 283 2118 317
rect 2152 283 2158 317
rect 2112 268 2158 283
rect 2208 1253 2254 1268
rect 2208 1219 2214 1253
rect 2248 1219 2254 1253
rect 2208 1181 2254 1219
rect 2208 1147 2214 1181
rect 2248 1147 2254 1181
rect 2208 1109 2254 1147
rect 2208 1075 2214 1109
rect 2248 1075 2254 1109
rect 2208 1037 2254 1075
rect 2208 1003 2214 1037
rect 2248 1003 2254 1037
rect 2208 965 2254 1003
rect 2208 931 2214 965
rect 2248 931 2254 965
rect 2208 893 2254 931
rect 2208 859 2214 893
rect 2248 859 2254 893
rect 2208 821 2254 859
rect 2208 787 2214 821
rect 2248 787 2254 821
rect 2208 749 2254 787
rect 2208 715 2214 749
rect 2248 715 2254 749
rect 2208 677 2254 715
rect 2208 643 2214 677
rect 2248 643 2254 677
rect 2208 605 2254 643
rect 2208 571 2214 605
rect 2248 571 2254 605
rect 2208 533 2254 571
rect 2208 499 2214 533
rect 2248 499 2254 533
rect 2208 461 2254 499
rect 2208 427 2214 461
rect 2248 427 2254 461
rect 2208 389 2254 427
rect 2208 355 2214 389
rect 2248 355 2254 389
rect 2208 317 2254 355
rect 2208 283 2214 317
rect 2248 283 2254 317
rect 2208 268 2254 283
rect 2304 1253 2350 1268
rect 2304 1219 2310 1253
rect 2344 1219 2350 1253
rect 2304 1181 2350 1219
rect 2304 1147 2310 1181
rect 2344 1147 2350 1181
rect 2304 1109 2350 1147
rect 2304 1075 2310 1109
rect 2344 1075 2350 1109
rect 2304 1037 2350 1075
rect 2304 1003 2310 1037
rect 2344 1003 2350 1037
rect 2304 965 2350 1003
rect 2304 931 2310 965
rect 2344 931 2350 965
rect 2304 893 2350 931
rect 2304 859 2310 893
rect 2344 859 2350 893
rect 2304 821 2350 859
rect 2304 787 2310 821
rect 2344 787 2350 821
rect 2304 749 2350 787
rect 2304 715 2310 749
rect 2344 715 2350 749
rect 2304 677 2350 715
rect 2304 643 2310 677
rect 2344 643 2350 677
rect 2304 605 2350 643
rect 2304 571 2310 605
rect 2344 571 2350 605
rect 2304 533 2350 571
rect 2304 499 2310 533
rect 2344 499 2350 533
rect 2304 461 2350 499
rect 2304 427 2310 461
rect 2344 427 2350 461
rect 2304 389 2350 427
rect 2304 355 2310 389
rect 2344 355 2350 389
rect 2304 317 2350 355
rect 2304 283 2310 317
rect 2344 283 2350 317
rect 2304 268 2350 283
rect 2400 1253 2446 1268
rect 2400 1219 2406 1253
rect 2440 1219 2446 1253
rect 2400 1181 2446 1219
rect 2400 1147 2406 1181
rect 2440 1147 2446 1181
rect 2400 1109 2446 1147
rect 2400 1075 2406 1109
rect 2440 1075 2446 1109
rect 2400 1037 2446 1075
rect 2400 1003 2406 1037
rect 2440 1003 2446 1037
rect 2400 965 2446 1003
rect 2400 931 2406 965
rect 2440 931 2446 965
rect 2400 893 2446 931
rect 2400 859 2406 893
rect 2440 859 2446 893
rect 2400 821 2446 859
rect 2400 787 2406 821
rect 2440 787 2446 821
rect 2400 749 2446 787
rect 2400 715 2406 749
rect 2440 715 2446 749
rect 2400 677 2446 715
rect 2400 643 2406 677
rect 2440 643 2446 677
rect 2400 605 2446 643
rect 2400 571 2406 605
rect 2440 571 2446 605
rect 2400 533 2446 571
rect 2400 499 2406 533
rect 2440 499 2446 533
rect 2400 461 2446 499
rect 2400 427 2406 461
rect 2440 427 2446 461
rect 2400 389 2446 427
rect 2400 355 2406 389
rect 2440 355 2446 389
rect 2400 317 2446 355
rect 2400 283 2406 317
rect 2440 283 2446 317
rect 2400 268 2446 283
rect 2496 1253 2542 1268
rect 2496 1219 2502 1253
rect 2536 1219 2542 1253
rect 2496 1181 2542 1219
rect 2496 1147 2502 1181
rect 2536 1147 2542 1181
rect 2496 1109 2542 1147
rect 2496 1075 2502 1109
rect 2536 1075 2542 1109
rect 2496 1037 2542 1075
rect 2496 1003 2502 1037
rect 2536 1003 2542 1037
rect 2496 965 2542 1003
rect 2496 931 2502 965
rect 2536 931 2542 965
rect 2496 893 2542 931
rect 2496 859 2502 893
rect 2536 859 2542 893
rect 2496 821 2542 859
rect 2496 787 2502 821
rect 2536 787 2542 821
rect 2496 749 2542 787
rect 2496 715 2502 749
rect 2536 715 2542 749
rect 2496 677 2542 715
rect 2496 643 2502 677
rect 2536 643 2542 677
rect 2496 605 2542 643
rect 2496 571 2502 605
rect 2536 571 2542 605
rect 2496 533 2542 571
rect 2496 499 2502 533
rect 2536 499 2542 533
rect 2496 461 2542 499
rect 2496 427 2502 461
rect 2536 427 2542 461
rect 2496 389 2542 427
rect 2496 355 2502 389
rect 2536 355 2542 389
rect 2496 317 2542 355
rect 2496 283 2502 317
rect 2536 283 2542 317
rect 2496 268 2542 283
rect 2592 1253 2638 1268
rect 2592 1219 2598 1253
rect 2632 1219 2638 1253
rect 2592 1181 2638 1219
rect 2592 1147 2598 1181
rect 2632 1147 2638 1181
rect 2592 1109 2638 1147
rect 2592 1075 2598 1109
rect 2632 1075 2638 1109
rect 2592 1037 2638 1075
rect 2592 1003 2598 1037
rect 2632 1003 2638 1037
rect 2592 965 2638 1003
rect 2592 931 2598 965
rect 2632 931 2638 965
rect 2592 893 2638 931
rect 2592 859 2598 893
rect 2632 859 2638 893
rect 2592 821 2638 859
rect 2592 787 2598 821
rect 2632 787 2638 821
rect 2592 749 2638 787
rect 2592 715 2598 749
rect 2632 715 2638 749
rect 2592 677 2638 715
rect 2592 643 2598 677
rect 2632 643 2638 677
rect 2592 605 2638 643
rect 2592 571 2598 605
rect 2632 571 2638 605
rect 2592 533 2638 571
rect 2592 499 2598 533
rect 2632 499 2638 533
rect 2592 461 2638 499
rect 2592 427 2598 461
rect 2632 427 2638 461
rect 2592 389 2638 427
rect 2592 355 2598 389
rect 2632 355 2638 389
rect 2592 317 2638 355
rect 2592 283 2598 317
rect 2632 283 2638 317
rect 2592 268 2638 283
rect 2688 1253 2734 1268
rect 2688 1219 2694 1253
rect 2728 1219 2734 1253
rect 2688 1181 2734 1219
rect 2688 1147 2694 1181
rect 2728 1147 2734 1181
rect 2688 1109 2734 1147
rect 2688 1075 2694 1109
rect 2728 1075 2734 1109
rect 2688 1037 2734 1075
rect 2688 1003 2694 1037
rect 2728 1003 2734 1037
rect 2688 965 2734 1003
rect 2688 931 2694 965
rect 2728 931 2734 965
rect 2688 893 2734 931
rect 2688 859 2694 893
rect 2728 859 2734 893
rect 2688 821 2734 859
rect 2688 787 2694 821
rect 2728 787 2734 821
rect 2688 749 2734 787
rect 2688 715 2694 749
rect 2728 715 2734 749
rect 2688 677 2734 715
rect 2688 643 2694 677
rect 2728 643 2734 677
rect 2688 605 2734 643
rect 2688 571 2694 605
rect 2728 571 2734 605
rect 2688 533 2734 571
rect 2688 499 2694 533
rect 2728 499 2734 533
rect 2688 461 2734 499
rect 2688 427 2694 461
rect 2728 427 2734 461
rect 2688 389 2734 427
rect 2688 355 2694 389
rect 2728 355 2734 389
rect 2688 317 2734 355
rect 2688 283 2694 317
rect 2728 283 2734 317
rect 2688 268 2734 283
rect 2784 1253 2830 1268
rect 2784 1219 2790 1253
rect 2824 1219 2830 1253
rect 2784 1181 2830 1219
rect 2784 1147 2790 1181
rect 2824 1147 2830 1181
rect 2784 1109 2830 1147
rect 2784 1075 2790 1109
rect 2824 1075 2830 1109
rect 2784 1037 2830 1075
rect 2784 1003 2790 1037
rect 2824 1003 2830 1037
rect 2784 965 2830 1003
rect 2784 931 2790 965
rect 2824 931 2830 965
rect 2784 893 2830 931
rect 2784 859 2790 893
rect 2824 859 2830 893
rect 2784 821 2830 859
rect 2784 787 2790 821
rect 2824 787 2830 821
rect 2784 749 2830 787
rect 2784 715 2790 749
rect 2824 715 2830 749
rect 2784 677 2830 715
rect 2784 643 2790 677
rect 2824 643 2830 677
rect 2784 605 2830 643
rect 2784 571 2790 605
rect 2824 571 2830 605
rect 2784 533 2830 571
rect 2784 499 2790 533
rect 2824 499 2830 533
rect 2784 461 2830 499
rect 2784 427 2790 461
rect 2824 427 2830 461
rect 2784 389 2830 427
rect 2784 355 2790 389
rect 2824 355 2830 389
rect 2784 317 2830 355
rect 2784 283 2790 317
rect 2824 283 2830 317
rect 2784 268 2830 283
rect 2880 1253 2926 1268
rect 2880 1219 2886 1253
rect 2920 1219 2926 1253
rect 2880 1181 2926 1219
rect 2880 1147 2886 1181
rect 2920 1147 2926 1181
rect 2880 1109 2926 1147
rect 2880 1075 2886 1109
rect 2920 1075 2926 1109
rect 2880 1037 2926 1075
rect 2880 1003 2886 1037
rect 2920 1003 2926 1037
rect 2880 965 2926 1003
rect 2880 931 2886 965
rect 2920 931 2926 965
rect 2880 893 2926 931
rect 2880 859 2886 893
rect 2920 859 2926 893
rect 2880 821 2926 859
rect 2880 787 2886 821
rect 2920 787 2926 821
rect 2880 749 2926 787
rect 2880 715 2886 749
rect 2920 715 2926 749
rect 2880 677 2926 715
rect 2880 643 2886 677
rect 2920 643 2926 677
rect 2880 605 2926 643
rect 2880 571 2886 605
rect 2920 571 2926 605
rect 2880 533 2926 571
rect 2880 499 2886 533
rect 2920 499 2926 533
rect 2880 461 2926 499
rect 2880 427 2886 461
rect 2920 427 2926 461
rect 2880 389 2926 427
rect 2880 355 2886 389
rect 2920 355 2926 389
rect 2880 317 2926 355
rect 2880 283 2886 317
rect 2920 283 2926 317
rect 2880 268 2926 283
rect 2976 1253 3022 1268
rect 2976 1219 2982 1253
rect 3016 1219 3022 1253
rect 15416 1257 15462 1300
rect 2976 1181 3022 1219
rect 2976 1147 2982 1181
rect 3016 1147 3022 1181
rect 2976 1109 3022 1147
rect 2976 1075 2982 1109
rect 3016 1075 3022 1109
rect 2976 1037 3022 1075
rect 2976 1003 2982 1037
rect 3016 1003 3022 1037
rect 2976 965 3022 1003
rect 2976 931 2982 965
rect 3016 931 3022 965
rect 2976 893 3022 931
rect 2976 859 2982 893
rect 3016 859 3022 893
rect 2976 821 3022 859
rect 2976 787 2982 821
rect 3016 787 3022 821
rect 2976 749 3022 787
rect 2976 715 2982 749
rect 3016 715 3022 749
rect 2976 677 3022 715
rect 2976 643 2982 677
rect 3016 643 3022 677
rect 2976 605 3022 643
rect 2976 571 2982 605
rect 3016 571 3022 605
rect 2976 533 3022 571
rect 2976 499 2982 533
rect 3016 499 3022 533
rect 2976 461 3022 499
rect 2976 427 2982 461
rect 3016 427 3022 461
rect 2976 389 3022 427
rect 2976 355 2982 389
rect 3016 355 3022 389
rect 2976 317 3022 355
rect 2976 283 2982 317
rect 3016 283 3022 317
rect 2976 268 3022 283
rect 3108 1237 3154 1252
rect 3108 1203 3114 1237
rect 3148 1203 3154 1237
rect 3108 1165 3154 1203
rect 3108 1131 3114 1165
rect 3148 1131 3154 1165
rect 3108 1093 3154 1131
rect 3108 1059 3114 1093
rect 3148 1059 3154 1093
rect 3108 1021 3154 1059
rect 3108 987 3114 1021
rect 3148 987 3154 1021
rect 3108 949 3154 987
rect 3108 915 3114 949
rect 3148 915 3154 949
rect 3108 877 3154 915
rect 3108 843 3114 877
rect 3148 843 3154 877
rect 3108 805 3154 843
rect 3108 771 3114 805
rect 3148 771 3154 805
rect 3108 733 3154 771
rect 3108 699 3114 733
rect 3148 699 3154 733
rect 3108 661 3154 699
rect 3108 627 3114 661
rect 3148 627 3154 661
rect 3108 589 3154 627
rect 3108 555 3114 589
rect 3148 555 3154 589
rect 3108 517 3154 555
rect 3108 483 3114 517
rect 3148 483 3154 517
rect 3108 445 3154 483
rect 3108 411 3114 445
rect 3148 411 3154 445
rect 3108 373 3154 411
rect 3108 339 3114 373
rect 3148 339 3154 373
rect 3108 301 3154 339
rect 3108 267 3114 301
rect 3148 267 3154 301
rect 3108 252 3154 267
rect 3204 1237 3250 1252
rect 3204 1203 3210 1237
rect 3244 1203 3250 1237
rect 3204 1165 3250 1203
rect 3204 1131 3210 1165
rect 3244 1131 3250 1165
rect 3204 1093 3250 1131
rect 3204 1059 3210 1093
rect 3244 1059 3250 1093
rect 3204 1021 3250 1059
rect 3204 987 3210 1021
rect 3244 987 3250 1021
rect 3204 949 3250 987
rect 3204 915 3210 949
rect 3244 915 3250 949
rect 3204 877 3250 915
rect 3204 843 3210 877
rect 3244 843 3250 877
rect 3204 805 3250 843
rect 3204 771 3210 805
rect 3244 771 3250 805
rect 3204 733 3250 771
rect 3204 699 3210 733
rect 3244 699 3250 733
rect 3204 661 3250 699
rect 3204 627 3210 661
rect 3244 627 3250 661
rect 3204 589 3250 627
rect 3204 555 3210 589
rect 3244 555 3250 589
rect 3204 517 3250 555
rect 3204 483 3210 517
rect 3244 483 3250 517
rect 3204 445 3250 483
rect 3204 411 3210 445
rect 3244 411 3250 445
rect 3204 373 3250 411
rect 3204 339 3210 373
rect 3244 339 3250 373
rect 3204 301 3250 339
rect 3204 267 3210 301
rect 3244 267 3250 301
rect 3204 252 3250 267
rect 3300 1237 3346 1252
rect 3300 1203 3306 1237
rect 3340 1203 3346 1237
rect 3300 1165 3346 1203
rect 3300 1131 3306 1165
rect 3340 1131 3346 1165
rect 3300 1093 3346 1131
rect 3300 1059 3306 1093
rect 3340 1059 3346 1093
rect 3300 1021 3346 1059
rect 3300 987 3306 1021
rect 3340 987 3346 1021
rect 3300 949 3346 987
rect 3300 915 3306 949
rect 3340 915 3346 949
rect 3300 877 3346 915
rect 3300 843 3306 877
rect 3340 843 3346 877
rect 3300 805 3346 843
rect 3300 771 3306 805
rect 3340 771 3346 805
rect 3300 733 3346 771
rect 3300 699 3306 733
rect 3340 699 3346 733
rect 3300 661 3346 699
rect 3300 627 3306 661
rect 3340 627 3346 661
rect 3300 589 3346 627
rect 3300 555 3306 589
rect 3340 555 3346 589
rect 3300 517 3346 555
rect 3300 483 3306 517
rect 3340 483 3346 517
rect 3300 445 3346 483
rect 3300 411 3306 445
rect 3340 411 3346 445
rect 3300 373 3346 411
rect 3300 339 3306 373
rect 3340 339 3346 373
rect 3300 301 3346 339
rect 3300 267 3306 301
rect 3340 267 3346 301
rect 3300 252 3346 267
rect 3396 1237 3442 1252
rect 3396 1203 3402 1237
rect 3436 1203 3442 1237
rect 3396 1165 3442 1203
rect 3396 1131 3402 1165
rect 3436 1131 3442 1165
rect 3396 1093 3442 1131
rect 3396 1059 3402 1093
rect 3436 1059 3442 1093
rect 3396 1021 3442 1059
rect 3396 987 3402 1021
rect 3436 987 3442 1021
rect 3396 949 3442 987
rect 3396 915 3402 949
rect 3436 915 3442 949
rect 3396 877 3442 915
rect 3396 843 3402 877
rect 3436 843 3442 877
rect 3396 805 3442 843
rect 3396 771 3402 805
rect 3436 771 3442 805
rect 3396 733 3442 771
rect 3396 699 3402 733
rect 3436 699 3442 733
rect 3396 661 3442 699
rect 3396 627 3402 661
rect 3436 627 3442 661
rect 3396 589 3442 627
rect 3396 555 3402 589
rect 3436 555 3442 589
rect 3396 517 3442 555
rect 3396 483 3402 517
rect 3436 483 3442 517
rect 3396 445 3442 483
rect 3396 411 3402 445
rect 3436 411 3442 445
rect 3396 373 3442 411
rect 3396 339 3402 373
rect 3436 339 3442 373
rect 3396 301 3442 339
rect 3396 267 3402 301
rect 3436 267 3442 301
rect 3396 252 3442 267
rect 3492 1237 3538 1252
rect 3492 1203 3498 1237
rect 3532 1203 3538 1237
rect 3492 1165 3538 1203
rect 3492 1131 3498 1165
rect 3532 1131 3538 1165
rect 3492 1093 3538 1131
rect 3492 1059 3498 1093
rect 3532 1059 3538 1093
rect 3492 1021 3538 1059
rect 3492 987 3498 1021
rect 3532 987 3538 1021
rect 3492 949 3538 987
rect 3492 915 3498 949
rect 3532 915 3538 949
rect 3492 877 3538 915
rect 3492 843 3498 877
rect 3532 843 3538 877
rect 3492 805 3538 843
rect 3492 771 3498 805
rect 3532 771 3538 805
rect 3492 733 3538 771
rect 3492 699 3498 733
rect 3532 699 3538 733
rect 3492 661 3538 699
rect 3492 627 3498 661
rect 3532 627 3538 661
rect 3492 589 3538 627
rect 3492 555 3498 589
rect 3532 555 3538 589
rect 3492 517 3538 555
rect 3492 483 3498 517
rect 3532 483 3538 517
rect 3492 445 3538 483
rect 3492 411 3498 445
rect 3532 411 3538 445
rect 3492 373 3538 411
rect 3492 339 3498 373
rect 3532 339 3538 373
rect 3492 301 3538 339
rect 3492 267 3498 301
rect 3532 267 3538 301
rect 3492 252 3538 267
rect 3588 1237 3634 1252
rect 3588 1203 3594 1237
rect 3628 1203 3634 1237
rect 3588 1165 3634 1203
rect 3588 1131 3594 1165
rect 3628 1131 3634 1165
rect 3588 1093 3634 1131
rect 3588 1059 3594 1093
rect 3628 1059 3634 1093
rect 3588 1021 3634 1059
rect 3588 987 3594 1021
rect 3628 987 3634 1021
rect 3588 949 3634 987
rect 3588 915 3594 949
rect 3628 915 3634 949
rect 3588 877 3634 915
rect 3588 843 3594 877
rect 3628 843 3634 877
rect 3588 805 3634 843
rect 3588 771 3594 805
rect 3628 771 3634 805
rect 3588 733 3634 771
rect 3588 699 3594 733
rect 3628 699 3634 733
rect 3588 661 3634 699
rect 3588 627 3594 661
rect 3628 627 3634 661
rect 3588 589 3634 627
rect 3588 555 3594 589
rect 3628 555 3634 589
rect 3588 517 3634 555
rect 3588 483 3594 517
rect 3628 483 3634 517
rect 3588 445 3634 483
rect 3588 411 3594 445
rect 3628 411 3634 445
rect 3588 373 3634 411
rect 3588 339 3594 373
rect 3628 339 3634 373
rect 3588 301 3634 339
rect 3588 267 3594 301
rect 3628 267 3634 301
rect 3588 252 3634 267
rect 3684 1237 3730 1252
rect 3684 1203 3690 1237
rect 3724 1203 3730 1237
rect 3684 1165 3730 1203
rect 3684 1131 3690 1165
rect 3724 1131 3730 1165
rect 3684 1093 3730 1131
rect 3684 1059 3690 1093
rect 3724 1059 3730 1093
rect 3684 1021 3730 1059
rect 3684 987 3690 1021
rect 3724 987 3730 1021
rect 3684 949 3730 987
rect 3684 915 3690 949
rect 3724 915 3730 949
rect 3684 877 3730 915
rect 3684 843 3690 877
rect 3724 843 3730 877
rect 3684 805 3730 843
rect 3684 771 3690 805
rect 3724 771 3730 805
rect 3684 733 3730 771
rect 3684 699 3690 733
rect 3724 699 3730 733
rect 3684 661 3730 699
rect 3684 627 3690 661
rect 3724 627 3730 661
rect 3684 589 3730 627
rect 3684 555 3690 589
rect 3724 555 3730 589
rect 3684 517 3730 555
rect 3684 483 3690 517
rect 3724 483 3730 517
rect 3684 445 3730 483
rect 3684 411 3690 445
rect 3724 411 3730 445
rect 3684 373 3730 411
rect 3684 339 3690 373
rect 3724 339 3730 373
rect 3684 301 3730 339
rect 3684 267 3690 301
rect 3724 267 3730 301
rect 3684 252 3730 267
rect 3780 1237 3826 1252
rect 3780 1203 3786 1237
rect 3820 1203 3826 1237
rect 3780 1165 3826 1203
rect 3780 1131 3786 1165
rect 3820 1131 3826 1165
rect 3780 1093 3826 1131
rect 3780 1059 3786 1093
rect 3820 1059 3826 1093
rect 3780 1021 3826 1059
rect 3780 987 3786 1021
rect 3820 987 3826 1021
rect 3780 949 3826 987
rect 3780 915 3786 949
rect 3820 915 3826 949
rect 3780 877 3826 915
rect 3780 843 3786 877
rect 3820 843 3826 877
rect 3780 805 3826 843
rect 3780 771 3786 805
rect 3820 771 3826 805
rect 3780 733 3826 771
rect 3780 699 3786 733
rect 3820 699 3826 733
rect 3780 661 3826 699
rect 3780 627 3786 661
rect 3820 627 3826 661
rect 3780 589 3826 627
rect 3780 555 3786 589
rect 3820 555 3826 589
rect 3780 517 3826 555
rect 3780 483 3786 517
rect 3820 483 3826 517
rect 3780 445 3826 483
rect 3780 411 3786 445
rect 3820 411 3826 445
rect 3780 373 3826 411
rect 3780 339 3786 373
rect 3820 339 3826 373
rect 3780 301 3826 339
rect 3780 267 3786 301
rect 3820 267 3826 301
rect 3780 252 3826 267
rect 3876 1237 3922 1252
rect 3876 1203 3882 1237
rect 3916 1203 3922 1237
rect 3876 1165 3922 1203
rect 3876 1131 3882 1165
rect 3916 1131 3922 1165
rect 3876 1093 3922 1131
rect 3876 1059 3882 1093
rect 3916 1059 3922 1093
rect 3876 1021 3922 1059
rect 3876 987 3882 1021
rect 3916 987 3922 1021
rect 3876 949 3922 987
rect 3876 915 3882 949
rect 3916 915 3922 949
rect 3876 877 3922 915
rect 3876 843 3882 877
rect 3916 843 3922 877
rect 3876 805 3922 843
rect 3876 771 3882 805
rect 3916 771 3922 805
rect 3876 733 3922 771
rect 3876 699 3882 733
rect 3916 699 3922 733
rect 3876 661 3922 699
rect 3876 627 3882 661
rect 3916 627 3922 661
rect 3876 589 3922 627
rect 3876 555 3882 589
rect 3916 555 3922 589
rect 3876 517 3922 555
rect 3876 483 3882 517
rect 3916 483 3922 517
rect 3876 445 3922 483
rect 3876 411 3882 445
rect 3916 411 3922 445
rect 3876 373 3922 411
rect 3876 339 3882 373
rect 3916 339 3922 373
rect 3876 301 3922 339
rect 3876 267 3882 301
rect 3916 267 3922 301
rect 3876 252 3922 267
rect 3972 1237 4018 1252
rect 3972 1203 3978 1237
rect 4012 1203 4018 1237
rect 3972 1165 4018 1203
rect 3972 1131 3978 1165
rect 4012 1131 4018 1165
rect 3972 1093 4018 1131
rect 3972 1059 3978 1093
rect 4012 1059 4018 1093
rect 3972 1021 4018 1059
rect 3972 987 3978 1021
rect 4012 987 4018 1021
rect 3972 949 4018 987
rect 3972 915 3978 949
rect 4012 915 4018 949
rect 3972 877 4018 915
rect 3972 843 3978 877
rect 4012 843 4018 877
rect 3972 805 4018 843
rect 3972 771 3978 805
rect 4012 771 4018 805
rect 3972 733 4018 771
rect 3972 699 3978 733
rect 4012 699 4018 733
rect 3972 661 4018 699
rect 3972 627 3978 661
rect 4012 627 4018 661
rect 3972 589 4018 627
rect 3972 555 3978 589
rect 4012 555 4018 589
rect 3972 517 4018 555
rect 3972 483 3978 517
rect 4012 483 4018 517
rect 3972 445 4018 483
rect 3972 411 3978 445
rect 4012 411 4018 445
rect 3972 373 4018 411
rect 3972 339 3978 373
rect 4012 339 4018 373
rect 3972 301 4018 339
rect 3972 267 3978 301
rect 4012 267 4018 301
rect 3972 252 4018 267
rect 4068 1237 4114 1252
rect 4068 1203 4074 1237
rect 4108 1203 4114 1237
rect 4068 1165 4114 1203
rect 4068 1131 4074 1165
rect 4108 1131 4114 1165
rect 4068 1093 4114 1131
rect 4068 1059 4074 1093
rect 4108 1059 4114 1093
rect 4068 1021 4114 1059
rect 4068 987 4074 1021
rect 4108 987 4114 1021
rect 4068 949 4114 987
rect 4068 915 4074 949
rect 4108 915 4114 949
rect 4068 877 4114 915
rect 4068 843 4074 877
rect 4108 843 4114 877
rect 4068 805 4114 843
rect 4068 771 4074 805
rect 4108 771 4114 805
rect 4068 733 4114 771
rect 4068 699 4074 733
rect 4108 699 4114 733
rect 4068 661 4114 699
rect 4068 627 4074 661
rect 4108 627 4114 661
rect 4068 589 4114 627
rect 4068 555 4074 589
rect 4108 555 4114 589
rect 4068 517 4114 555
rect 4068 483 4074 517
rect 4108 483 4114 517
rect 4068 445 4114 483
rect 4068 411 4074 445
rect 4108 411 4114 445
rect 4068 373 4114 411
rect 4068 339 4074 373
rect 4108 339 4114 373
rect 4068 301 4114 339
rect 4068 267 4074 301
rect 4108 267 4114 301
rect 4068 252 4114 267
rect 4164 1237 4210 1252
rect 4164 1203 4170 1237
rect 4204 1203 4210 1237
rect 4164 1165 4210 1203
rect 4164 1131 4170 1165
rect 4204 1131 4210 1165
rect 4164 1093 4210 1131
rect 4164 1059 4170 1093
rect 4204 1059 4210 1093
rect 4164 1021 4210 1059
rect 4164 987 4170 1021
rect 4204 987 4210 1021
rect 4164 949 4210 987
rect 4164 915 4170 949
rect 4204 915 4210 949
rect 4164 877 4210 915
rect 4164 843 4170 877
rect 4204 843 4210 877
rect 4164 805 4210 843
rect 4164 771 4170 805
rect 4204 771 4210 805
rect 4164 733 4210 771
rect 4164 699 4170 733
rect 4204 699 4210 733
rect 4164 661 4210 699
rect 4164 627 4170 661
rect 4204 627 4210 661
rect 4164 589 4210 627
rect 4164 555 4170 589
rect 4204 555 4210 589
rect 4164 517 4210 555
rect 4164 483 4170 517
rect 4204 483 4210 517
rect 4164 445 4210 483
rect 4164 411 4170 445
rect 4204 411 4210 445
rect 4164 373 4210 411
rect 4164 339 4170 373
rect 4204 339 4210 373
rect 4164 301 4210 339
rect 4164 267 4170 301
rect 4204 267 4210 301
rect 4164 252 4210 267
rect 4260 1237 4306 1252
rect 4260 1203 4266 1237
rect 4300 1203 4306 1237
rect 4260 1165 4306 1203
rect 4260 1131 4266 1165
rect 4300 1131 4306 1165
rect 4260 1093 4306 1131
rect 4260 1059 4266 1093
rect 4300 1059 4306 1093
rect 4260 1021 4306 1059
rect 4260 987 4266 1021
rect 4300 987 4306 1021
rect 4260 949 4306 987
rect 4260 915 4266 949
rect 4300 915 4306 949
rect 4260 877 4306 915
rect 4260 843 4266 877
rect 4300 843 4306 877
rect 4260 805 4306 843
rect 4260 771 4266 805
rect 4300 771 4306 805
rect 4260 733 4306 771
rect 4260 699 4266 733
rect 4300 699 4306 733
rect 4260 661 4306 699
rect 4260 627 4266 661
rect 4300 627 4306 661
rect 4260 589 4306 627
rect 4260 555 4266 589
rect 4300 555 4306 589
rect 4260 517 4306 555
rect 4260 483 4266 517
rect 4300 483 4306 517
rect 4260 445 4306 483
rect 4260 411 4266 445
rect 4300 411 4306 445
rect 4260 373 4306 411
rect 4260 339 4266 373
rect 4300 339 4306 373
rect 4260 301 4306 339
rect 4260 267 4266 301
rect 4300 267 4306 301
rect 4260 252 4306 267
rect 4876 1237 4922 1252
rect 4876 1203 4882 1237
rect 4916 1203 4922 1237
rect 4876 1165 4922 1203
rect 4876 1131 4882 1165
rect 4916 1131 4922 1165
rect 4876 1093 4922 1131
rect 4876 1059 4882 1093
rect 4916 1059 4922 1093
rect 4876 1021 4922 1059
rect 4876 987 4882 1021
rect 4916 987 4922 1021
rect 4876 949 4922 987
rect 4876 915 4882 949
rect 4916 915 4922 949
rect 4876 877 4922 915
rect 4876 843 4882 877
rect 4916 843 4922 877
rect 4876 805 4922 843
rect 4876 771 4882 805
rect 4916 771 4922 805
rect 4876 733 4922 771
rect 4876 699 4882 733
rect 4916 699 4922 733
rect 4876 661 4922 699
rect 4876 627 4882 661
rect 4916 627 4922 661
rect 4876 589 4922 627
rect 4876 555 4882 589
rect 4916 555 4922 589
rect 4876 517 4922 555
rect 4876 483 4882 517
rect 4916 483 4922 517
rect 4876 445 4922 483
rect 4876 411 4882 445
rect 4916 411 4922 445
rect 4876 373 4922 411
rect 4876 339 4882 373
rect 4916 339 4922 373
rect 4876 301 4922 339
rect 4876 267 4882 301
rect 4916 267 4922 301
rect 4876 252 4922 267
rect 4972 1237 5018 1252
rect 4972 1203 4978 1237
rect 5012 1203 5018 1237
rect 4972 1165 5018 1203
rect 4972 1131 4978 1165
rect 5012 1131 5018 1165
rect 4972 1093 5018 1131
rect 4972 1059 4978 1093
rect 5012 1059 5018 1093
rect 4972 1021 5018 1059
rect 4972 987 4978 1021
rect 5012 987 5018 1021
rect 4972 949 5018 987
rect 4972 915 4978 949
rect 5012 915 5018 949
rect 4972 877 5018 915
rect 4972 843 4978 877
rect 5012 843 5018 877
rect 4972 805 5018 843
rect 4972 771 4978 805
rect 5012 771 5018 805
rect 4972 733 5018 771
rect 4972 699 4978 733
rect 5012 699 5018 733
rect 4972 661 5018 699
rect 4972 627 4978 661
rect 5012 627 5018 661
rect 4972 589 5018 627
rect 4972 555 4978 589
rect 5012 555 5018 589
rect 4972 517 5018 555
rect 4972 483 4978 517
rect 5012 483 5018 517
rect 4972 445 5018 483
rect 4972 411 4978 445
rect 5012 411 5018 445
rect 4972 373 5018 411
rect 4972 339 4978 373
rect 5012 339 5018 373
rect 4972 301 5018 339
rect 4972 267 4978 301
rect 5012 267 5018 301
rect 4972 252 5018 267
rect 5068 1237 5114 1252
rect 5068 1203 5074 1237
rect 5108 1203 5114 1237
rect 5068 1165 5114 1203
rect 5068 1131 5074 1165
rect 5108 1131 5114 1165
rect 5068 1093 5114 1131
rect 5068 1059 5074 1093
rect 5108 1059 5114 1093
rect 5068 1021 5114 1059
rect 5068 987 5074 1021
rect 5108 987 5114 1021
rect 5068 949 5114 987
rect 5068 915 5074 949
rect 5108 915 5114 949
rect 5068 877 5114 915
rect 5068 843 5074 877
rect 5108 843 5114 877
rect 5068 805 5114 843
rect 5068 771 5074 805
rect 5108 771 5114 805
rect 5068 733 5114 771
rect 5068 699 5074 733
rect 5108 699 5114 733
rect 5068 661 5114 699
rect 5068 627 5074 661
rect 5108 627 5114 661
rect 5068 589 5114 627
rect 5068 555 5074 589
rect 5108 555 5114 589
rect 5068 517 5114 555
rect 5068 483 5074 517
rect 5108 483 5114 517
rect 5068 445 5114 483
rect 5068 411 5074 445
rect 5108 411 5114 445
rect 5068 373 5114 411
rect 5068 339 5074 373
rect 5108 339 5114 373
rect 5068 301 5114 339
rect 5068 267 5074 301
rect 5108 267 5114 301
rect 5068 252 5114 267
rect 5164 1237 5210 1252
rect 5164 1203 5170 1237
rect 5204 1203 5210 1237
rect 5164 1165 5210 1203
rect 5164 1131 5170 1165
rect 5204 1131 5210 1165
rect 5164 1093 5210 1131
rect 5164 1059 5170 1093
rect 5204 1059 5210 1093
rect 5164 1021 5210 1059
rect 5164 987 5170 1021
rect 5204 987 5210 1021
rect 5164 949 5210 987
rect 5164 915 5170 949
rect 5204 915 5210 949
rect 5164 877 5210 915
rect 5164 843 5170 877
rect 5204 843 5210 877
rect 5164 805 5210 843
rect 5164 771 5170 805
rect 5204 771 5210 805
rect 5164 733 5210 771
rect 5164 699 5170 733
rect 5204 699 5210 733
rect 5164 661 5210 699
rect 5164 627 5170 661
rect 5204 627 5210 661
rect 5164 589 5210 627
rect 5164 555 5170 589
rect 5204 555 5210 589
rect 5164 517 5210 555
rect 5164 483 5170 517
rect 5204 483 5210 517
rect 5164 445 5210 483
rect 5164 411 5170 445
rect 5204 411 5210 445
rect 5164 373 5210 411
rect 5164 339 5170 373
rect 5204 339 5210 373
rect 5164 301 5210 339
rect 5164 267 5170 301
rect 5204 267 5210 301
rect 5164 252 5210 267
rect 5260 1237 5306 1252
rect 5260 1203 5266 1237
rect 5300 1203 5306 1237
rect 5260 1165 5306 1203
rect 5260 1131 5266 1165
rect 5300 1131 5306 1165
rect 5260 1093 5306 1131
rect 5260 1059 5266 1093
rect 5300 1059 5306 1093
rect 5260 1021 5306 1059
rect 5260 987 5266 1021
rect 5300 987 5306 1021
rect 5260 949 5306 987
rect 5260 915 5266 949
rect 5300 915 5306 949
rect 5260 877 5306 915
rect 5260 843 5266 877
rect 5300 843 5306 877
rect 5260 805 5306 843
rect 5260 771 5266 805
rect 5300 771 5306 805
rect 5260 733 5306 771
rect 5260 699 5266 733
rect 5300 699 5306 733
rect 5260 661 5306 699
rect 5260 627 5266 661
rect 5300 627 5306 661
rect 5260 589 5306 627
rect 5260 555 5266 589
rect 5300 555 5306 589
rect 5260 517 5306 555
rect 5260 483 5266 517
rect 5300 483 5306 517
rect 5260 445 5306 483
rect 5260 411 5266 445
rect 5300 411 5306 445
rect 5260 373 5306 411
rect 5260 339 5266 373
rect 5300 339 5306 373
rect 5260 301 5306 339
rect 5260 267 5266 301
rect 5300 267 5306 301
rect 5260 252 5306 267
rect 5356 1237 5402 1252
rect 5356 1203 5362 1237
rect 5396 1203 5402 1237
rect 5356 1165 5402 1203
rect 5356 1131 5362 1165
rect 5396 1131 5402 1165
rect 5356 1093 5402 1131
rect 5356 1059 5362 1093
rect 5396 1059 5402 1093
rect 5356 1021 5402 1059
rect 5356 987 5362 1021
rect 5396 987 5402 1021
rect 5356 949 5402 987
rect 5356 915 5362 949
rect 5396 915 5402 949
rect 5356 877 5402 915
rect 5356 843 5362 877
rect 5396 843 5402 877
rect 5356 805 5402 843
rect 5356 771 5362 805
rect 5396 771 5402 805
rect 5356 733 5402 771
rect 5356 699 5362 733
rect 5396 699 5402 733
rect 5356 661 5402 699
rect 5356 627 5362 661
rect 5396 627 5402 661
rect 5356 589 5402 627
rect 5356 555 5362 589
rect 5396 555 5402 589
rect 5356 517 5402 555
rect 5356 483 5362 517
rect 5396 483 5402 517
rect 5356 445 5402 483
rect 5356 411 5362 445
rect 5396 411 5402 445
rect 5356 373 5402 411
rect 5356 339 5362 373
rect 5396 339 5402 373
rect 5356 301 5402 339
rect 5356 267 5362 301
rect 5396 267 5402 301
rect 5356 252 5402 267
rect 5452 1237 5498 1252
rect 5452 1203 5458 1237
rect 5492 1203 5498 1237
rect 5452 1165 5498 1203
rect 5452 1131 5458 1165
rect 5492 1131 5498 1165
rect 5452 1093 5498 1131
rect 5452 1059 5458 1093
rect 5492 1059 5498 1093
rect 5452 1021 5498 1059
rect 5452 987 5458 1021
rect 5492 987 5498 1021
rect 5452 949 5498 987
rect 5452 915 5458 949
rect 5492 915 5498 949
rect 5452 877 5498 915
rect 5452 843 5458 877
rect 5492 843 5498 877
rect 5452 805 5498 843
rect 5452 771 5458 805
rect 5492 771 5498 805
rect 5452 733 5498 771
rect 5452 699 5458 733
rect 5492 699 5498 733
rect 5452 661 5498 699
rect 5452 627 5458 661
rect 5492 627 5498 661
rect 5452 589 5498 627
rect 5452 555 5458 589
rect 5492 555 5498 589
rect 5452 517 5498 555
rect 5452 483 5458 517
rect 5492 483 5498 517
rect 5452 445 5498 483
rect 5452 411 5458 445
rect 5492 411 5498 445
rect 5452 373 5498 411
rect 5452 339 5458 373
rect 5492 339 5498 373
rect 5452 301 5498 339
rect 5452 267 5458 301
rect 5492 267 5498 301
rect 5452 252 5498 267
rect 5548 1237 5594 1252
rect 5548 1203 5554 1237
rect 5588 1203 5594 1237
rect 5548 1165 5594 1203
rect 5548 1131 5554 1165
rect 5588 1131 5594 1165
rect 5548 1093 5594 1131
rect 5548 1059 5554 1093
rect 5588 1059 5594 1093
rect 5548 1021 5594 1059
rect 5548 987 5554 1021
rect 5588 987 5594 1021
rect 5548 949 5594 987
rect 5548 915 5554 949
rect 5588 915 5594 949
rect 5548 877 5594 915
rect 5548 843 5554 877
rect 5588 843 5594 877
rect 5548 805 5594 843
rect 5548 771 5554 805
rect 5588 771 5594 805
rect 5548 733 5594 771
rect 5548 699 5554 733
rect 5588 699 5594 733
rect 5548 661 5594 699
rect 5548 627 5554 661
rect 5588 627 5594 661
rect 5548 589 5594 627
rect 5548 555 5554 589
rect 5588 555 5594 589
rect 5548 517 5594 555
rect 5548 483 5554 517
rect 5588 483 5594 517
rect 5548 445 5594 483
rect 5548 411 5554 445
rect 5588 411 5594 445
rect 5548 373 5594 411
rect 5548 339 5554 373
rect 5588 339 5594 373
rect 5548 301 5594 339
rect 5548 267 5554 301
rect 5588 267 5594 301
rect 5548 252 5594 267
rect 5644 1237 5690 1252
rect 5644 1203 5650 1237
rect 5684 1203 5690 1237
rect 5644 1165 5690 1203
rect 5644 1131 5650 1165
rect 5684 1131 5690 1165
rect 5644 1093 5690 1131
rect 5644 1059 5650 1093
rect 5684 1059 5690 1093
rect 5644 1021 5690 1059
rect 5644 987 5650 1021
rect 5684 987 5690 1021
rect 5644 949 5690 987
rect 5644 915 5650 949
rect 5684 915 5690 949
rect 5644 877 5690 915
rect 5644 843 5650 877
rect 5684 843 5690 877
rect 5644 805 5690 843
rect 5644 771 5650 805
rect 5684 771 5690 805
rect 5644 733 5690 771
rect 5644 699 5650 733
rect 5684 699 5690 733
rect 5644 661 5690 699
rect 5644 627 5650 661
rect 5684 627 5690 661
rect 5644 589 5690 627
rect 5644 555 5650 589
rect 5684 555 5690 589
rect 5644 517 5690 555
rect 5644 483 5650 517
rect 5684 483 5690 517
rect 5644 445 5690 483
rect 5644 411 5650 445
rect 5684 411 5690 445
rect 5644 373 5690 411
rect 5644 339 5650 373
rect 5684 339 5690 373
rect 5644 301 5690 339
rect 5644 267 5650 301
rect 5684 267 5690 301
rect 5644 252 5690 267
rect 5740 1237 5786 1252
rect 5740 1203 5746 1237
rect 5780 1203 5786 1237
rect 5740 1165 5786 1203
rect 5740 1131 5746 1165
rect 5780 1131 5786 1165
rect 5740 1093 5786 1131
rect 5740 1059 5746 1093
rect 5780 1059 5786 1093
rect 5740 1021 5786 1059
rect 5740 987 5746 1021
rect 5780 987 5786 1021
rect 5740 949 5786 987
rect 5740 915 5746 949
rect 5780 915 5786 949
rect 5740 877 5786 915
rect 5740 843 5746 877
rect 5780 843 5786 877
rect 5740 805 5786 843
rect 5740 771 5746 805
rect 5780 771 5786 805
rect 5740 733 5786 771
rect 5740 699 5746 733
rect 5780 699 5786 733
rect 5740 661 5786 699
rect 5740 627 5746 661
rect 5780 627 5786 661
rect 5740 589 5786 627
rect 5740 555 5746 589
rect 5780 555 5786 589
rect 5740 517 5786 555
rect 5740 483 5746 517
rect 5780 483 5786 517
rect 5740 445 5786 483
rect 5740 411 5746 445
rect 5780 411 5786 445
rect 5740 373 5786 411
rect 5740 339 5746 373
rect 5780 339 5786 373
rect 5740 301 5786 339
rect 5740 267 5746 301
rect 5780 267 5786 301
rect 5740 252 5786 267
rect 5836 1237 5882 1252
rect 5836 1203 5842 1237
rect 5876 1203 5882 1237
rect 5836 1165 5882 1203
rect 5836 1131 5842 1165
rect 5876 1131 5882 1165
rect 5836 1093 5882 1131
rect 5836 1059 5842 1093
rect 5876 1059 5882 1093
rect 5836 1021 5882 1059
rect 5836 987 5842 1021
rect 5876 987 5882 1021
rect 5836 949 5882 987
rect 5836 915 5842 949
rect 5876 915 5882 949
rect 5836 877 5882 915
rect 5836 843 5842 877
rect 5876 843 5882 877
rect 5836 805 5882 843
rect 5836 771 5842 805
rect 5876 771 5882 805
rect 5836 733 5882 771
rect 5836 699 5842 733
rect 5876 699 5882 733
rect 5836 661 5882 699
rect 5836 627 5842 661
rect 5876 627 5882 661
rect 5836 589 5882 627
rect 5836 555 5842 589
rect 5876 555 5882 589
rect 5836 517 5882 555
rect 5836 483 5842 517
rect 5876 483 5882 517
rect 5836 445 5882 483
rect 5836 411 5842 445
rect 5876 411 5882 445
rect 5836 373 5882 411
rect 5836 339 5842 373
rect 5876 339 5882 373
rect 5836 301 5882 339
rect 5836 267 5842 301
rect 5876 267 5882 301
rect 5836 252 5882 267
rect 5932 1237 5978 1252
rect 5932 1203 5938 1237
rect 5972 1203 5978 1237
rect 5932 1165 5978 1203
rect 5932 1131 5938 1165
rect 5972 1131 5978 1165
rect 5932 1093 5978 1131
rect 5932 1059 5938 1093
rect 5972 1059 5978 1093
rect 5932 1021 5978 1059
rect 5932 987 5938 1021
rect 5972 987 5978 1021
rect 5932 949 5978 987
rect 5932 915 5938 949
rect 5972 915 5978 949
rect 5932 877 5978 915
rect 5932 843 5938 877
rect 5972 843 5978 877
rect 5932 805 5978 843
rect 5932 771 5938 805
rect 5972 771 5978 805
rect 5932 733 5978 771
rect 5932 699 5938 733
rect 5972 699 5978 733
rect 5932 661 5978 699
rect 5932 627 5938 661
rect 5972 627 5978 661
rect 5932 589 5978 627
rect 5932 555 5938 589
rect 5972 555 5978 589
rect 5932 517 5978 555
rect 5932 483 5938 517
rect 5972 483 5978 517
rect 5932 445 5978 483
rect 5932 411 5938 445
rect 5972 411 5978 445
rect 5932 373 5978 411
rect 5932 339 5938 373
rect 5972 339 5978 373
rect 5932 301 5978 339
rect 5932 267 5938 301
rect 5972 267 5978 301
rect 5932 252 5978 267
rect 6138 1237 6184 1252
rect 6138 1203 6144 1237
rect 6178 1203 6184 1237
rect 6138 1165 6184 1203
rect 6138 1131 6144 1165
rect 6178 1131 6184 1165
rect 6138 1093 6184 1131
rect 6138 1059 6144 1093
rect 6178 1059 6184 1093
rect 6138 1021 6184 1059
rect 6138 987 6144 1021
rect 6178 987 6184 1021
rect 6138 949 6184 987
rect 6138 915 6144 949
rect 6178 915 6184 949
rect 6138 877 6184 915
rect 6138 843 6144 877
rect 6178 843 6184 877
rect 6138 805 6184 843
rect 6138 771 6144 805
rect 6178 771 6184 805
rect 6138 733 6184 771
rect 6138 699 6144 733
rect 6178 699 6184 733
rect 6138 661 6184 699
rect 6138 627 6144 661
rect 6178 627 6184 661
rect 6138 589 6184 627
rect 6138 555 6144 589
rect 6178 555 6184 589
rect 6138 517 6184 555
rect 6138 483 6144 517
rect 6178 483 6184 517
rect 6138 445 6184 483
rect 6138 411 6144 445
rect 6178 411 6184 445
rect 6138 373 6184 411
rect 6138 339 6144 373
rect 6178 339 6184 373
rect 6138 301 6184 339
rect 6138 267 6144 301
rect 6178 267 6184 301
rect 6138 252 6184 267
rect 6234 1237 6280 1252
rect 6234 1203 6240 1237
rect 6274 1203 6280 1237
rect 6234 1165 6280 1203
rect 6234 1131 6240 1165
rect 6274 1131 6280 1165
rect 6234 1093 6280 1131
rect 6234 1059 6240 1093
rect 6274 1059 6280 1093
rect 6234 1021 6280 1059
rect 6234 987 6240 1021
rect 6274 987 6280 1021
rect 6234 949 6280 987
rect 6234 915 6240 949
rect 6274 915 6280 949
rect 6234 877 6280 915
rect 6234 843 6240 877
rect 6274 843 6280 877
rect 6234 805 6280 843
rect 6234 771 6240 805
rect 6274 771 6280 805
rect 6234 733 6280 771
rect 6234 699 6240 733
rect 6274 699 6280 733
rect 6234 661 6280 699
rect 6234 627 6240 661
rect 6274 627 6280 661
rect 6234 589 6280 627
rect 6234 555 6240 589
rect 6274 555 6280 589
rect 6234 517 6280 555
rect 6234 483 6240 517
rect 6274 483 6280 517
rect 6234 445 6280 483
rect 6234 411 6240 445
rect 6274 411 6280 445
rect 6234 373 6280 411
rect 6234 339 6240 373
rect 6274 339 6280 373
rect 6234 301 6280 339
rect 6234 267 6240 301
rect 6274 267 6280 301
rect 6234 252 6280 267
rect 6330 1237 6376 1252
rect 6330 1203 6336 1237
rect 6370 1203 6376 1237
rect 6330 1165 6376 1203
rect 6330 1131 6336 1165
rect 6370 1131 6376 1165
rect 6330 1093 6376 1131
rect 6330 1059 6336 1093
rect 6370 1059 6376 1093
rect 6330 1021 6376 1059
rect 6330 987 6336 1021
rect 6370 987 6376 1021
rect 6330 949 6376 987
rect 6330 915 6336 949
rect 6370 915 6376 949
rect 6330 877 6376 915
rect 6330 843 6336 877
rect 6370 843 6376 877
rect 6330 805 6376 843
rect 6330 771 6336 805
rect 6370 771 6376 805
rect 6330 733 6376 771
rect 6330 699 6336 733
rect 6370 699 6376 733
rect 6330 661 6376 699
rect 6330 627 6336 661
rect 6370 627 6376 661
rect 6330 589 6376 627
rect 6330 555 6336 589
rect 6370 555 6376 589
rect 6330 517 6376 555
rect 6330 483 6336 517
rect 6370 483 6376 517
rect 6330 445 6376 483
rect 6330 411 6336 445
rect 6370 411 6376 445
rect 6330 373 6376 411
rect 6330 339 6336 373
rect 6370 339 6376 373
rect 6330 301 6376 339
rect 6330 267 6336 301
rect 6370 267 6376 301
rect 6330 252 6376 267
rect 6426 1237 6472 1252
rect 6426 1203 6432 1237
rect 6466 1203 6472 1237
rect 6426 1165 6472 1203
rect 6426 1131 6432 1165
rect 6466 1131 6472 1165
rect 6426 1093 6472 1131
rect 6426 1059 6432 1093
rect 6466 1059 6472 1093
rect 6426 1021 6472 1059
rect 6426 987 6432 1021
rect 6466 987 6472 1021
rect 6426 949 6472 987
rect 6426 915 6432 949
rect 6466 915 6472 949
rect 6426 877 6472 915
rect 6426 843 6432 877
rect 6466 843 6472 877
rect 6426 805 6472 843
rect 6426 771 6432 805
rect 6466 771 6472 805
rect 6426 733 6472 771
rect 6426 699 6432 733
rect 6466 699 6472 733
rect 6426 661 6472 699
rect 6426 627 6432 661
rect 6466 627 6472 661
rect 6426 589 6472 627
rect 6426 555 6432 589
rect 6466 555 6472 589
rect 6426 517 6472 555
rect 6426 483 6432 517
rect 6466 483 6472 517
rect 6426 445 6472 483
rect 6426 411 6432 445
rect 6466 411 6472 445
rect 6426 373 6472 411
rect 6426 339 6432 373
rect 6466 339 6472 373
rect 6426 301 6472 339
rect 6426 267 6432 301
rect 6466 267 6472 301
rect 6426 252 6472 267
rect 6522 1237 6568 1252
rect 6522 1203 6528 1237
rect 6562 1203 6568 1237
rect 6522 1165 6568 1203
rect 6522 1131 6528 1165
rect 6562 1131 6568 1165
rect 6522 1093 6568 1131
rect 6522 1059 6528 1093
rect 6562 1059 6568 1093
rect 6522 1021 6568 1059
rect 6522 987 6528 1021
rect 6562 987 6568 1021
rect 6522 949 6568 987
rect 6522 915 6528 949
rect 6562 915 6568 949
rect 6522 877 6568 915
rect 6522 843 6528 877
rect 6562 843 6568 877
rect 6522 805 6568 843
rect 6522 771 6528 805
rect 6562 771 6568 805
rect 6522 733 6568 771
rect 6522 699 6528 733
rect 6562 699 6568 733
rect 6522 661 6568 699
rect 6522 627 6528 661
rect 6562 627 6568 661
rect 6522 589 6568 627
rect 6522 555 6528 589
rect 6562 555 6568 589
rect 6522 517 6568 555
rect 6522 483 6528 517
rect 6562 483 6568 517
rect 6522 445 6568 483
rect 6522 411 6528 445
rect 6562 411 6568 445
rect 6522 373 6568 411
rect 6522 339 6528 373
rect 6562 339 6568 373
rect 6522 301 6568 339
rect 6522 267 6528 301
rect 6562 267 6568 301
rect 6522 252 6568 267
rect 6618 1237 6664 1252
rect 6618 1203 6624 1237
rect 6658 1203 6664 1237
rect 6618 1165 6664 1203
rect 6618 1131 6624 1165
rect 6658 1131 6664 1165
rect 6618 1093 6664 1131
rect 6618 1059 6624 1093
rect 6658 1059 6664 1093
rect 6618 1021 6664 1059
rect 6618 987 6624 1021
rect 6658 987 6664 1021
rect 6618 949 6664 987
rect 6618 915 6624 949
rect 6658 915 6664 949
rect 6618 877 6664 915
rect 6618 843 6624 877
rect 6658 843 6664 877
rect 6618 805 6664 843
rect 6618 771 6624 805
rect 6658 771 6664 805
rect 6618 733 6664 771
rect 6618 699 6624 733
rect 6658 699 6664 733
rect 6618 661 6664 699
rect 6618 627 6624 661
rect 6658 627 6664 661
rect 6618 589 6664 627
rect 6618 555 6624 589
rect 6658 555 6664 589
rect 6618 517 6664 555
rect 6618 483 6624 517
rect 6658 483 6664 517
rect 6618 445 6664 483
rect 6618 411 6624 445
rect 6658 411 6664 445
rect 6618 373 6664 411
rect 6618 339 6624 373
rect 6658 339 6664 373
rect 6618 301 6664 339
rect 6618 267 6624 301
rect 6658 267 6664 301
rect 6618 252 6664 267
rect 6714 1237 6760 1252
rect 6714 1203 6720 1237
rect 6754 1203 6760 1237
rect 6714 1165 6760 1203
rect 6714 1131 6720 1165
rect 6754 1131 6760 1165
rect 6714 1093 6760 1131
rect 6714 1059 6720 1093
rect 6754 1059 6760 1093
rect 6714 1021 6760 1059
rect 6714 987 6720 1021
rect 6754 987 6760 1021
rect 6714 949 6760 987
rect 6714 915 6720 949
rect 6754 915 6760 949
rect 6714 877 6760 915
rect 6714 843 6720 877
rect 6754 843 6760 877
rect 6714 805 6760 843
rect 6714 771 6720 805
rect 6754 771 6760 805
rect 6714 733 6760 771
rect 6714 699 6720 733
rect 6754 699 6760 733
rect 6714 661 6760 699
rect 6714 627 6720 661
rect 6754 627 6760 661
rect 6714 589 6760 627
rect 6714 555 6720 589
rect 6754 555 6760 589
rect 6714 517 6760 555
rect 6714 483 6720 517
rect 6754 483 6760 517
rect 6714 445 6760 483
rect 6714 411 6720 445
rect 6754 411 6760 445
rect 6714 373 6760 411
rect 6714 339 6720 373
rect 6754 339 6760 373
rect 6714 301 6760 339
rect 6714 267 6720 301
rect 6754 267 6760 301
rect 6714 252 6760 267
rect 6810 1237 6856 1252
rect 6810 1203 6816 1237
rect 6850 1203 6856 1237
rect 6810 1165 6856 1203
rect 6810 1131 6816 1165
rect 6850 1131 6856 1165
rect 6810 1093 6856 1131
rect 6810 1059 6816 1093
rect 6850 1059 6856 1093
rect 6810 1021 6856 1059
rect 6810 987 6816 1021
rect 6850 987 6856 1021
rect 6810 949 6856 987
rect 6810 915 6816 949
rect 6850 915 6856 949
rect 6810 877 6856 915
rect 6810 843 6816 877
rect 6850 843 6856 877
rect 6810 805 6856 843
rect 6810 771 6816 805
rect 6850 771 6856 805
rect 6810 733 6856 771
rect 6810 699 6816 733
rect 6850 699 6856 733
rect 6810 661 6856 699
rect 6810 627 6816 661
rect 6850 627 6856 661
rect 6810 589 6856 627
rect 6810 555 6816 589
rect 6850 555 6856 589
rect 6810 517 6856 555
rect 6810 483 6816 517
rect 6850 483 6856 517
rect 6810 445 6856 483
rect 6810 411 6816 445
rect 6850 411 6856 445
rect 6810 373 6856 411
rect 6810 339 6816 373
rect 6850 339 6856 373
rect 6810 301 6856 339
rect 6810 267 6816 301
rect 6850 267 6856 301
rect 6810 252 6856 267
rect 6906 1237 6952 1252
rect 6906 1203 6912 1237
rect 6946 1203 6952 1237
rect 6906 1165 6952 1203
rect 6906 1131 6912 1165
rect 6946 1131 6952 1165
rect 6906 1093 6952 1131
rect 6906 1059 6912 1093
rect 6946 1059 6952 1093
rect 6906 1021 6952 1059
rect 6906 987 6912 1021
rect 6946 987 6952 1021
rect 6906 949 6952 987
rect 6906 915 6912 949
rect 6946 915 6952 949
rect 6906 877 6952 915
rect 6906 843 6912 877
rect 6946 843 6952 877
rect 6906 805 6952 843
rect 6906 771 6912 805
rect 6946 771 6952 805
rect 6906 733 6952 771
rect 6906 699 6912 733
rect 6946 699 6952 733
rect 6906 661 6952 699
rect 6906 627 6912 661
rect 6946 627 6952 661
rect 6906 589 6952 627
rect 6906 555 6912 589
rect 6946 555 6952 589
rect 6906 517 6952 555
rect 6906 483 6912 517
rect 6946 483 6952 517
rect 6906 445 6952 483
rect 6906 411 6912 445
rect 6946 411 6952 445
rect 6906 373 6952 411
rect 6906 339 6912 373
rect 6946 339 6952 373
rect 6906 301 6952 339
rect 6906 267 6912 301
rect 6946 267 6952 301
rect 6906 252 6952 267
rect 7002 1237 7048 1252
rect 7002 1203 7008 1237
rect 7042 1203 7048 1237
rect 7002 1165 7048 1203
rect 7002 1131 7008 1165
rect 7042 1131 7048 1165
rect 7002 1093 7048 1131
rect 7002 1059 7008 1093
rect 7042 1059 7048 1093
rect 7002 1021 7048 1059
rect 7002 987 7008 1021
rect 7042 987 7048 1021
rect 7002 949 7048 987
rect 7002 915 7008 949
rect 7042 915 7048 949
rect 7002 877 7048 915
rect 7002 843 7008 877
rect 7042 843 7048 877
rect 7002 805 7048 843
rect 7002 771 7008 805
rect 7042 771 7048 805
rect 7002 733 7048 771
rect 7002 699 7008 733
rect 7042 699 7048 733
rect 7002 661 7048 699
rect 7002 627 7008 661
rect 7042 627 7048 661
rect 7002 589 7048 627
rect 7002 555 7008 589
rect 7042 555 7048 589
rect 7002 517 7048 555
rect 7002 483 7008 517
rect 7042 483 7048 517
rect 7002 445 7048 483
rect 7002 411 7008 445
rect 7042 411 7048 445
rect 7002 373 7048 411
rect 7002 339 7008 373
rect 7042 339 7048 373
rect 7002 301 7048 339
rect 7002 267 7008 301
rect 7042 267 7048 301
rect 7002 252 7048 267
rect 7098 1237 7144 1252
rect 7098 1203 7104 1237
rect 7138 1203 7144 1237
rect 7098 1165 7144 1203
rect 7098 1131 7104 1165
rect 7138 1131 7144 1165
rect 7098 1093 7144 1131
rect 7098 1059 7104 1093
rect 7138 1059 7144 1093
rect 7098 1021 7144 1059
rect 7098 987 7104 1021
rect 7138 987 7144 1021
rect 7098 949 7144 987
rect 7098 915 7104 949
rect 7138 915 7144 949
rect 7098 877 7144 915
rect 7098 843 7104 877
rect 7138 843 7144 877
rect 7098 805 7144 843
rect 7098 771 7104 805
rect 7138 771 7144 805
rect 7098 733 7144 771
rect 7098 699 7104 733
rect 7138 699 7144 733
rect 7098 661 7144 699
rect 7098 627 7104 661
rect 7138 627 7144 661
rect 7098 589 7144 627
rect 7098 555 7104 589
rect 7138 555 7144 589
rect 7098 517 7144 555
rect 7098 483 7104 517
rect 7138 483 7144 517
rect 7098 445 7144 483
rect 7098 411 7104 445
rect 7138 411 7144 445
rect 7098 373 7144 411
rect 7098 339 7104 373
rect 7138 339 7144 373
rect 7098 301 7144 339
rect 7098 267 7104 301
rect 7138 267 7144 301
rect 7098 252 7144 267
rect 7194 1237 7240 1252
rect 7194 1203 7200 1237
rect 7234 1203 7240 1237
rect 7194 1165 7240 1203
rect 7194 1131 7200 1165
rect 7234 1131 7240 1165
rect 7194 1093 7240 1131
rect 7194 1059 7200 1093
rect 7234 1059 7240 1093
rect 7194 1021 7240 1059
rect 7194 987 7200 1021
rect 7234 987 7240 1021
rect 7194 949 7240 987
rect 7194 915 7200 949
rect 7234 915 7240 949
rect 7194 877 7240 915
rect 7194 843 7200 877
rect 7234 843 7240 877
rect 7194 805 7240 843
rect 7194 771 7200 805
rect 7234 771 7240 805
rect 7194 733 7240 771
rect 7194 699 7200 733
rect 7234 699 7240 733
rect 7194 661 7240 699
rect 7194 627 7200 661
rect 7234 627 7240 661
rect 7194 589 7240 627
rect 7194 555 7200 589
rect 7234 555 7240 589
rect 7194 517 7240 555
rect 7194 483 7200 517
rect 7234 483 7240 517
rect 7194 445 7240 483
rect 7194 411 7200 445
rect 7234 411 7240 445
rect 7194 373 7240 411
rect 7194 339 7200 373
rect 7234 339 7240 373
rect 7194 301 7240 339
rect 7194 267 7200 301
rect 7234 267 7240 301
rect 7194 252 7240 267
rect 7290 1237 7336 1252
rect 7290 1203 7296 1237
rect 7330 1203 7336 1237
rect 7290 1165 7336 1203
rect 7290 1131 7296 1165
rect 7330 1131 7336 1165
rect 7290 1093 7336 1131
rect 7290 1059 7296 1093
rect 7330 1059 7336 1093
rect 7290 1021 7336 1059
rect 7290 987 7296 1021
rect 7330 987 7336 1021
rect 7290 949 7336 987
rect 7290 915 7296 949
rect 7330 915 7336 949
rect 7290 877 7336 915
rect 7290 843 7296 877
rect 7330 843 7336 877
rect 7290 805 7336 843
rect 7290 771 7296 805
rect 7330 771 7336 805
rect 7290 733 7336 771
rect 7290 699 7296 733
rect 7330 699 7336 733
rect 7290 661 7336 699
rect 7290 627 7296 661
rect 7330 627 7336 661
rect 7290 589 7336 627
rect 7290 555 7296 589
rect 7330 555 7336 589
rect 7290 517 7336 555
rect 7290 483 7296 517
rect 7330 483 7336 517
rect 7290 445 7336 483
rect 7290 411 7296 445
rect 7330 411 7336 445
rect 7290 373 7336 411
rect 7290 339 7296 373
rect 7330 339 7336 373
rect 7290 301 7336 339
rect 7290 267 7296 301
rect 7330 267 7336 301
rect 7290 252 7336 267
rect 7906 1237 7952 1252
rect 7906 1203 7912 1237
rect 7946 1203 7952 1237
rect 7906 1165 7952 1203
rect 7906 1131 7912 1165
rect 7946 1131 7952 1165
rect 7906 1093 7952 1131
rect 7906 1059 7912 1093
rect 7946 1059 7952 1093
rect 7906 1021 7952 1059
rect 7906 987 7912 1021
rect 7946 987 7952 1021
rect 7906 949 7952 987
rect 7906 915 7912 949
rect 7946 915 7952 949
rect 7906 877 7952 915
rect 7906 843 7912 877
rect 7946 843 7952 877
rect 7906 805 7952 843
rect 7906 771 7912 805
rect 7946 771 7952 805
rect 7906 733 7952 771
rect 7906 699 7912 733
rect 7946 699 7952 733
rect 7906 661 7952 699
rect 7906 627 7912 661
rect 7946 627 7952 661
rect 7906 589 7952 627
rect 7906 555 7912 589
rect 7946 555 7952 589
rect 7906 517 7952 555
rect 7906 483 7912 517
rect 7946 483 7952 517
rect 7906 445 7952 483
rect 7906 411 7912 445
rect 7946 411 7952 445
rect 7906 373 7952 411
rect 7906 339 7912 373
rect 7946 339 7952 373
rect 7906 301 7952 339
rect 7906 267 7912 301
rect 7946 267 7952 301
rect 7906 252 7952 267
rect 8002 1237 8048 1252
rect 8002 1203 8008 1237
rect 8042 1203 8048 1237
rect 8002 1165 8048 1203
rect 8002 1131 8008 1165
rect 8042 1131 8048 1165
rect 8002 1093 8048 1131
rect 8002 1059 8008 1093
rect 8042 1059 8048 1093
rect 8002 1021 8048 1059
rect 8002 987 8008 1021
rect 8042 987 8048 1021
rect 8002 949 8048 987
rect 8002 915 8008 949
rect 8042 915 8048 949
rect 8002 877 8048 915
rect 8002 843 8008 877
rect 8042 843 8048 877
rect 8002 805 8048 843
rect 8002 771 8008 805
rect 8042 771 8048 805
rect 8002 733 8048 771
rect 8002 699 8008 733
rect 8042 699 8048 733
rect 8002 661 8048 699
rect 8002 627 8008 661
rect 8042 627 8048 661
rect 8002 589 8048 627
rect 8002 555 8008 589
rect 8042 555 8048 589
rect 8002 517 8048 555
rect 8002 483 8008 517
rect 8042 483 8048 517
rect 8002 445 8048 483
rect 8002 411 8008 445
rect 8042 411 8048 445
rect 8002 373 8048 411
rect 8002 339 8008 373
rect 8042 339 8048 373
rect 8002 301 8048 339
rect 8002 267 8008 301
rect 8042 267 8048 301
rect 8002 252 8048 267
rect 8098 1237 8144 1252
rect 8098 1203 8104 1237
rect 8138 1203 8144 1237
rect 8098 1165 8144 1203
rect 8098 1131 8104 1165
rect 8138 1131 8144 1165
rect 8098 1093 8144 1131
rect 8098 1059 8104 1093
rect 8138 1059 8144 1093
rect 8098 1021 8144 1059
rect 8098 987 8104 1021
rect 8138 987 8144 1021
rect 8098 949 8144 987
rect 8098 915 8104 949
rect 8138 915 8144 949
rect 8098 877 8144 915
rect 8098 843 8104 877
rect 8138 843 8144 877
rect 8098 805 8144 843
rect 8098 771 8104 805
rect 8138 771 8144 805
rect 8098 733 8144 771
rect 8098 699 8104 733
rect 8138 699 8144 733
rect 8098 661 8144 699
rect 8098 627 8104 661
rect 8138 627 8144 661
rect 8098 589 8144 627
rect 8098 555 8104 589
rect 8138 555 8144 589
rect 8098 517 8144 555
rect 8098 483 8104 517
rect 8138 483 8144 517
rect 8098 445 8144 483
rect 8098 411 8104 445
rect 8138 411 8144 445
rect 8098 373 8144 411
rect 8098 339 8104 373
rect 8138 339 8144 373
rect 8098 301 8144 339
rect 8098 267 8104 301
rect 8138 267 8144 301
rect 8098 252 8144 267
rect 8194 1237 8240 1252
rect 8194 1203 8200 1237
rect 8234 1203 8240 1237
rect 8194 1165 8240 1203
rect 8194 1131 8200 1165
rect 8234 1131 8240 1165
rect 8194 1093 8240 1131
rect 8194 1059 8200 1093
rect 8234 1059 8240 1093
rect 8194 1021 8240 1059
rect 8194 987 8200 1021
rect 8234 987 8240 1021
rect 8194 949 8240 987
rect 8194 915 8200 949
rect 8234 915 8240 949
rect 8194 877 8240 915
rect 8194 843 8200 877
rect 8234 843 8240 877
rect 8194 805 8240 843
rect 8194 771 8200 805
rect 8234 771 8240 805
rect 8194 733 8240 771
rect 8194 699 8200 733
rect 8234 699 8240 733
rect 8194 661 8240 699
rect 8194 627 8200 661
rect 8234 627 8240 661
rect 8194 589 8240 627
rect 8194 555 8200 589
rect 8234 555 8240 589
rect 8194 517 8240 555
rect 8194 483 8200 517
rect 8234 483 8240 517
rect 8194 445 8240 483
rect 8194 411 8200 445
rect 8234 411 8240 445
rect 8194 373 8240 411
rect 8194 339 8200 373
rect 8234 339 8240 373
rect 8194 301 8240 339
rect 8194 267 8200 301
rect 8234 267 8240 301
rect 8194 252 8240 267
rect 8290 1237 8336 1252
rect 8290 1203 8296 1237
rect 8330 1203 8336 1237
rect 8290 1165 8336 1203
rect 8290 1131 8296 1165
rect 8330 1131 8336 1165
rect 8290 1093 8336 1131
rect 8290 1059 8296 1093
rect 8330 1059 8336 1093
rect 8290 1021 8336 1059
rect 8290 987 8296 1021
rect 8330 987 8336 1021
rect 8290 949 8336 987
rect 8290 915 8296 949
rect 8330 915 8336 949
rect 8290 877 8336 915
rect 8290 843 8296 877
rect 8330 843 8336 877
rect 8290 805 8336 843
rect 8290 771 8296 805
rect 8330 771 8336 805
rect 8290 733 8336 771
rect 8290 699 8296 733
rect 8330 699 8336 733
rect 8290 661 8336 699
rect 8290 627 8296 661
rect 8330 627 8336 661
rect 8290 589 8336 627
rect 8290 555 8296 589
rect 8330 555 8336 589
rect 8290 517 8336 555
rect 8290 483 8296 517
rect 8330 483 8336 517
rect 8290 445 8336 483
rect 8290 411 8296 445
rect 8330 411 8336 445
rect 8290 373 8336 411
rect 8290 339 8296 373
rect 8330 339 8336 373
rect 8290 301 8336 339
rect 8290 267 8296 301
rect 8330 267 8336 301
rect 8290 252 8336 267
rect 8386 1237 8432 1252
rect 8386 1203 8392 1237
rect 8426 1203 8432 1237
rect 8386 1165 8432 1203
rect 8386 1131 8392 1165
rect 8426 1131 8432 1165
rect 8386 1093 8432 1131
rect 8386 1059 8392 1093
rect 8426 1059 8432 1093
rect 8386 1021 8432 1059
rect 8386 987 8392 1021
rect 8426 987 8432 1021
rect 8386 949 8432 987
rect 8386 915 8392 949
rect 8426 915 8432 949
rect 8386 877 8432 915
rect 8386 843 8392 877
rect 8426 843 8432 877
rect 8386 805 8432 843
rect 8386 771 8392 805
rect 8426 771 8432 805
rect 8386 733 8432 771
rect 8386 699 8392 733
rect 8426 699 8432 733
rect 8386 661 8432 699
rect 8386 627 8392 661
rect 8426 627 8432 661
rect 8386 589 8432 627
rect 8386 555 8392 589
rect 8426 555 8432 589
rect 8386 517 8432 555
rect 8386 483 8392 517
rect 8426 483 8432 517
rect 8386 445 8432 483
rect 8386 411 8392 445
rect 8426 411 8432 445
rect 8386 373 8432 411
rect 8386 339 8392 373
rect 8426 339 8432 373
rect 8386 301 8432 339
rect 8386 267 8392 301
rect 8426 267 8432 301
rect 8386 252 8432 267
rect 8482 1237 8528 1252
rect 8482 1203 8488 1237
rect 8522 1203 8528 1237
rect 8482 1165 8528 1203
rect 8482 1131 8488 1165
rect 8522 1131 8528 1165
rect 8482 1093 8528 1131
rect 8482 1059 8488 1093
rect 8522 1059 8528 1093
rect 8482 1021 8528 1059
rect 8482 987 8488 1021
rect 8522 987 8528 1021
rect 8482 949 8528 987
rect 8482 915 8488 949
rect 8522 915 8528 949
rect 8482 877 8528 915
rect 8482 843 8488 877
rect 8522 843 8528 877
rect 8482 805 8528 843
rect 8482 771 8488 805
rect 8522 771 8528 805
rect 8482 733 8528 771
rect 8482 699 8488 733
rect 8522 699 8528 733
rect 8482 661 8528 699
rect 8482 627 8488 661
rect 8522 627 8528 661
rect 8482 589 8528 627
rect 8482 555 8488 589
rect 8522 555 8528 589
rect 8482 517 8528 555
rect 8482 483 8488 517
rect 8522 483 8528 517
rect 8482 445 8528 483
rect 8482 411 8488 445
rect 8522 411 8528 445
rect 8482 373 8528 411
rect 8482 339 8488 373
rect 8522 339 8528 373
rect 8482 301 8528 339
rect 8482 267 8488 301
rect 8522 267 8528 301
rect 8482 252 8528 267
rect 8578 1237 8624 1252
rect 8578 1203 8584 1237
rect 8618 1203 8624 1237
rect 8578 1165 8624 1203
rect 8578 1131 8584 1165
rect 8618 1131 8624 1165
rect 8578 1093 8624 1131
rect 8578 1059 8584 1093
rect 8618 1059 8624 1093
rect 8578 1021 8624 1059
rect 8578 987 8584 1021
rect 8618 987 8624 1021
rect 8578 949 8624 987
rect 8578 915 8584 949
rect 8618 915 8624 949
rect 8578 877 8624 915
rect 8578 843 8584 877
rect 8618 843 8624 877
rect 8578 805 8624 843
rect 8578 771 8584 805
rect 8618 771 8624 805
rect 8578 733 8624 771
rect 8578 699 8584 733
rect 8618 699 8624 733
rect 8578 661 8624 699
rect 8578 627 8584 661
rect 8618 627 8624 661
rect 8578 589 8624 627
rect 8578 555 8584 589
rect 8618 555 8624 589
rect 8578 517 8624 555
rect 8578 483 8584 517
rect 8618 483 8624 517
rect 8578 445 8624 483
rect 8578 411 8584 445
rect 8618 411 8624 445
rect 8578 373 8624 411
rect 8578 339 8584 373
rect 8618 339 8624 373
rect 8578 301 8624 339
rect 8578 267 8584 301
rect 8618 267 8624 301
rect 8578 252 8624 267
rect 8674 1237 8720 1252
rect 8674 1203 8680 1237
rect 8714 1203 8720 1237
rect 8674 1165 8720 1203
rect 8674 1131 8680 1165
rect 8714 1131 8720 1165
rect 8674 1093 8720 1131
rect 8674 1059 8680 1093
rect 8714 1059 8720 1093
rect 8674 1021 8720 1059
rect 8674 987 8680 1021
rect 8714 987 8720 1021
rect 8674 949 8720 987
rect 8674 915 8680 949
rect 8714 915 8720 949
rect 8674 877 8720 915
rect 8674 843 8680 877
rect 8714 843 8720 877
rect 8674 805 8720 843
rect 8674 771 8680 805
rect 8714 771 8720 805
rect 8674 733 8720 771
rect 8674 699 8680 733
rect 8714 699 8720 733
rect 8674 661 8720 699
rect 8674 627 8680 661
rect 8714 627 8720 661
rect 8674 589 8720 627
rect 8674 555 8680 589
rect 8714 555 8720 589
rect 8674 517 8720 555
rect 8674 483 8680 517
rect 8714 483 8720 517
rect 8674 445 8720 483
rect 8674 411 8680 445
rect 8714 411 8720 445
rect 8674 373 8720 411
rect 8674 339 8680 373
rect 8714 339 8720 373
rect 8674 301 8720 339
rect 8674 267 8680 301
rect 8714 267 8720 301
rect 8674 252 8720 267
rect 8770 1237 8816 1252
rect 8770 1203 8776 1237
rect 8810 1203 8816 1237
rect 8770 1165 8816 1203
rect 8770 1131 8776 1165
rect 8810 1131 8816 1165
rect 8770 1093 8816 1131
rect 8770 1059 8776 1093
rect 8810 1059 8816 1093
rect 8770 1021 8816 1059
rect 8770 987 8776 1021
rect 8810 987 8816 1021
rect 8770 949 8816 987
rect 8770 915 8776 949
rect 8810 915 8816 949
rect 8770 877 8816 915
rect 8770 843 8776 877
rect 8810 843 8816 877
rect 8770 805 8816 843
rect 8770 771 8776 805
rect 8810 771 8816 805
rect 8770 733 8816 771
rect 8770 699 8776 733
rect 8810 699 8816 733
rect 8770 661 8816 699
rect 8770 627 8776 661
rect 8810 627 8816 661
rect 8770 589 8816 627
rect 8770 555 8776 589
rect 8810 555 8816 589
rect 8770 517 8816 555
rect 8770 483 8776 517
rect 8810 483 8816 517
rect 8770 445 8816 483
rect 8770 411 8776 445
rect 8810 411 8816 445
rect 8770 373 8816 411
rect 8770 339 8776 373
rect 8810 339 8816 373
rect 8770 301 8816 339
rect 8770 267 8776 301
rect 8810 267 8816 301
rect 8770 252 8816 267
rect 8866 1237 8912 1252
rect 8866 1203 8872 1237
rect 8906 1203 8912 1237
rect 8866 1165 8912 1203
rect 8866 1131 8872 1165
rect 8906 1131 8912 1165
rect 8866 1093 8912 1131
rect 8866 1059 8872 1093
rect 8906 1059 8912 1093
rect 8866 1021 8912 1059
rect 8866 987 8872 1021
rect 8906 987 8912 1021
rect 8866 949 8912 987
rect 8866 915 8872 949
rect 8906 915 8912 949
rect 8866 877 8912 915
rect 8866 843 8872 877
rect 8906 843 8912 877
rect 8866 805 8912 843
rect 8866 771 8872 805
rect 8906 771 8912 805
rect 8866 733 8912 771
rect 8866 699 8872 733
rect 8906 699 8912 733
rect 8866 661 8912 699
rect 8866 627 8872 661
rect 8906 627 8912 661
rect 8866 589 8912 627
rect 8866 555 8872 589
rect 8906 555 8912 589
rect 8866 517 8912 555
rect 8866 483 8872 517
rect 8906 483 8912 517
rect 8866 445 8912 483
rect 8866 411 8872 445
rect 8906 411 8912 445
rect 8866 373 8912 411
rect 8866 339 8872 373
rect 8906 339 8912 373
rect 8866 301 8912 339
rect 8866 267 8872 301
rect 8906 267 8912 301
rect 8866 252 8912 267
rect 8962 1237 9008 1252
rect 8962 1203 8968 1237
rect 9002 1203 9008 1237
rect 8962 1165 9008 1203
rect 8962 1131 8968 1165
rect 9002 1131 9008 1165
rect 8962 1093 9008 1131
rect 8962 1059 8968 1093
rect 9002 1059 9008 1093
rect 8962 1021 9008 1059
rect 8962 987 8968 1021
rect 9002 987 9008 1021
rect 8962 949 9008 987
rect 8962 915 8968 949
rect 9002 915 9008 949
rect 8962 877 9008 915
rect 8962 843 8968 877
rect 9002 843 9008 877
rect 8962 805 9008 843
rect 8962 771 8968 805
rect 9002 771 9008 805
rect 8962 733 9008 771
rect 8962 699 8968 733
rect 9002 699 9008 733
rect 8962 661 9008 699
rect 8962 627 8968 661
rect 9002 627 9008 661
rect 8962 589 9008 627
rect 8962 555 8968 589
rect 9002 555 9008 589
rect 8962 517 9008 555
rect 8962 483 8968 517
rect 9002 483 9008 517
rect 8962 445 9008 483
rect 8962 411 8968 445
rect 9002 411 9008 445
rect 8962 373 9008 411
rect 8962 339 8968 373
rect 9002 339 9008 373
rect 8962 301 9008 339
rect 8962 267 8968 301
rect 9002 267 9008 301
rect 8962 252 9008 267
rect 9226 1235 9272 1250
rect 9226 1201 9232 1235
rect 9266 1201 9272 1235
rect 9226 1163 9272 1201
rect 9226 1129 9232 1163
rect 9266 1129 9272 1163
rect 9226 1091 9272 1129
rect 9226 1057 9232 1091
rect 9266 1057 9272 1091
rect 9226 1019 9272 1057
rect 9226 985 9232 1019
rect 9266 985 9272 1019
rect 9226 947 9272 985
rect 9226 913 9232 947
rect 9266 913 9272 947
rect 9226 875 9272 913
rect 9226 841 9232 875
rect 9266 841 9272 875
rect 9226 803 9272 841
rect 9226 769 9232 803
rect 9266 769 9272 803
rect 9226 731 9272 769
rect 9226 697 9232 731
rect 9266 697 9272 731
rect 9226 659 9272 697
rect 9226 625 9232 659
rect 9266 625 9272 659
rect 9226 587 9272 625
rect 9226 553 9232 587
rect 9266 553 9272 587
rect 9226 515 9272 553
rect 9226 481 9232 515
rect 9266 481 9272 515
rect 9226 443 9272 481
rect 9226 409 9232 443
rect 9266 409 9272 443
rect 9226 371 9272 409
rect 9226 337 9232 371
rect 9266 337 9272 371
rect 9226 299 9272 337
rect 9226 265 9232 299
rect 9266 265 9272 299
rect 9226 250 9272 265
rect 9322 1235 9368 1250
rect 9322 1201 9328 1235
rect 9362 1201 9368 1235
rect 9322 1163 9368 1201
rect 9322 1129 9328 1163
rect 9362 1129 9368 1163
rect 9322 1091 9368 1129
rect 9322 1057 9328 1091
rect 9362 1057 9368 1091
rect 9322 1019 9368 1057
rect 9322 985 9328 1019
rect 9362 985 9368 1019
rect 9322 947 9368 985
rect 9322 913 9328 947
rect 9362 913 9368 947
rect 9322 875 9368 913
rect 9322 841 9328 875
rect 9362 841 9368 875
rect 9322 803 9368 841
rect 9322 769 9328 803
rect 9362 769 9368 803
rect 9322 731 9368 769
rect 9322 697 9328 731
rect 9362 697 9368 731
rect 9322 659 9368 697
rect 9322 625 9328 659
rect 9362 625 9368 659
rect 9322 587 9368 625
rect 9322 553 9328 587
rect 9362 553 9368 587
rect 9322 515 9368 553
rect 9322 481 9328 515
rect 9362 481 9368 515
rect 9322 443 9368 481
rect 9322 409 9328 443
rect 9362 409 9368 443
rect 9322 371 9368 409
rect 9322 337 9328 371
rect 9362 337 9368 371
rect 9322 299 9368 337
rect 9322 265 9328 299
rect 9362 265 9368 299
rect 9322 250 9368 265
rect 9418 1235 9464 1250
rect 9418 1201 9424 1235
rect 9458 1201 9464 1235
rect 9418 1163 9464 1201
rect 9418 1129 9424 1163
rect 9458 1129 9464 1163
rect 9418 1091 9464 1129
rect 9418 1057 9424 1091
rect 9458 1057 9464 1091
rect 9418 1019 9464 1057
rect 9418 985 9424 1019
rect 9458 985 9464 1019
rect 9418 947 9464 985
rect 9418 913 9424 947
rect 9458 913 9464 947
rect 9418 875 9464 913
rect 9418 841 9424 875
rect 9458 841 9464 875
rect 9418 803 9464 841
rect 9418 769 9424 803
rect 9458 769 9464 803
rect 9418 731 9464 769
rect 9418 697 9424 731
rect 9458 697 9464 731
rect 9418 659 9464 697
rect 9418 625 9424 659
rect 9458 625 9464 659
rect 9418 587 9464 625
rect 9418 553 9424 587
rect 9458 553 9464 587
rect 9418 515 9464 553
rect 9418 481 9424 515
rect 9458 481 9464 515
rect 9418 443 9464 481
rect 9418 409 9424 443
rect 9458 409 9464 443
rect 9418 371 9464 409
rect 9418 337 9424 371
rect 9458 337 9464 371
rect 9418 299 9464 337
rect 9418 265 9424 299
rect 9458 265 9464 299
rect 9418 250 9464 265
rect 9514 1235 9560 1250
rect 9514 1201 9520 1235
rect 9554 1201 9560 1235
rect 9514 1163 9560 1201
rect 9514 1129 9520 1163
rect 9554 1129 9560 1163
rect 9514 1091 9560 1129
rect 9514 1057 9520 1091
rect 9554 1057 9560 1091
rect 9514 1019 9560 1057
rect 9514 985 9520 1019
rect 9554 985 9560 1019
rect 9514 947 9560 985
rect 9514 913 9520 947
rect 9554 913 9560 947
rect 9514 875 9560 913
rect 9514 841 9520 875
rect 9554 841 9560 875
rect 9514 803 9560 841
rect 9514 769 9520 803
rect 9554 769 9560 803
rect 9514 731 9560 769
rect 9514 697 9520 731
rect 9554 697 9560 731
rect 9514 659 9560 697
rect 9514 625 9520 659
rect 9554 625 9560 659
rect 9514 587 9560 625
rect 9514 553 9520 587
rect 9554 553 9560 587
rect 9514 515 9560 553
rect 9514 481 9520 515
rect 9554 481 9560 515
rect 9514 443 9560 481
rect 9514 409 9520 443
rect 9554 409 9560 443
rect 9514 371 9560 409
rect 9514 337 9520 371
rect 9554 337 9560 371
rect 9514 299 9560 337
rect 9514 265 9520 299
rect 9554 265 9560 299
rect 9514 250 9560 265
rect 9610 1235 9656 1250
rect 9610 1201 9616 1235
rect 9650 1201 9656 1235
rect 9610 1163 9656 1201
rect 9610 1129 9616 1163
rect 9650 1129 9656 1163
rect 9610 1091 9656 1129
rect 9610 1057 9616 1091
rect 9650 1057 9656 1091
rect 9610 1019 9656 1057
rect 9610 985 9616 1019
rect 9650 985 9656 1019
rect 9610 947 9656 985
rect 9610 913 9616 947
rect 9650 913 9656 947
rect 9610 875 9656 913
rect 9610 841 9616 875
rect 9650 841 9656 875
rect 9610 803 9656 841
rect 9610 769 9616 803
rect 9650 769 9656 803
rect 9610 731 9656 769
rect 9610 697 9616 731
rect 9650 697 9656 731
rect 9610 659 9656 697
rect 9610 625 9616 659
rect 9650 625 9656 659
rect 9610 587 9656 625
rect 9610 553 9616 587
rect 9650 553 9656 587
rect 9610 515 9656 553
rect 9610 481 9616 515
rect 9650 481 9656 515
rect 9610 443 9656 481
rect 9610 409 9616 443
rect 9650 409 9656 443
rect 9610 371 9656 409
rect 9610 337 9616 371
rect 9650 337 9656 371
rect 9610 299 9656 337
rect 9610 265 9616 299
rect 9650 265 9656 299
rect 9610 250 9656 265
rect 9706 1235 9752 1250
rect 9706 1201 9712 1235
rect 9746 1201 9752 1235
rect 9706 1163 9752 1201
rect 9706 1129 9712 1163
rect 9746 1129 9752 1163
rect 9706 1091 9752 1129
rect 9706 1057 9712 1091
rect 9746 1057 9752 1091
rect 9706 1019 9752 1057
rect 9706 985 9712 1019
rect 9746 985 9752 1019
rect 9706 947 9752 985
rect 9706 913 9712 947
rect 9746 913 9752 947
rect 9706 875 9752 913
rect 9706 841 9712 875
rect 9746 841 9752 875
rect 9706 803 9752 841
rect 9706 769 9712 803
rect 9746 769 9752 803
rect 9706 731 9752 769
rect 9706 697 9712 731
rect 9746 697 9752 731
rect 9706 659 9752 697
rect 9706 625 9712 659
rect 9746 625 9752 659
rect 9706 587 9752 625
rect 9706 553 9712 587
rect 9746 553 9752 587
rect 9706 515 9752 553
rect 9706 481 9712 515
rect 9746 481 9752 515
rect 9706 443 9752 481
rect 9706 409 9712 443
rect 9746 409 9752 443
rect 9706 371 9752 409
rect 9706 337 9712 371
rect 9746 337 9752 371
rect 9706 299 9752 337
rect 9706 265 9712 299
rect 9746 265 9752 299
rect 9706 250 9752 265
rect 9802 1235 9848 1250
rect 9802 1201 9808 1235
rect 9842 1201 9848 1235
rect 9802 1163 9848 1201
rect 9802 1129 9808 1163
rect 9842 1129 9848 1163
rect 9802 1091 9848 1129
rect 9802 1057 9808 1091
rect 9842 1057 9848 1091
rect 9802 1019 9848 1057
rect 9802 985 9808 1019
rect 9842 985 9848 1019
rect 9802 947 9848 985
rect 9802 913 9808 947
rect 9842 913 9848 947
rect 9802 875 9848 913
rect 9802 841 9808 875
rect 9842 841 9848 875
rect 9802 803 9848 841
rect 9802 769 9808 803
rect 9842 769 9848 803
rect 9802 731 9848 769
rect 9802 697 9808 731
rect 9842 697 9848 731
rect 9802 659 9848 697
rect 9802 625 9808 659
rect 9842 625 9848 659
rect 9802 587 9848 625
rect 9802 553 9808 587
rect 9842 553 9848 587
rect 9802 515 9848 553
rect 9802 481 9808 515
rect 9842 481 9848 515
rect 9802 443 9848 481
rect 9802 409 9808 443
rect 9842 409 9848 443
rect 9802 371 9848 409
rect 9802 337 9808 371
rect 9842 337 9848 371
rect 9802 299 9848 337
rect 9802 265 9808 299
rect 9842 265 9848 299
rect 9802 250 9848 265
rect 9898 1235 9944 1250
rect 9898 1201 9904 1235
rect 9938 1201 9944 1235
rect 9898 1163 9944 1201
rect 9898 1129 9904 1163
rect 9938 1129 9944 1163
rect 9898 1091 9944 1129
rect 9898 1057 9904 1091
rect 9938 1057 9944 1091
rect 9898 1019 9944 1057
rect 9898 985 9904 1019
rect 9938 985 9944 1019
rect 9898 947 9944 985
rect 9898 913 9904 947
rect 9938 913 9944 947
rect 9898 875 9944 913
rect 9898 841 9904 875
rect 9938 841 9944 875
rect 9898 803 9944 841
rect 9898 769 9904 803
rect 9938 769 9944 803
rect 9898 731 9944 769
rect 9898 697 9904 731
rect 9938 697 9944 731
rect 9898 659 9944 697
rect 9898 625 9904 659
rect 9938 625 9944 659
rect 9898 587 9944 625
rect 9898 553 9904 587
rect 9938 553 9944 587
rect 9898 515 9944 553
rect 9898 481 9904 515
rect 9938 481 9944 515
rect 9898 443 9944 481
rect 9898 409 9904 443
rect 9938 409 9944 443
rect 9898 371 9944 409
rect 9898 337 9904 371
rect 9938 337 9944 371
rect 9898 299 9944 337
rect 9898 265 9904 299
rect 9938 265 9944 299
rect 9898 250 9944 265
rect 9994 1235 10040 1250
rect 9994 1201 10000 1235
rect 10034 1201 10040 1235
rect 9994 1163 10040 1201
rect 9994 1129 10000 1163
rect 10034 1129 10040 1163
rect 9994 1091 10040 1129
rect 9994 1057 10000 1091
rect 10034 1057 10040 1091
rect 9994 1019 10040 1057
rect 9994 985 10000 1019
rect 10034 985 10040 1019
rect 9994 947 10040 985
rect 9994 913 10000 947
rect 10034 913 10040 947
rect 9994 875 10040 913
rect 9994 841 10000 875
rect 10034 841 10040 875
rect 9994 803 10040 841
rect 9994 769 10000 803
rect 10034 769 10040 803
rect 9994 731 10040 769
rect 9994 697 10000 731
rect 10034 697 10040 731
rect 9994 659 10040 697
rect 9994 625 10000 659
rect 10034 625 10040 659
rect 9994 587 10040 625
rect 9994 553 10000 587
rect 10034 553 10040 587
rect 9994 515 10040 553
rect 9994 481 10000 515
rect 10034 481 10040 515
rect 9994 443 10040 481
rect 9994 409 10000 443
rect 10034 409 10040 443
rect 9994 371 10040 409
rect 9994 337 10000 371
rect 10034 337 10040 371
rect 9994 299 10040 337
rect 9994 265 10000 299
rect 10034 265 10040 299
rect 9994 250 10040 265
rect 10090 1235 10136 1250
rect 10090 1201 10096 1235
rect 10130 1201 10136 1235
rect 10090 1163 10136 1201
rect 10090 1129 10096 1163
rect 10130 1129 10136 1163
rect 10090 1091 10136 1129
rect 10090 1057 10096 1091
rect 10130 1057 10136 1091
rect 10090 1019 10136 1057
rect 10090 985 10096 1019
rect 10130 985 10136 1019
rect 10090 947 10136 985
rect 10090 913 10096 947
rect 10130 913 10136 947
rect 10090 875 10136 913
rect 10090 841 10096 875
rect 10130 841 10136 875
rect 10090 803 10136 841
rect 10090 769 10096 803
rect 10130 769 10136 803
rect 10090 731 10136 769
rect 10090 697 10096 731
rect 10130 697 10136 731
rect 10090 659 10136 697
rect 10090 625 10096 659
rect 10130 625 10136 659
rect 10090 587 10136 625
rect 10090 553 10096 587
rect 10130 553 10136 587
rect 10090 515 10136 553
rect 10090 481 10096 515
rect 10130 481 10136 515
rect 10090 443 10136 481
rect 10090 409 10096 443
rect 10130 409 10136 443
rect 10090 371 10136 409
rect 10090 337 10096 371
rect 10130 337 10136 371
rect 10090 299 10136 337
rect 10090 265 10096 299
rect 10130 265 10136 299
rect 10090 250 10136 265
rect 10186 1235 10232 1250
rect 10186 1201 10192 1235
rect 10226 1201 10232 1235
rect 10186 1163 10232 1201
rect 10186 1129 10192 1163
rect 10226 1129 10232 1163
rect 10186 1091 10232 1129
rect 10186 1057 10192 1091
rect 10226 1057 10232 1091
rect 10186 1019 10232 1057
rect 10186 985 10192 1019
rect 10226 985 10232 1019
rect 10186 947 10232 985
rect 10186 913 10192 947
rect 10226 913 10232 947
rect 10186 875 10232 913
rect 10186 841 10192 875
rect 10226 841 10232 875
rect 10186 803 10232 841
rect 10186 769 10192 803
rect 10226 769 10232 803
rect 10186 731 10232 769
rect 10186 697 10192 731
rect 10226 697 10232 731
rect 10186 659 10232 697
rect 10186 625 10192 659
rect 10226 625 10232 659
rect 10186 587 10232 625
rect 10186 553 10192 587
rect 10226 553 10232 587
rect 10186 515 10232 553
rect 10186 481 10192 515
rect 10226 481 10232 515
rect 10186 443 10232 481
rect 10186 409 10192 443
rect 10226 409 10232 443
rect 10186 371 10232 409
rect 10186 337 10192 371
rect 10226 337 10232 371
rect 10186 299 10232 337
rect 10186 265 10192 299
rect 10226 265 10232 299
rect 10186 250 10232 265
rect 10282 1235 10328 1250
rect 10282 1201 10288 1235
rect 10322 1201 10328 1235
rect 10282 1163 10328 1201
rect 10282 1129 10288 1163
rect 10322 1129 10328 1163
rect 10282 1091 10328 1129
rect 10282 1057 10288 1091
rect 10322 1057 10328 1091
rect 10282 1019 10328 1057
rect 10282 985 10288 1019
rect 10322 985 10328 1019
rect 10282 947 10328 985
rect 10282 913 10288 947
rect 10322 913 10328 947
rect 10282 875 10328 913
rect 10282 841 10288 875
rect 10322 841 10328 875
rect 10282 803 10328 841
rect 10282 769 10288 803
rect 10322 769 10328 803
rect 10282 731 10328 769
rect 10282 697 10288 731
rect 10322 697 10328 731
rect 10282 659 10328 697
rect 10282 625 10288 659
rect 10322 625 10328 659
rect 10282 587 10328 625
rect 10282 553 10288 587
rect 10322 553 10328 587
rect 10282 515 10328 553
rect 10282 481 10288 515
rect 10322 481 10328 515
rect 10282 443 10328 481
rect 10282 409 10288 443
rect 10322 409 10328 443
rect 10282 371 10328 409
rect 10282 337 10288 371
rect 10322 337 10328 371
rect 10282 299 10328 337
rect 10282 265 10288 299
rect 10322 265 10328 299
rect 10282 250 10328 265
rect 10378 1235 10424 1250
rect 10378 1201 10384 1235
rect 10418 1201 10424 1235
rect 10378 1163 10424 1201
rect 10378 1129 10384 1163
rect 10418 1129 10424 1163
rect 10378 1091 10424 1129
rect 10378 1057 10384 1091
rect 10418 1057 10424 1091
rect 10378 1019 10424 1057
rect 10378 985 10384 1019
rect 10418 985 10424 1019
rect 10378 947 10424 985
rect 10378 913 10384 947
rect 10418 913 10424 947
rect 10378 875 10424 913
rect 10378 841 10384 875
rect 10418 841 10424 875
rect 10378 803 10424 841
rect 10378 769 10384 803
rect 10418 769 10424 803
rect 10378 731 10424 769
rect 10378 697 10384 731
rect 10418 697 10424 731
rect 10378 659 10424 697
rect 10378 625 10384 659
rect 10418 625 10424 659
rect 10378 587 10424 625
rect 10378 553 10384 587
rect 10418 553 10424 587
rect 10378 515 10424 553
rect 10378 481 10384 515
rect 10418 481 10424 515
rect 10378 443 10424 481
rect 10378 409 10384 443
rect 10418 409 10424 443
rect 10378 371 10424 409
rect 10378 337 10384 371
rect 10418 337 10424 371
rect 10378 299 10424 337
rect 10378 265 10384 299
rect 10418 265 10424 299
rect 10378 250 10424 265
rect 10994 1235 11040 1250
rect 10994 1201 11000 1235
rect 11034 1201 11040 1235
rect 10994 1163 11040 1201
rect 10994 1129 11000 1163
rect 11034 1129 11040 1163
rect 10994 1091 11040 1129
rect 10994 1057 11000 1091
rect 11034 1057 11040 1091
rect 10994 1019 11040 1057
rect 10994 985 11000 1019
rect 11034 985 11040 1019
rect 10994 947 11040 985
rect 10994 913 11000 947
rect 11034 913 11040 947
rect 10994 875 11040 913
rect 10994 841 11000 875
rect 11034 841 11040 875
rect 10994 803 11040 841
rect 10994 769 11000 803
rect 11034 769 11040 803
rect 10994 731 11040 769
rect 10994 697 11000 731
rect 11034 697 11040 731
rect 10994 659 11040 697
rect 10994 625 11000 659
rect 11034 625 11040 659
rect 10994 587 11040 625
rect 10994 553 11000 587
rect 11034 553 11040 587
rect 10994 515 11040 553
rect 10994 481 11000 515
rect 11034 481 11040 515
rect 10994 443 11040 481
rect 10994 409 11000 443
rect 11034 409 11040 443
rect 10994 371 11040 409
rect 10994 337 11000 371
rect 11034 337 11040 371
rect 10994 299 11040 337
rect 10994 265 11000 299
rect 11034 265 11040 299
rect 10994 250 11040 265
rect 11090 1235 11136 1250
rect 11090 1201 11096 1235
rect 11130 1201 11136 1235
rect 11090 1163 11136 1201
rect 11090 1129 11096 1163
rect 11130 1129 11136 1163
rect 11090 1091 11136 1129
rect 11090 1057 11096 1091
rect 11130 1057 11136 1091
rect 11090 1019 11136 1057
rect 11090 985 11096 1019
rect 11130 985 11136 1019
rect 11090 947 11136 985
rect 11090 913 11096 947
rect 11130 913 11136 947
rect 11090 875 11136 913
rect 11090 841 11096 875
rect 11130 841 11136 875
rect 11090 803 11136 841
rect 11090 769 11096 803
rect 11130 769 11136 803
rect 11090 731 11136 769
rect 11090 697 11096 731
rect 11130 697 11136 731
rect 11090 659 11136 697
rect 11090 625 11096 659
rect 11130 625 11136 659
rect 11090 587 11136 625
rect 11090 553 11096 587
rect 11130 553 11136 587
rect 11090 515 11136 553
rect 11090 481 11096 515
rect 11130 481 11136 515
rect 11090 443 11136 481
rect 11090 409 11096 443
rect 11130 409 11136 443
rect 11090 371 11136 409
rect 11090 337 11096 371
rect 11130 337 11136 371
rect 11090 299 11136 337
rect 11090 265 11096 299
rect 11130 265 11136 299
rect 11090 250 11136 265
rect 11186 1235 11232 1250
rect 11186 1201 11192 1235
rect 11226 1201 11232 1235
rect 11186 1163 11232 1201
rect 11186 1129 11192 1163
rect 11226 1129 11232 1163
rect 11186 1091 11232 1129
rect 11186 1057 11192 1091
rect 11226 1057 11232 1091
rect 11186 1019 11232 1057
rect 11186 985 11192 1019
rect 11226 985 11232 1019
rect 11186 947 11232 985
rect 11186 913 11192 947
rect 11226 913 11232 947
rect 11186 875 11232 913
rect 11186 841 11192 875
rect 11226 841 11232 875
rect 11186 803 11232 841
rect 11186 769 11192 803
rect 11226 769 11232 803
rect 11186 731 11232 769
rect 11186 697 11192 731
rect 11226 697 11232 731
rect 11186 659 11232 697
rect 11186 625 11192 659
rect 11226 625 11232 659
rect 11186 587 11232 625
rect 11186 553 11192 587
rect 11226 553 11232 587
rect 11186 515 11232 553
rect 11186 481 11192 515
rect 11226 481 11232 515
rect 11186 443 11232 481
rect 11186 409 11192 443
rect 11226 409 11232 443
rect 11186 371 11232 409
rect 11186 337 11192 371
rect 11226 337 11232 371
rect 11186 299 11232 337
rect 11186 265 11192 299
rect 11226 265 11232 299
rect 11186 250 11232 265
rect 11282 1235 11328 1250
rect 11282 1201 11288 1235
rect 11322 1201 11328 1235
rect 11282 1163 11328 1201
rect 11282 1129 11288 1163
rect 11322 1129 11328 1163
rect 11282 1091 11328 1129
rect 11282 1057 11288 1091
rect 11322 1057 11328 1091
rect 11282 1019 11328 1057
rect 11282 985 11288 1019
rect 11322 985 11328 1019
rect 11282 947 11328 985
rect 11282 913 11288 947
rect 11322 913 11328 947
rect 11282 875 11328 913
rect 11282 841 11288 875
rect 11322 841 11328 875
rect 11282 803 11328 841
rect 11282 769 11288 803
rect 11322 769 11328 803
rect 11282 731 11328 769
rect 11282 697 11288 731
rect 11322 697 11328 731
rect 11282 659 11328 697
rect 11282 625 11288 659
rect 11322 625 11328 659
rect 11282 587 11328 625
rect 11282 553 11288 587
rect 11322 553 11328 587
rect 11282 515 11328 553
rect 11282 481 11288 515
rect 11322 481 11328 515
rect 11282 443 11328 481
rect 11282 409 11288 443
rect 11322 409 11328 443
rect 11282 371 11328 409
rect 11282 337 11288 371
rect 11322 337 11328 371
rect 11282 299 11328 337
rect 11282 265 11288 299
rect 11322 265 11328 299
rect 11282 250 11328 265
rect 11378 1235 11424 1250
rect 11378 1201 11384 1235
rect 11418 1201 11424 1235
rect 11378 1163 11424 1201
rect 11378 1129 11384 1163
rect 11418 1129 11424 1163
rect 11378 1091 11424 1129
rect 11378 1057 11384 1091
rect 11418 1057 11424 1091
rect 11378 1019 11424 1057
rect 11378 985 11384 1019
rect 11418 985 11424 1019
rect 11378 947 11424 985
rect 11378 913 11384 947
rect 11418 913 11424 947
rect 11378 875 11424 913
rect 11378 841 11384 875
rect 11418 841 11424 875
rect 11378 803 11424 841
rect 11378 769 11384 803
rect 11418 769 11424 803
rect 11378 731 11424 769
rect 11378 697 11384 731
rect 11418 697 11424 731
rect 11378 659 11424 697
rect 11378 625 11384 659
rect 11418 625 11424 659
rect 11378 587 11424 625
rect 11378 553 11384 587
rect 11418 553 11424 587
rect 11378 515 11424 553
rect 11378 481 11384 515
rect 11418 481 11424 515
rect 11378 443 11424 481
rect 11378 409 11384 443
rect 11418 409 11424 443
rect 11378 371 11424 409
rect 11378 337 11384 371
rect 11418 337 11424 371
rect 11378 299 11424 337
rect 11378 265 11384 299
rect 11418 265 11424 299
rect 11378 250 11424 265
rect 11474 1235 11520 1250
rect 11474 1201 11480 1235
rect 11514 1201 11520 1235
rect 11474 1163 11520 1201
rect 11474 1129 11480 1163
rect 11514 1129 11520 1163
rect 11474 1091 11520 1129
rect 11474 1057 11480 1091
rect 11514 1057 11520 1091
rect 11474 1019 11520 1057
rect 11474 985 11480 1019
rect 11514 985 11520 1019
rect 11474 947 11520 985
rect 11474 913 11480 947
rect 11514 913 11520 947
rect 11474 875 11520 913
rect 11474 841 11480 875
rect 11514 841 11520 875
rect 11474 803 11520 841
rect 11474 769 11480 803
rect 11514 769 11520 803
rect 11474 731 11520 769
rect 11474 697 11480 731
rect 11514 697 11520 731
rect 11474 659 11520 697
rect 11474 625 11480 659
rect 11514 625 11520 659
rect 11474 587 11520 625
rect 11474 553 11480 587
rect 11514 553 11520 587
rect 11474 515 11520 553
rect 11474 481 11480 515
rect 11514 481 11520 515
rect 11474 443 11520 481
rect 11474 409 11480 443
rect 11514 409 11520 443
rect 11474 371 11520 409
rect 11474 337 11480 371
rect 11514 337 11520 371
rect 11474 299 11520 337
rect 11474 265 11480 299
rect 11514 265 11520 299
rect 11474 250 11520 265
rect 11570 1235 11616 1250
rect 11570 1201 11576 1235
rect 11610 1201 11616 1235
rect 11570 1163 11616 1201
rect 11570 1129 11576 1163
rect 11610 1129 11616 1163
rect 11570 1091 11616 1129
rect 11570 1057 11576 1091
rect 11610 1057 11616 1091
rect 11570 1019 11616 1057
rect 11570 985 11576 1019
rect 11610 985 11616 1019
rect 11570 947 11616 985
rect 11570 913 11576 947
rect 11610 913 11616 947
rect 11570 875 11616 913
rect 11570 841 11576 875
rect 11610 841 11616 875
rect 11570 803 11616 841
rect 11570 769 11576 803
rect 11610 769 11616 803
rect 11570 731 11616 769
rect 11570 697 11576 731
rect 11610 697 11616 731
rect 11570 659 11616 697
rect 11570 625 11576 659
rect 11610 625 11616 659
rect 11570 587 11616 625
rect 11570 553 11576 587
rect 11610 553 11616 587
rect 11570 515 11616 553
rect 11570 481 11576 515
rect 11610 481 11616 515
rect 11570 443 11616 481
rect 11570 409 11576 443
rect 11610 409 11616 443
rect 11570 371 11616 409
rect 11570 337 11576 371
rect 11610 337 11616 371
rect 11570 299 11616 337
rect 11570 265 11576 299
rect 11610 265 11616 299
rect 11570 250 11616 265
rect 11666 1235 11712 1250
rect 11666 1201 11672 1235
rect 11706 1201 11712 1235
rect 11666 1163 11712 1201
rect 11666 1129 11672 1163
rect 11706 1129 11712 1163
rect 11666 1091 11712 1129
rect 11666 1057 11672 1091
rect 11706 1057 11712 1091
rect 11666 1019 11712 1057
rect 11666 985 11672 1019
rect 11706 985 11712 1019
rect 11666 947 11712 985
rect 11666 913 11672 947
rect 11706 913 11712 947
rect 11666 875 11712 913
rect 11666 841 11672 875
rect 11706 841 11712 875
rect 11666 803 11712 841
rect 11666 769 11672 803
rect 11706 769 11712 803
rect 11666 731 11712 769
rect 11666 697 11672 731
rect 11706 697 11712 731
rect 11666 659 11712 697
rect 11666 625 11672 659
rect 11706 625 11712 659
rect 11666 587 11712 625
rect 11666 553 11672 587
rect 11706 553 11712 587
rect 11666 515 11712 553
rect 11666 481 11672 515
rect 11706 481 11712 515
rect 11666 443 11712 481
rect 11666 409 11672 443
rect 11706 409 11712 443
rect 11666 371 11712 409
rect 11666 337 11672 371
rect 11706 337 11712 371
rect 11666 299 11712 337
rect 11666 265 11672 299
rect 11706 265 11712 299
rect 11666 250 11712 265
rect 11762 1235 11808 1250
rect 11762 1201 11768 1235
rect 11802 1201 11808 1235
rect 11762 1163 11808 1201
rect 11762 1129 11768 1163
rect 11802 1129 11808 1163
rect 11762 1091 11808 1129
rect 11762 1057 11768 1091
rect 11802 1057 11808 1091
rect 11762 1019 11808 1057
rect 11762 985 11768 1019
rect 11802 985 11808 1019
rect 11762 947 11808 985
rect 11762 913 11768 947
rect 11802 913 11808 947
rect 11762 875 11808 913
rect 11762 841 11768 875
rect 11802 841 11808 875
rect 11762 803 11808 841
rect 11762 769 11768 803
rect 11802 769 11808 803
rect 11762 731 11808 769
rect 11762 697 11768 731
rect 11802 697 11808 731
rect 11762 659 11808 697
rect 11762 625 11768 659
rect 11802 625 11808 659
rect 11762 587 11808 625
rect 11762 553 11768 587
rect 11802 553 11808 587
rect 11762 515 11808 553
rect 11762 481 11768 515
rect 11802 481 11808 515
rect 11762 443 11808 481
rect 11762 409 11768 443
rect 11802 409 11808 443
rect 11762 371 11808 409
rect 11762 337 11768 371
rect 11802 337 11808 371
rect 11762 299 11808 337
rect 11762 265 11768 299
rect 11802 265 11808 299
rect 11762 250 11808 265
rect 11858 1235 11904 1250
rect 11858 1201 11864 1235
rect 11898 1201 11904 1235
rect 11858 1163 11904 1201
rect 11858 1129 11864 1163
rect 11898 1129 11904 1163
rect 11858 1091 11904 1129
rect 11858 1057 11864 1091
rect 11898 1057 11904 1091
rect 11858 1019 11904 1057
rect 11858 985 11864 1019
rect 11898 985 11904 1019
rect 11858 947 11904 985
rect 11858 913 11864 947
rect 11898 913 11904 947
rect 11858 875 11904 913
rect 11858 841 11864 875
rect 11898 841 11904 875
rect 11858 803 11904 841
rect 11858 769 11864 803
rect 11898 769 11904 803
rect 11858 731 11904 769
rect 11858 697 11864 731
rect 11898 697 11904 731
rect 11858 659 11904 697
rect 11858 625 11864 659
rect 11898 625 11904 659
rect 11858 587 11904 625
rect 11858 553 11864 587
rect 11898 553 11904 587
rect 11858 515 11904 553
rect 11858 481 11864 515
rect 11898 481 11904 515
rect 11858 443 11904 481
rect 11858 409 11864 443
rect 11898 409 11904 443
rect 11858 371 11904 409
rect 11858 337 11864 371
rect 11898 337 11904 371
rect 11858 299 11904 337
rect 11858 265 11864 299
rect 11898 265 11904 299
rect 11858 250 11904 265
rect 11954 1235 12000 1250
rect 11954 1201 11960 1235
rect 11994 1201 12000 1235
rect 11954 1163 12000 1201
rect 11954 1129 11960 1163
rect 11994 1129 12000 1163
rect 11954 1091 12000 1129
rect 11954 1057 11960 1091
rect 11994 1057 12000 1091
rect 11954 1019 12000 1057
rect 11954 985 11960 1019
rect 11994 985 12000 1019
rect 11954 947 12000 985
rect 11954 913 11960 947
rect 11994 913 12000 947
rect 11954 875 12000 913
rect 11954 841 11960 875
rect 11994 841 12000 875
rect 11954 803 12000 841
rect 11954 769 11960 803
rect 11994 769 12000 803
rect 11954 731 12000 769
rect 11954 697 11960 731
rect 11994 697 12000 731
rect 11954 659 12000 697
rect 11954 625 11960 659
rect 11994 625 12000 659
rect 11954 587 12000 625
rect 11954 553 11960 587
rect 11994 553 12000 587
rect 11954 515 12000 553
rect 11954 481 11960 515
rect 11994 481 12000 515
rect 11954 443 12000 481
rect 11954 409 11960 443
rect 11994 409 12000 443
rect 11954 371 12000 409
rect 11954 337 11960 371
rect 11994 337 12000 371
rect 11954 299 12000 337
rect 11954 265 11960 299
rect 11994 265 12000 299
rect 11954 250 12000 265
rect 12050 1235 12096 1250
rect 12050 1201 12056 1235
rect 12090 1201 12096 1235
rect 12050 1163 12096 1201
rect 12050 1129 12056 1163
rect 12090 1129 12096 1163
rect 12050 1091 12096 1129
rect 12050 1057 12056 1091
rect 12090 1057 12096 1091
rect 12050 1019 12096 1057
rect 12050 985 12056 1019
rect 12090 985 12096 1019
rect 12050 947 12096 985
rect 12050 913 12056 947
rect 12090 913 12096 947
rect 12050 875 12096 913
rect 12050 841 12056 875
rect 12090 841 12096 875
rect 12050 803 12096 841
rect 12050 769 12056 803
rect 12090 769 12096 803
rect 12050 731 12096 769
rect 12050 697 12056 731
rect 12090 697 12096 731
rect 12050 659 12096 697
rect 12050 625 12056 659
rect 12090 625 12096 659
rect 12050 587 12096 625
rect 12050 553 12056 587
rect 12090 553 12096 587
rect 12050 515 12096 553
rect 12050 481 12056 515
rect 12090 481 12096 515
rect 12050 443 12096 481
rect 12050 409 12056 443
rect 12090 409 12096 443
rect 12050 371 12096 409
rect 12050 337 12056 371
rect 12090 337 12096 371
rect 12050 299 12096 337
rect 12050 265 12056 299
rect 12090 265 12096 299
rect 12050 250 12096 265
rect 12382 1209 12428 1224
rect 12382 1175 12388 1209
rect 12422 1175 12428 1209
rect 12382 1137 12428 1175
rect 12382 1103 12388 1137
rect 12422 1103 12428 1137
rect 12382 1065 12428 1103
rect 12382 1031 12388 1065
rect 12422 1031 12428 1065
rect 12382 993 12428 1031
rect 12382 959 12388 993
rect 12422 959 12428 993
rect 12382 921 12428 959
rect 12382 887 12388 921
rect 12422 887 12428 921
rect 12382 849 12428 887
rect 12382 815 12388 849
rect 12422 815 12428 849
rect 12382 777 12428 815
rect 12382 743 12388 777
rect 12422 743 12428 777
rect 12382 705 12428 743
rect 12382 671 12388 705
rect 12422 671 12428 705
rect 12382 633 12428 671
rect 12382 599 12388 633
rect 12422 599 12428 633
rect 12382 561 12428 599
rect 12382 527 12388 561
rect 12422 527 12428 561
rect 12382 489 12428 527
rect 12382 455 12388 489
rect 12422 455 12428 489
rect 12382 417 12428 455
rect 12382 383 12388 417
rect 12422 383 12428 417
rect 12382 345 12428 383
rect 12382 311 12388 345
rect 12422 311 12428 345
rect 12382 273 12428 311
rect 12382 239 12388 273
rect 12422 239 12428 273
rect 12382 224 12428 239
rect 12478 1209 12524 1224
rect 12478 1175 12484 1209
rect 12518 1175 12524 1209
rect 12478 1137 12524 1175
rect 12478 1103 12484 1137
rect 12518 1103 12524 1137
rect 12478 1065 12524 1103
rect 12478 1031 12484 1065
rect 12518 1031 12524 1065
rect 12478 993 12524 1031
rect 12478 959 12484 993
rect 12518 959 12524 993
rect 12478 921 12524 959
rect 12478 887 12484 921
rect 12518 887 12524 921
rect 12478 849 12524 887
rect 12478 815 12484 849
rect 12518 815 12524 849
rect 12478 777 12524 815
rect 12478 743 12484 777
rect 12518 743 12524 777
rect 12478 705 12524 743
rect 12478 671 12484 705
rect 12518 671 12524 705
rect 12478 633 12524 671
rect 12478 599 12484 633
rect 12518 599 12524 633
rect 12478 561 12524 599
rect 12478 527 12484 561
rect 12518 527 12524 561
rect 12478 489 12524 527
rect 12478 455 12484 489
rect 12518 455 12524 489
rect 12478 417 12524 455
rect 12478 383 12484 417
rect 12518 383 12524 417
rect 12478 345 12524 383
rect 12478 311 12484 345
rect 12518 311 12524 345
rect 12478 273 12524 311
rect 12478 239 12484 273
rect 12518 239 12524 273
rect 12478 224 12524 239
rect 12574 1209 12620 1224
rect 12574 1175 12580 1209
rect 12614 1175 12620 1209
rect 12574 1137 12620 1175
rect 12574 1103 12580 1137
rect 12614 1103 12620 1137
rect 12574 1065 12620 1103
rect 12574 1031 12580 1065
rect 12614 1031 12620 1065
rect 12574 993 12620 1031
rect 12574 959 12580 993
rect 12614 959 12620 993
rect 12574 921 12620 959
rect 12574 887 12580 921
rect 12614 887 12620 921
rect 12574 849 12620 887
rect 12574 815 12580 849
rect 12614 815 12620 849
rect 12574 777 12620 815
rect 12574 743 12580 777
rect 12614 743 12620 777
rect 12574 705 12620 743
rect 12574 671 12580 705
rect 12614 671 12620 705
rect 12574 633 12620 671
rect 12574 599 12580 633
rect 12614 599 12620 633
rect 12574 561 12620 599
rect 12574 527 12580 561
rect 12614 527 12620 561
rect 12574 489 12620 527
rect 12574 455 12580 489
rect 12614 455 12620 489
rect 12574 417 12620 455
rect 12574 383 12580 417
rect 12614 383 12620 417
rect 12574 345 12620 383
rect 12574 311 12580 345
rect 12614 311 12620 345
rect 12574 273 12620 311
rect 12574 239 12580 273
rect 12614 239 12620 273
rect 12574 224 12620 239
rect 12670 1209 12716 1224
rect 12670 1175 12676 1209
rect 12710 1175 12716 1209
rect 12670 1137 12716 1175
rect 12670 1103 12676 1137
rect 12710 1103 12716 1137
rect 12670 1065 12716 1103
rect 12670 1031 12676 1065
rect 12710 1031 12716 1065
rect 12670 993 12716 1031
rect 12670 959 12676 993
rect 12710 959 12716 993
rect 12670 921 12716 959
rect 12670 887 12676 921
rect 12710 887 12716 921
rect 12670 849 12716 887
rect 12670 815 12676 849
rect 12710 815 12716 849
rect 12670 777 12716 815
rect 12670 743 12676 777
rect 12710 743 12716 777
rect 12670 705 12716 743
rect 12670 671 12676 705
rect 12710 671 12716 705
rect 12670 633 12716 671
rect 12670 599 12676 633
rect 12710 599 12716 633
rect 12670 561 12716 599
rect 12670 527 12676 561
rect 12710 527 12716 561
rect 12670 489 12716 527
rect 12670 455 12676 489
rect 12710 455 12716 489
rect 12670 417 12716 455
rect 12670 383 12676 417
rect 12710 383 12716 417
rect 12670 345 12716 383
rect 12670 311 12676 345
rect 12710 311 12716 345
rect 12670 273 12716 311
rect 12670 239 12676 273
rect 12710 239 12716 273
rect 12670 224 12716 239
rect 12766 1209 12812 1224
rect 12766 1175 12772 1209
rect 12806 1175 12812 1209
rect 12766 1137 12812 1175
rect 12766 1103 12772 1137
rect 12806 1103 12812 1137
rect 12766 1065 12812 1103
rect 12766 1031 12772 1065
rect 12806 1031 12812 1065
rect 12766 993 12812 1031
rect 12766 959 12772 993
rect 12806 959 12812 993
rect 12766 921 12812 959
rect 12766 887 12772 921
rect 12806 887 12812 921
rect 12766 849 12812 887
rect 12766 815 12772 849
rect 12806 815 12812 849
rect 12766 777 12812 815
rect 12766 743 12772 777
rect 12806 743 12812 777
rect 12766 705 12812 743
rect 12766 671 12772 705
rect 12806 671 12812 705
rect 12766 633 12812 671
rect 12766 599 12772 633
rect 12806 599 12812 633
rect 12766 561 12812 599
rect 12766 527 12772 561
rect 12806 527 12812 561
rect 12766 489 12812 527
rect 12766 455 12772 489
rect 12806 455 12812 489
rect 12766 417 12812 455
rect 12766 383 12772 417
rect 12806 383 12812 417
rect 12766 345 12812 383
rect 12766 311 12772 345
rect 12806 311 12812 345
rect 12766 273 12812 311
rect 12766 239 12772 273
rect 12806 239 12812 273
rect 12766 224 12812 239
rect 12862 1209 12908 1224
rect 12862 1175 12868 1209
rect 12902 1175 12908 1209
rect 12862 1137 12908 1175
rect 12862 1103 12868 1137
rect 12902 1103 12908 1137
rect 12862 1065 12908 1103
rect 12862 1031 12868 1065
rect 12902 1031 12908 1065
rect 12862 993 12908 1031
rect 12862 959 12868 993
rect 12902 959 12908 993
rect 12862 921 12908 959
rect 12862 887 12868 921
rect 12902 887 12908 921
rect 12862 849 12908 887
rect 12862 815 12868 849
rect 12902 815 12908 849
rect 12862 777 12908 815
rect 12862 743 12868 777
rect 12902 743 12908 777
rect 12862 705 12908 743
rect 12862 671 12868 705
rect 12902 671 12908 705
rect 12862 633 12908 671
rect 12862 599 12868 633
rect 12902 599 12908 633
rect 12862 561 12908 599
rect 12862 527 12868 561
rect 12902 527 12908 561
rect 12862 489 12908 527
rect 12862 455 12868 489
rect 12902 455 12908 489
rect 12862 417 12908 455
rect 12862 383 12868 417
rect 12902 383 12908 417
rect 12862 345 12908 383
rect 12862 311 12868 345
rect 12902 311 12908 345
rect 12862 273 12908 311
rect 12862 239 12868 273
rect 12902 239 12908 273
rect 12862 224 12908 239
rect 12958 1209 13004 1224
rect 12958 1175 12964 1209
rect 12998 1175 13004 1209
rect 12958 1137 13004 1175
rect 12958 1103 12964 1137
rect 12998 1103 13004 1137
rect 12958 1065 13004 1103
rect 12958 1031 12964 1065
rect 12998 1031 13004 1065
rect 12958 993 13004 1031
rect 12958 959 12964 993
rect 12998 959 13004 993
rect 12958 921 13004 959
rect 12958 887 12964 921
rect 12998 887 13004 921
rect 12958 849 13004 887
rect 12958 815 12964 849
rect 12998 815 13004 849
rect 12958 777 13004 815
rect 12958 743 12964 777
rect 12998 743 13004 777
rect 12958 705 13004 743
rect 12958 671 12964 705
rect 12998 671 13004 705
rect 12958 633 13004 671
rect 12958 599 12964 633
rect 12998 599 13004 633
rect 12958 561 13004 599
rect 12958 527 12964 561
rect 12998 527 13004 561
rect 12958 489 13004 527
rect 12958 455 12964 489
rect 12998 455 13004 489
rect 12958 417 13004 455
rect 12958 383 12964 417
rect 12998 383 13004 417
rect 12958 345 13004 383
rect 12958 311 12964 345
rect 12998 311 13004 345
rect 12958 273 13004 311
rect 12958 239 12964 273
rect 12998 239 13004 273
rect 12958 224 13004 239
rect 13054 1209 13100 1224
rect 13054 1175 13060 1209
rect 13094 1175 13100 1209
rect 13054 1137 13100 1175
rect 13054 1103 13060 1137
rect 13094 1103 13100 1137
rect 13054 1065 13100 1103
rect 13054 1031 13060 1065
rect 13094 1031 13100 1065
rect 13054 993 13100 1031
rect 13054 959 13060 993
rect 13094 959 13100 993
rect 13054 921 13100 959
rect 13054 887 13060 921
rect 13094 887 13100 921
rect 13054 849 13100 887
rect 13054 815 13060 849
rect 13094 815 13100 849
rect 13054 777 13100 815
rect 13054 743 13060 777
rect 13094 743 13100 777
rect 13054 705 13100 743
rect 13054 671 13060 705
rect 13094 671 13100 705
rect 13054 633 13100 671
rect 13054 599 13060 633
rect 13094 599 13100 633
rect 13054 561 13100 599
rect 13054 527 13060 561
rect 13094 527 13100 561
rect 13054 489 13100 527
rect 13054 455 13060 489
rect 13094 455 13100 489
rect 13054 417 13100 455
rect 13054 383 13060 417
rect 13094 383 13100 417
rect 13054 345 13100 383
rect 13054 311 13060 345
rect 13094 311 13100 345
rect 13054 273 13100 311
rect 13054 239 13060 273
rect 13094 239 13100 273
rect 13054 224 13100 239
rect 13150 1209 13196 1224
rect 13150 1175 13156 1209
rect 13190 1175 13196 1209
rect 13150 1137 13196 1175
rect 13150 1103 13156 1137
rect 13190 1103 13196 1137
rect 13150 1065 13196 1103
rect 13150 1031 13156 1065
rect 13190 1031 13196 1065
rect 13150 993 13196 1031
rect 13150 959 13156 993
rect 13190 959 13196 993
rect 13150 921 13196 959
rect 13150 887 13156 921
rect 13190 887 13196 921
rect 13150 849 13196 887
rect 13150 815 13156 849
rect 13190 815 13196 849
rect 13150 777 13196 815
rect 13150 743 13156 777
rect 13190 743 13196 777
rect 13150 705 13196 743
rect 13150 671 13156 705
rect 13190 671 13196 705
rect 13150 633 13196 671
rect 13150 599 13156 633
rect 13190 599 13196 633
rect 13150 561 13196 599
rect 13150 527 13156 561
rect 13190 527 13196 561
rect 13150 489 13196 527
rect 13150 455 13156 489
rect 13190 455 13196 489
rect 13150 417 13196 455
rect 13150 383 13156 417
rect 13190 383 13196 417
rect 13150 345 13196 383
rect 13150 311 13156 345
rect 13190 311 13196 345
rect 13150 273 13196 311
rect 13150 239 13156 273
rect 13190 239 13196 273
rect 13150 224 13196 239
rect 13246 1209 13292 1224
rect 13246 1175 13252 1209
rect 13286 1175 13292 1209
rect 13246 1137 13292 1175
rect 13246 1103 13252 1137
rect 13286 1103 13292 1137
rect 13246 1065 13292 1103
rect 13246 1031 13252 1065
rect 13286 1031 13292 1065
rect 13246 993 13292 1031
rect 13246 959 13252 993
rect 13286 959 13292 993
rect 13246 921 13292 959
rect 13246 887 13252 921
rect 13286 887 13292 921
rect 13246 849 13292 887
rect 13246 815 13252 849
rect 13286 815 13292 849
rect 13246 777 13292 815
rect 13246 743 13252 777
rect 13286 743 13292 777
rect 13246 705 13292 743
rect 13246 671 13252 705
rect 13286 671 13292 705
rect 13246 633 13292 671
rect 13246 599 13252 633
rect 13286 599 13292 633
rect 13246 561 13292 599
rect 13246 527 13252 561
rect 13286 527 13292 561
rect 13246 489 13292 527
rect 13246 455 13252 489
rect 13286 455 13292 489
rect 13246 417 13292 455
rect 13246 383 13252 417
rect 13286 383 13292 417
rect 13246 345 13292 383
rect 13246 311 13252 345
rect 13286 311 13292 345
rect 13246 273 13292 311
rect 13246 239 13252 273
rect 13286 239 13292 273
rect 13246 224 13292 239
rect 13342 1209 13388 1224
rect 13342 1175 13348 1209
rect 13382 1175 13388 1209
rect 13342 1137 13388 1175
rect 13342 1103 13348 1137
rect 13382 1103 13388 1137
rect 13342 1065 13388 1103
rect 13342 1031 13348 1065
rect 13382 1031 13388 1065
rect 13342 993 13388 1031
rect 13342 959 13348 993
rect 13382 959 13388 993
rect 13342 921 13388 959
rect 13342 887 13348 921
rect 13382 887 13388 921
rect 13342 849 13388 887
rect 13342 815 13348 849
rect 13382 815 13388 849
rect 13342 777 13388 815
rect 13342 743 13348 777
rect 13382 743 13388 777
rect 13342 705 13388 743
rect 13342 671 13348 705
rect 13382 671 13388 705
rect 13342 633 13388 671
rect 13342 599 13348 633
rect 13382 599 13388 633
rect 13342 561 13388 599
rect 13342 527 13348 561
rect 13382 527 13388 561
rect 13342 489 13388 527
rect 13342 455 13348 489
rect 13382 455 13388 489
rect 13342 417 13388 455
rect 13342 383 13348 417
rect 13382 383 13388 417
rect 13342 345 13388 383
rect 13342 311 13348 345
rect 13382 311 13388 345
rect 13342 273 13388 311
rect 13342 239 13348 273
rect 13382 239 13388 273
rect 13342 224 13388 239
rect 13438 1209 13484 1224
rect 13438 1175 13444 1209
rect 13478 1175 13484 1209
rect 13438 1137 13484 1175
rect 13438 1103 13444 1137
rect 13478 1103 13484 1137
rect 13438 1065 13484 1103
rect 13438 1031 13444 1065
rect 13478 1031 13484 1065
rect 13438 993 13484 1031
rect 13438 959 13444 993
rect 13478 959 13484 993
rect 13438 921 13484 959
rect 13438 887 13444 921
rect 13478 887 13484 921
rect 13438 849 13484 887
rect 13438 815 13444 849
rect 13478 815 13484 849
rect 13438 777 13484 815
rect 13438 743 13444 777
rect 13478 743 13484 777
rect 13438 705 13484 743
rect 13438 671 13444 705
rect 13478 671 13484 705
rect 13438 633 13484 671
rect 13438 599 13444 633
rect 13478 599 13484 633
rect 13438 561 13484 599
rect 13438 527 13444 561
rect 13478 527 13484 561
rect 13438 489 13484 527
rect 13438 455 13444 489
rect 13478 455 13484 489
rect 13438 417 13484 455
rect 13438 383 13444 417
rect 13478 383 13484 417
rect 13438 345 13484 383
rect 13438 311 13444 345
rect 13478 311 13484 345
rect 13438 273 13484 311
rect 13438 239 13444 273
rect 13478 239 13484 273
rect 13438 224 13484 239
rect 13534 1209 13580 1224
rect 13534 1175 13540 1209
rect 13574 1175 13580 1209
rect 13534 1137 13580 1175
rect 13534 1103 13540 1137
rect 13574 1103 13580 1137
rect 13534 1065 13580 1103
rect 13534 1031 13540 1065
rect 13574 1031 13580 1065
rect 13534 993 13580 1031
rect 13534 959 13540 993
rect 13574 959 13580 993
rect 13534 921 13580 959
rect 13534 887 13540 921
rect 13574 887 13580 921
rect 13534 849 13580 887
rect 13534 815 13540 849
rect 13574 815 13580 849
rect 13534 777 13580 815
rect 13534 743 13540 777
rect 13574 743 13580 777
rect 13534 705 13580 743
rect 13534 671 13540 705
rect 13574 671 13580 705
rect 13534 633 13580 671
rect 13534 599 13540 633
rect 13574 599 13580 633
rect 13534 561 13580 599
rect 13534 527 13540 561
rect 13574 527 13580 561
rect 13534 489 13580 527
rect 13534 455 13540 489
rect 13574 455 13580 489
rect 13534 417 13580 455
rect 13534 383 13540 417
rect 13574 383 13580 417
rect 13534 345 13580 383
rect 13534 311 13540 345
rect 13574 311 13580 345
rect 13534 273 13580 311
rect 13534 239 13540 273
rect 13574 239 13580 273
rect 13534 224 13580 239
rect 14150 1209 14196 1224
rect 14150 1175 14156 1209
rect 14190 1175 14196 1209
rect 14150 1137 14196 1175
rect 14150 1103 14156 1137
rect 14190 1103 14196 1137
rect 14150 1065 14196 1103
rect 14150 1031 14156 1065
rect 14190 1031 14196 1065
rect 14150 993 14196 1031
rect 14150 959 14156 993
rect 14190 959 14196 993
rect 14150 921 14196 959
rect 14150 887 14156 921
rect 14190 887 14196 921
rect 14150 849 14196 887
rect 14150 815 14156 849
rect 14190 815 14196 849
rect 14150 777 14196 815
rect 14150 743 14156 777
rect 14190 743 14196 777
rect 14150 705 14196 743
rect 14150 671 14156 705
rect 14190 671 14196 705
rect 14150 633 14196 671
rect 14150 599 14156 633
rect 14190 599 14196 633
rect 14150 561 14196 599
rect 14150 527 14156 561
rect 14190 527 14196 561
rect 14150 489 14196 527
rect 14150 455 14156 489
rect 14190 455 14196 489
rect 14150 417 14196 455
rect 14150 383 14156 417
rect 14190 383 14196 417
rect 14150 345 14196 383
rect 14150 311 14156 345
rect 14190 311 14196 345
rect 14150 273 14196 311
rect 14150 239 14156 273
rect 14190 239 14196 273
rect 14150 224 14196 239
rect 14246 1209 14292 1224
rect 14246 1175 14252 1209
rect 14286 1175 14292 1209
rect 14246 1137 14292 1175
rect 14246 1103 14252 1137
rect 14286 1103 14292 1137
rect 14246 1065 14292 1103
rect 14246 1031 14252 1065
rect 14286 1031 14292 1065
rect 14246 993 14292 1031
rect 14246 959 14252 993
rect 14286 959 14292 993
rect 14246 921 14292 959
rect 14246 887 14252 921
rect 14286 887 14292 921
rect 14246 849 14292 887
rect 14246 815 14252 849
rect 14286 815 14292 849
rect 14246 777 14292 815
rect 14246 743 14252 777
rect 14286 743 14292 777
rect 14246 705 14292 743
rect 14246 671 14252 705
rect 14286 671 14292 705
rect 14246 633 14292 671
rect 14246 599 14252 633
rect 14286 599 14292 633
rect 14246 561 14292 599
rect 14246 527 14252 561
rect 14286 527 14292 561
rect 14246 489 14292 527
rect 14246 455 14252 489
rect 14286 455 14292 489
rect 14246 417 14292 455
rect 14246 383 14252 417
rect 14286 383 14292 417
rect 14246 345 14292 383
rect 14246 311 14252 345
rect 14286 311 14292 345
rect 14246 273 14292 311
rect 14246 239 14252 273
rect 14286 239 14292 273
rect 14246 224 14292 239
rect 14342 1209 14388 1224
rect 14342 1175 14348 1209
rect 14382 1175 14388 1209
rect 14342 1137 14388 1175
rect 14342 1103 14348 1137
rect 14382 1103 14388 1137
rect 14342 1065 14388 1103
rect 14342 1031 14348 1065
rect 14382 1031 14388 1065
rect 14342 993 14388 1031
rect 14342 959 14348 993
rect 14382 959 14388 993
rect 14342 921 14388 959
rect 14342 887 14348 921
rect 14382 887 14388 921
rect 14342 849 14388 887
rect 14342 815 14348 849
rect 14382 815 14388 849
rect 14342 777 14388 815
rect 14342 743 14348 777
rect 14382 743 14388 777
rect 14342 705 14388 743
rect 14342 671 14348 705
rect 14382 671 14388 705
rect 14342 633 14388 671
rect 14342 599 14348 633
rect 14382 599 14388 633
rect 14342 561 14388 599
rect 14342 527 14348 561
rect 14382 527 14388 561
rect 14342 489 14388 527
rect 14342 455 14348 489
rect 14382 455 14388 489
rect 14342 417 14388 455
rect 14342 383 14348 417
rect 14382 383 14388 417
rect 14342 345 14388 383
rect 14342 311 14348 345
rect 14382 311 14388 345
rect 14342 273 14388 311
rect 14342 239 14348 273
rect 14382 239 14388 273
rect 14342 224 14388 239
rect 14438 1209 14484 1224
rect 14438 1175 14444 1209
rect 14478 1175 14484 1209
rect 14438 1137 14484 1175
rect 14438 1103 14444 1137
rect 14478 1103 14484 1137
rect 14438 1065 14484 1103
rect 14438 1031 14444 1065
rect 14478 1031 14484 1065
rect 14438 993 14484 1031
rect 14438 959 14444 993
rect 14478 959 14484 993
rect 14438 921 14484 959
rect 14438 887 14444 921
rect 14478 887 14484 921
rect 14438 849 14484 887
rect 14438 815 14444 849
rect 14478 815 14484 849
rect 14438 777 14484 815
rect 14438 743 14444 777
rect 14478 743 14484 777
rect 14438 705 14484 743
rect 14438 671 14444 705
rect 14478 671 14484 705
rect 14438 633 14484 671
rect 14438 599 14444 633
rect 14478 599 14484 633
rect 14438 561 14484 599
rect 14438 527 14444 561
rect 14478 527 14484 561
rect 14438 489 14484 527
rect 14438 455 14444 489
rect 14478 455 14484 489
rect 14438 417 14484 455
rect 14438 383 14444 417
rect 14478 383 14484 417
rect 14438 345 14484 383
rect 14438 311 14444 345
rect 14478 311 14484 345
rect 14438 273 14484 311
rect 14438 239 14444 273
rect 14478 239 14484 273
rect 14438 224 14484 239
rect 14534 1209 14580 1224
rect 14534 1175 14540 1209
rect 14574 1175 14580 1209
rect 14534 1137 14580 1175
rect 14534 1103 14540 1137
rect 14574 1103 14580 1137
rect 14534 1065 14580 1103
rect 14534 1031 14540 1065
rect 14574 1031 14580 1065
rect 14534 993 14580 1031
rect 14534 959 14540 993
rect 14574 959 14580 993
rect 14534 921 14580 959
rect 14534 887 14540 921
rect 14574 887 14580 921
rect 14534 849 14580 887
rect 14534 815 14540 849
rect 14574 815 14580 849
rect 14534 777 14580 815
rect 14534 743 14540 777
rect 14574 743 14580 777
rect 14534 705 14580 743
rect 14534 671 14540 705
rect 14574 671 14580 705
rect 14534 633 14580 671
rect 14534 599 14540 633
rect 14574 599 14580 633
rect 14534 561 14580 599
rect 14534 527 14540 561
rect 14574 527 14580 561
rect 14534 489 14580 527
rect 14534 455 14540 489
rect 14574 455 14580 489
rect 14534 417 14580 455
rect 14534 383 14540 417
rect 14574 383 14580 417
rect 14534 345 14580 383
rect 14534 311 14540 345
rect 14574 311 14580 345
rect 14534 273 14580 311
rect 14534 239 14540 273
rect 14574 239 14580 273
rect 14534 224 14580 239
rect 14630 1209 14676 1224
rect 14630 1175 14636 1209
rect 14670 1175 14676 1209
rect 14630 1137 14676 1175
rect 14630 1103 14636 1137
rect 14670 1103 14676 1137
rect 14630 1065 14676 1103
rect 14630 1031 14636 1065
rect 14670 1031 14676 1065
rect 14630 993 14676 1031
rect 14630 959 14636 993
rect 14670 959 14676 993
rect 14630 921 14676 959
rect 14630 887 14636 921
rect 14670 887 14676 921
rect 14630 849 14676 887
rect 14630 815 14636 849
rect 14670 815 14676 849
rect 14630 777 14676 815
rect 14630 743 14636 777
rect 14670 743 14676 777
rect 14630 705 14676 743
rect 14630 671 14636 705
rect 14670 671 14676 705
rect 14630 633 14676 671
rect 14630 599 14636 633
rect 14670 599 14676 633
rect 14630 561 14676 599
rect 14630 527 14636 561
rect 14670 527 14676 561
rect 14630 489 14676 527
rect 14630 455 14636 489
rect 14670 455 14676 489
rect 14630 417 14676 455
rect 14630 383 14636 417
rect 14670 383 14676 417
rect 14630 345 14676 383
rect 14630 311 14636 345
rect 14670 311 14676 345
rect 14630 273 14676 311
rect 14630 239 14636 273
rect 14670 239 14676 273
rect 14630 224 14676 239
rect 14726 1209 14772 1224
rect 14726 1175 14732 1209
rect 14766 1175 14772 1209
rect 14726 1137 14772 1175
rect 14726 1103 14732 1137
rect 14766 1103 14772 1137
rect 14726 1065 14772 1103
rect 14726 1031 14732 1065
rect 14766 1031 14772 1065
rect 14726 993 14772 1031
rect 14726 959 14732 993
rect 14766 959 14772 993
rect 14726 921 14772 959
rect 14726 887 14732 921
rect 14766 887 14772 921
rect 14726 849 14772 887
rect 14726 815 14732 849
rect 14766 815 14772 849
rect 14726 777 14772 815
rect 14726 743 14732 777
rect 14766 743 14772 777
rect 14726 705 14772 743
rect 14726 671 14732 705
rect 14766 671 14772 705
rect 14726 633 14772 671
rect 14726 599 14732 633
rect 14766 599 14772 633
rect 14726 561 14772 599
rect 14726 527 14732 561
rect 14766 527 14772 561
rect 14726 489 14772 527
rect 14726 455 14732 489
rect 14766 455 14772 489
rect 14726 417 14772 455
rect 14726 383 14732 417
rect 14766 383 14772 417
rect 14726 345 14772 383
rect 14726 311 14732 345
rect 14766 311 14772 345
rect 14726 273 14772 311
rect 14726 239 14732 273
rect 14766 239 14772 273
rect 14726 224 14772 239
rect 14822 1209 14868 1224
rect 14822 1175 14828 1209
rect 14862 1175 14868 1209
rect 14822 1137 14868 1175
rect 14822 1103 14828 1137
rect 14862 1103 14868 1137
rect 14822 1065 14868 1103
rect 14822 1031 14828 1065
rect 14862 1031 14868 1065
rect 14822 993 14868 1031
rect 14822 959 14828 993
rect 14862 959 14868 993
rect 14822 921 14868 959
rect 14822 887 14828 921
rect 14862 887 14868 921
rect 14822 849 14868 887
rect 14822 815 14828 849
rect 14862 815 14868 849
rect 14822 777 14868 815
rect 14822 743 14828 777
rect 14862 743 14868 777
rect 14822 705 14868 743
rect 14822 671 14828 705
rect 14862 671 14868 705
rect 14822 633 14868 671
rect 14822 599 14828 633
rect 14862 599 14868 633
rect 14822 561 14868 599
rect 14822 527 14828 561
rect 14862 527 14868 561
rect 14822 489 14868 527
rect 14822 455 14828 489
rect 14862 455 14868 489
rect 14822 417 14868 455
rect 14822 383 14828 417
rect 14862 383 14868 417
rect 14822 345 14868 383
rect 14822 311 14828 345
rect 14862 311 14868 345
rect 14822 273 14868 311
rect 14822 239 14828 273
rect 14862 239 14868 273
rect 14822 224 14868 239
rect 14918 1209 14964 1224
rect 14918 1175 14924 1209
rect 14958 1175 14964 1209
rect 14918 1137 14964 1175
rect 14918 1103 14924 1137
rect 14958 1103 14964 1137
rect 14918 1065 14964 1103
rect 14918 1031 14924 1065
rect 14958 1031 14964 1065
rect 14918 993 14964 1031
rect 14918 959 14924 993
rect 14958 959 14964 993
rect 14918 921 14964 959
rect 14918 887 14924 921
rect 14958 887 14964 921
rect 14918 849 14964 887
rect 14918 815 14924 849
rect 14958 815 14964 849
rect 14918 777 14964 815
rect 14918 743 14924 777
rect 14958 743 14964 777
rect 14918 705 14964 743
rect 14918 671 14924 705
rect 14958 671 14964 705
rect 14918 633 14964 671
rect 14918 599 14924 633
rect 14958 599 14964 633
rect 14918 561 14964 599
rect 14918 527 14924 561
rect 14958 527 14964 561
rect 14918 489 14964 527
rect 14918 455 14924 489
rect 14958 455 14964 489
rect 14918 417 14964 455
rect 14918 383 14924 417
rect 14958 383 14964 417
rect 14918 345 14964 383
rect 14918 311 14924 345
rect 14958 311 14964 345
rect 14918 273 14964 311
rect 14918 239 14924 273
rect 14958 239 14964 273
rect 14918 224 14964 239
rect 15014 1209 15060 1224
rect 15014 1175 15020 1209
rect 15054 1175 15060 1209
rect 15014 1137 15060 1175
rect 15014 1103 15020 1137
rect 15054 1103 15060 1137
rect 15014 1065 15060 1103
rect 15014 1031 15020 1065
rect 15054 1031 15060 1065
rect 15014 993 15060 1031
rect 15014 959 15020 993
rect 15054 959 15060 993
rect 15014 921 15060 959
rect 15014 887 15020 921
rect 15054 887 15060 921
rect 15014 849 15060 887
rect 15014 815 15020 849
rect 15054 815 15060 849
rect 15014 777 15060 815
rect 15014 743 15020 777
rect 15054 743 15060 777
rect 15014 705 15060 743
rect 15014 671 15020 705
rect 15054 671 15060 705
rect 15014 633 15060 671
rect 15014 599 15020 633
rect 15054 599 15060 633
rect 15014 561 15060 599
rect 15014 527 15020 561
rect 15054 527 15060 561
rect 15014 489 15060 527
rect 15014 455 15020 489
rect 15054 455 15060 489
rect 15014 417 15060 455
rect 15014 383 15020 417
rect 15054 383 15060 417
rect 15014 345 15060 383
rect 15014 311 15020 345
rect 15054 311 15060 345
rect 15014 273 15060 311
rect 15014 239 15020 273
rect 15054 239 15060 273
rect 15014 224 15060 239
rect 15110 1209 15156 1224
rect 15110 1175 15116 1209
rect 15150 1175 15156 1209
rect 15110 1137 15156 1175
rect 15110 1103 15116 1137
rect 15150 1103 15156 1137
rect 15110 1065 15156 1103
rect 15110 1031 15116 1065
rect 15150 1031 15156 1065
rect 15110 993 15156 1031
rect 15110 959 15116 993
rect 15150 959 15156 993
rect 15110 921 15156 959
rect 15110 887 15116 921
rect 15150 887 15156 921
rect 15110 849 15156 887
rect 15110 815 15116 849
rect 15150 815 15156 849
rect 15110 777 15156 815
rect 15110 743 15116 777
rect 15150 743 15156 777
rect 15110 705 15156 743
rect 15110 671 15116 705
rect 15150 671 15156 705
rect 15110 633 15156 671
rect 15110 599 15116 633
rect 15150 599 15156 633
rect 15110 561 15156 599
rect 15110 527 15116 561
rect 15150 527 15156 561
rect 15110 489 15156 527
rect 15110 455 15116 489
rect 15150 455 15156 489
rect 15110 417 15156 455
rect 15110 383 15116 417
rect 15150 383 15156 417
rect 15110 345 15156 383
rect 15110 311 15116 345
rect 15150 311 15156 345
rect 15110 273 15156 311
rect 15110 239 15116 273
rect 15150 239 15156 273
rect 15110 224 15156 239
rect 15206 1209 15252 1224
rect 15206 1175 15212 1209
rect 15246 1175 15252 1209
rect 15206 1137 15252 1175
rect 15206 1103 15212 1137
rect 15246 1103 15252 1137
rect 15206 1065 15252 1103
rect 15206 1031 15212 1065
rect 15246 1031 15252 1065
rect 15206 993 15252 1031
rect 15206 959 15212 993
rect 15246 959 15252 993
rect 15206 921 15252 959
rect 15206 887 15212 921
rect 15246 887 15252 921
rect 15206 849 15252 887
rect 15206 815 15212 849
rect 15246 815 15252 849
rect 15206 777 15252 815
rect 15206 743 15212 777
rect 15246 743 15252 777
rect 15206 705 15252 743
rect 15206 671 15212 705
rect 15246 671 15252 705
rect 15206 633 15252 671
rect 15206 599 15212 633
rect 15246 599 15252 633
rect 15206 561 15252 599
rect 15206 527 15212 561
rect 15246 527 15252 561
rect 15206 489 15252 527
rect 15206 455 15212 489
rect 15246 455 15252 489
rect 15206 417 15252 455
rect 15206 383 15212 417
rect 15246 383 15252 417
rect 15206 345 15252 383
rect 15206 311 15212 345
rect 15246 311 15252 345
rect 15206 273 15252 311
rect 15206 239 15212 273
rect 15246 239 15252 273
rect 15206 224 15252 239
rect 15416 1223 15422 1257
rect 15456 1223 15462 1257
rect 15416 1185 15462 1223
rect 15416 1151 15422 1185
rect 15456 1151 15462 1185
rect 15416 1113 15462 1151
rect 15416 1079 15422 1113
rect 15456 1079 15462 1113
rect 15416 1041 15462 1079
rect 15416 1007 15422 1041
rect 15456 1007 15462 1041
rect 15416 969 15462 1007
rect 15416 935 15422 969
rect 15456 935 15462 969
rect 15416 897 15462 935
rect 15416 863 15422 897
rect 15456 863 15462 897
rect 15416 825 15462 863
rect 15416 791 15422 825
rect 15456 791 15462 825
rect 15416 753 15462 791
rect 15416 719 15422 753
rect 15456 719 15462 753
rect 15416 681 15462 719
rect 15416 647 15422 681
rect 15456 647 15462 681
rect 15416 609 15462 647
rect 15416 575 15422 609
rect 15456 575 15462 609
rect 15416 537 15462 575
rect 15416 503 15422 537
rect 15456 503 15462 537
rect 15416 465 15462 503
rect 15416 431 15422 465
rect 15456 431 15462 465
rect 15416 393 15462 431
rect 15416 359 15422 393
rect 15456 359 15462 393
rect 15416 321 15462 359
rect 15416 287 15422 321
rect 15456 287 15462 321
rect 15416 249 15462 287
rect 15416 215 15422 249
rect 15456 215 15462 249
rect 15416 177 15462 215
rect 2482 146 2540 160
rect 142 130 204 144
rect 142 96 156 130
rect 190 96 204 130
rect 142 -76 204 96
rect 818 120 876 130
rect 818 86 830 120
rect 864 86 876 120
rect 818 40 876 86
rect 2482 112 2494 146
rect 2528 112 2540 146
rect 2482 40 2540 112
rect 2774 130 2836 144
rect 2774 96 2788 130
rect 2822 96 2836 130
rect 5438 130 5496 144
rect 818 30 2544 40
rect 818 -6 1498 30
rect 1720 -6 2544 30
rect 818 -20 2544 -6
rect 2774 -15 2836 96
rect 2774 -67 2779 -15
rect 2831 -67 2836 -15
rect 142 -126 206 -76
rect 2774 -82 2836 -67
rect 3098 114 3160 128
rect 3098 80 3112 114
rect 3146 80 3160 114
rect 3098 -76 3160 80
rect 3774 104 3832 114
rect 3774 70 3786 104
rect 3820 70 3832 104
rect 3774 24 3832 70
rect 5438 96 5450 130
rect 5484 96 5496 130
rect 8468 130 8526 144
rect 15416 143 15422 177
rect 15456 143 15462 177
rect 5438 24 5496 96
rect 5730 122 5790 124
rect 5730 114 5792 122
rect 5730 80 5744 114
rect 5778 80 5792 114
rect 3774 12 5500 24
rect 3774 -24 4584 12
rect 4806 -24 5500 12
rect 3774 -36 5500 -24
rect 5730 -11 5792 80
rect 5730 -63 5735 -11
rect 5787 -63 5792 -11
rect 3098 -126 3162 -76
rect 5730 -78 5792 -63
rect 6128 114 6190 126
rect 6128 80 6142 114
rect 6176 80 6190 114
rect 6128 -78 6190 80
rect 6804 104 6862 114
rect 6804 70 6816 104
rect 6850 70 6862 104
rect 6804 24 6862 70
rect 8468 96 8480 130
rect 8514 96 8526 130
rect 11556 128 11614 142
rect 8468 24 8526 96
rect 8760 122 8820 124
rect 8760 114 8822 122
rect 8760 80 8774 114
rect 8808 80 8822 114
rect 6804 18 8530 24
rect 6804 -16 7632 18
rect 7854 -16 8530 18
rect 6804 -36 8530 -16
rect 8760 -25 8822 80
rect 6126 -126 6190 -78
rect 8760 -77 8765 -25
rect 8817 -77 8822 -25
rect 8760 -92 8822 -77
rect 9214 112 9276 128
rect 9214 78 9230 112
rect 9264 78 9276 112
rect 9214 -76 9276 78
rect 9892 102 9950 112
rect 9892 68 9904 102
rect 9938 68 9950 102
rect 9892 22 9950 68
rect 11556 94 11568 128
rect 11602 94 11614 128
rect 11556 22 11614 94
rect 11848 112 11910 122
rect 11848 78 11862 112
rect 11896 78 11910 112
rect 9892 12 11618 22
rect 9892 -24 10562 12
rect 10796 -24 11618 12
rect 9892 -38 11618 -24
rect 11848 -25 11910 78
rect 9214 -126 9278 -76
rect 11848 -77 11853 -25
rect 11905 -77 11910 -25
rect 11848 -92 11910 -77
rect 12346 86 12464 104
rect 14712 102 14770 116
rect 12346 52 12386 86
rect 12420 52 12464 86
rect 12346 -126 12464 52
rect 13048 76 13106 86
rect 13048 42 13060 76
rect 13094 42 13106 76
rect 13048 -4 13106 42
rect 14712 68 14724 102
rect 14758 68 14770 102
rect 15416 100 15462 143
rect 15504 1257 15550 1300
rect 15504 1223 15510 1257
rect 15544 1223 15550 1257
rect 15504 1185 15550 1223
rect 15504 1151 15510 1185
rect 15544 1151 15550 1185
rect 15504 1113 15550 1151
rect 15504 1079 15510 1113
rect 15544 1079 15550 1113
rect 15504 1041 15550 1079
rect 15504 1007 15510 1041
rect 15544 1007 15550 1041
rect 15504 969 15550 1007
rect 15504 935 15510 969
rect 15544 935 15550 969
rect 15504 897 15550 935
rect 15504 863 15510 897
rect 15544 863 15550 897
rect 15504 825 15550 863
rect 15504 791 15510 825
rect 15544 791 15550 825
rect 15504 753 15550 791
rect 15504 719 15510 753
rect 15544 719 15550 753
rect 15504 681 15550 719
rect 15504 647 15510 681
rect 15544 647 15550 681
rect 15504 609 15550 647
rect 15504 575 15510 609
rect 15544 575 15550 609
rect 15504 537 15550 575
rect 15504 503 15510 537
rect 15544 503 15550 537
rect 15504 465 15550 503
rect 15504 431 15510 465
rect 15544 431 15550 465
rect 15504 393 15550 431
rect 15504 359 15510 393
rect 15544 359 15550 393
rect 15504 321 15550 359
rect 15504 287 15510 321
rect 15544 287 15550 321
rect 15504 249 15550 287
rect 15504 215 15510 249
rect 15544 215 15550 249
rect 15504 177 15550 215
rect 15504 143 15510 177
rect 15544 143 15550 177
rect 15504 100 15550 143
rect 14712 -4 14770 68
rect 15002 86 15064 98
rect 15002 52 15018 86
rect 15052 52 15064 86
rect 13048 -14 14774 -4
rect 13048 -50 13856 -14
rect 14090 -50 14774 -14
rect 13048 -64 14774 -50
rect -564 -280 12464 -126
rect 15002 -66 15064 52
rect 15322 52 15554 64
rect 15322 18 15510 52
rect 15544 18 15554 52
rect 15322 2 15554 18
rect 15322 -66 15384 2
rect 15002 -128 15384 -66
rect 15320 -258 15384 -128
rect 15698 -258 15760 3726
rect 16796 3706 16894 3742
rect 16796 3672 16830 3706
rect 16864 3672 16894 3706
rect 17498 3736 17578 3770
rect 17736 3819 18788 3850
rect 20348 3949 20460 3994
rect 20348 3915 20386 3949
rect 20420 3915 20460 3949
rect 20348 3832 20460 3915
rect 23284 3941 23382 3968
rect 23284 3907 23318 3941
rect 23352 3907 23382 3941
rect 23284 3844 23382 3907
rect 17736 3785 17790 3819
rect 17824 3785 18788 3819
rect 17736 3754 18788 3785
rect 17498 3702 17522 3736
rect 17556 3702 17578 3736
rect 17498 3680 17578 3702
rect 18688 3692 18788 3754
rect 19390 3806 20460 3832
rect 19390 3772 19443 3806
rect 19477 3772 20460 3806
rect 19390 3748 20460 3772
rect 21590 3804 22722 3824
rect 21590 3770 21646 3804
rect 21680 3770 22722 3804
rect 21590 3752 22722 3770
rect 16796 3646 16894 3672
rect 18688 3658 18720 3692
rect 18754 3658 18788 3692
rect 18688 3632 18788 3658
rect 20348 3690 20460 3748
rect 20348 3656 20388 3690
rect 20422 3656 20460 3690
rect 20348 3616 20460 3656
rect 16680 3519 16726 3534
rect 16680 3485 16686 3519
rect 16720 3485 16726 3519
rect 16680 3447 16726 3485
rect 16680 3413 16686 3447
rect 16720 3413 16726 3447
rect 16680 3375 16726 3413
rect 16680 3341 16686 3375
rect 16720 3341 16726 3375
rect 16680 3303 16726 3341
rect 16680 3269 16686 3303
rect 16720 3269 16726 3303
rect 16680 3231 16726 3269
rect 16680 3197 16686 3231
rect 16720 3197 16726 3231
rect 16680 3159 16726 3197
rect 16680 3125 16686 3159
rect 16720 3125 16726 3159
rect 16680 3087 16726 3125
rect 16680 3053 16686 3087
rect 16720 3053 16726 3087
rect 16680 3015 16726 3053
rect 16680 2981 16686 3015
rect 16720 2981 16726 3015
rect 16680 2943 16726 2981
rect 16680 2909 16686 2943
rect 16720 2909 16726 2943
rect 16680 2871 16726 2909
rect 16680 2837 16686 2871
rect 16720 2837 16726 2871
rect 16680 2799 16726 2837
rect 16680 2765 16686 2799
rect 16720 2765 16726 2799
rect 16680 2727 16726 2765
rect 16680 2693 16686 2727
rect 16720 2693 16726 2727
rect 16680 2655 16726 2693
rect 16680 2621 16686 2655
rect 16720 2621 16726 2655
rect 16680 2583 16726 2621
rect 16680 2549 16686 2583
rect 16720 2549 16726 2583
rect 16680 2534 16726 2549
rect 16776 3519 16822 3534
rect 16776 3485 16782 3519
rect 16816 3485 16822 3519
rect 16776 3447 16822 3485
rect 16776 3413 16782 3447
rect 16816 3413 16822 3447
rect 16776 3375 16822 3413
rect 16776 3341 16782 3375
rect 16816 3341 16822 3375
rect 16776 3303 16822 3341
rect 16776 3269 16782 3303
rect 16816 3269 16822 3303
rect 16776 3231 16822 3269
rect 16776 3197 16782 3231
rect 16816 3197 16822 3231
rect 16776 3159 16822 3197
rect 16776 3125 16782 3159
rect 16816 3125 16822 3159
rect 16776 3087 16822 3125
rect 16776 3053 16782 3087
rect 16816 3053 16822 3087
rect 16776 3015 16822 3053
rect 16776 2981 16782 3015
rect 16816 2981 16822 3015
rect 16776 2943 16822 2981
rect 16776 2909 16782 2943
rect 16816 2909 16822 2943
rect 16776 2871 16822 2909
rect 16776 2837 16782 2871
rect 16816 2837 16822 2871
rect 16776 2799 16822 2837
rect 16776 2765 16782 2799
rect 16816 2765 16822 2799
rect 16776 2727 16822 2765
rect 16776 2693 16782 2727
rect 16816 2693 16822 2727
rect 16776 2655 16822 2693
rect 16776 2621 16782 2655
rect 16816 2621 16822 2655
rect 16776 2583 16822 2621
rect 16776 2549 16782 2583
rect 16816 2549 16822 2583
rect 16776 2534 16822 2549
rect 16872 3519 16918 3534
rect 16872 3485 16878 3519
rect 16912 3485 16918 3519
rect 16872 3447 16918 3485
rect 16872 3413 16878 3447
rect 16912 3413 16918 3447
rect 16872 3375 16918 3413
rect 16872 3341 16878 3375
rect 16912 3341 16918 3375
rect 16872 3303 16918 3341
rect 16872 3269 16878 3303
rect 16912 3269 16918 3303
rect 16872 3231 16918 3269
rect 16872 3197 16878 3231
rect 16912 3197 16918 3231
rect 16872 3159 16918 3197
rect 16872 3125 16878 3159
rect 16912 3125 16918 3159
rect 16872 3087 16918 3125
rect 16872 3053 16878 3087
rect 16912 3053 16918 3087
rect 16872 3015 16918 3053
rect 16872 2981 16878 3015
rect 16912 2981 16918 3015
rect 16872 2943 16918 2981
rect 16872 2909 16878 2943
rect 16912 2909 16918 2943
rect 16872 2871 16918 2909
rect 16872 2837 16878 2871
rect 16912 2837 16918 2871
rect 16872 2799 16918 2837
rect 16872 2765 16878 2799
rect 16912 2765 16918 2799
rect 16872 2727 16918 2765
rect 16872 2693 16878 2727
rect 16912 2693 16918 2727
rect 16872 2655 16918 2693
rect 16872 2621 16878 2655
rect 16912 2621 16918 2655
rect 16872 2583 16918 2621
rect 16872 2549 16878 2583
rect 16912 2549 16918 2583
rect 16872 2534 16918 2549
rect 16968 3519 17014 3534
rect 16968 3485 16974 3519
rect 17008 3485 17014 3519
rect 16968 3447 17014 3485
rect 16968 3413 16974 3447
rect 17008 3413 17014 3447
rect 16968 3375 17014 3413
rect 16968 3341 16974 3375
rect 17008 3341 17014 3375
rect 16968 3303 17014 3341
rect 16968 3269 16974 3303
rect 17008 3269 17014 3303
rect 16968 3231 17014 3269
rect 16968 3197 16974 3231
rect 17008 3197 17014 3231
rect 16968 3159 17014 3197
rect 16968 3125 16974 3159
rect 17008 3125 17014 3159
rect 16968 3087 17014 3125
rect 16968 3053 16974 3087
rect 17008 3053 17014 3087
rect 16968 3015 17014 3053
rect 16968 2981 16974 3015
rect 17008 2981 17014 3015
rect 16968 2943 17014 2981
rect 16968 2909 16974 2943
rect 17008 2909 17014 2943
rect 16968 2871 17014 2909
rect 16968 2837 16974 2871
rect 17008 2837 17014 2871
rect 16968 2799 17014 2837
rect 16968 2765 16974 2799
rect 17008 2765 17014 2799
rect 16968 2727 17014 2765
rect 16968 2693 16974 2727
rect 17008 2693 17014 2727
rect 16968 2655 17014 2693
rect 16968 2621 16974 2655
rect 17008 2621 17014 2655
rect 16968 2583 17014 2621
rect 16968 2549 16974 2583
rect 17008 2549 17014 2583
rect 16968 2534 17014 2549
rect 17064 3519 17110 3534
rect 17064 3485 17070 3519
rect 17104 3485 17110 3519
rect 17064 3447 17110 3485
rect 17064 3413 17070 3447
rect 17104 3413 17110 3447
rect 17064 3375 17110 3413
rect 17064 3341 17070 3375
rect 17104 3341 17110 3375
rect 17064 3303 17110 3341
rect 17064 3269 17070 3303
rect 17104 3269 17110 3303
rect 17064 3231 17110 3269
rect 17064 3197 17070 3231
rect 17104 3197 17110 3231
rect 17064 3159 17110 3197
rect 17064 3125 17070 3159
rect 17104 3125 17110 3159
rect 17064 3087 17110 3125
rect 17064 3053 17070 3087
rect 17104 3053 17110 3087
rect 17064 3015 17110 3053
rect 17064 2981 17070 3015
rect 17104 2981 17110 3015
rect 17064 2943 17110 2981
rect 17064 2909 17070 2943
rect 17104 2909 17110 2943
rect 17064 2871 17110 2909
rect 17064 2837 17070 2871
rect 17104 2837 17110 2871
rect 17064 2799 17110 2837
rect 17064 2765 17070 2799
rect 17104 2765 17110 2799
rect 17064 2727 17110 2765
rect 17064 2693 17070 2727
rect 17104 2693 17110 2727
rect 17064 2655 17110 2693
rect 17064 2621 17070 2655
rect 17104 2621 17110 2655
rect 17064 2583 17110 2621
rect 17064 2549 17070 2583
rect 17104 2549 17110 2583
rect 17064 2534 17110 2549
rect 17160 3519 17206 3534
rect 17160 3485 17166 3519
rect 17200 3485 17206 3519
rect 17160 3447 17206 3485
rect 17160 3413 17166 3447
rect 17200 3413 17206 3447
rect 17160 3375 17206 3413
rect 17160 3341 17166 3375
rect 17200 3341 17206 3375
rect 17160 3303 17206 3341
rect 17160 3269 17166 3303
rect 17200 3269 17206 3303
rect 17160 3231 17206 3269
rect 17160 3197 17166 3231
rect 17200 3197 17206 3231
rect 17160 3159 17206 3197
rect 17160 3125 17166 3159
rect 17200 3125 17206 3159
rect 17160 3087 17206 3125
rect 17160 3053 17166 3087
rect 17200 3053 17206 3087
rect 17160 3015 17206 3053
rect 17160 2981 17166 3015
rect 17200 2981 17206 3015
rect 17160 2943 17206 2981
rect 17160 2909 17166 2943
rect 17200 2909 17206 2943
rect 17160 2871 17206 2909
rect 17160 2837 17166 2871
rect 17200 2837 17206 2871
rect 17160 2799 17206 2837
rect 17160 2765 17166 2799
rect 17200 2765 17206 2799
rect 17160 2727 17206 2765
rect 17160 2693 17166 2727
rect 17200 2693 17206 2727
rect 17160 2655 17206 2693
rect 17160 2621 17166 2655
rect 17200 2621 17206 2655
rect 17160 2583 17206 2621
rect 17160 2549 17166 2583
rect 17200 2549 17206 2583
rect 17160 2534 17206 2549
rect 17372 3509 17418 3524
rect 17372 3475 17378 3509
rect 17412 3475 17418 3509
rect 17372 3437 17418 3475
rect 17372 3403 17378 3437
rect 17412 3403 17418 3437
rect 17372 3365 17418 3403
rect 17372 3331 17378 3365
rect 17412 3331 17418 3365
rect 17372 3293 17418 3331
rect 17372 3259 17378 3293
rect 17412 3259 17418 3293
rect 17372 3221 17418 3259
rect 17372 3187 17378 3221
rect 17412 3187 17418 3221
rect 17372 3149 17418 3187
rect 17372 3115 17378 3149
rect 17412 3115 17418 3149
rect 17372 3077 17418 3115
rect 17372 3043 17378 3077
rect 17412 3043 17418 3077
rect 17372 3005 17418 3043
rect 17372 2971 17378 3005
rect 17412 2971 17418 3005
rect 17372 2933 17418 2971
rect 17372 2899 17378 2933
rect 17412 2899 17418 2933
rect 17372 2861 17418 2899
rect 17372 2827 17378 2861
rect 17412 2827 17418 2861
rect 17372 2789 17418 2827
rect 17372 2755 17378 2789
rect 17412 2755 17418 2789
rect 17372 2717 17418 2755
rect 17372 2683 17378 2717
rect 17412 2683 17418 2717
rect 17372 2645 17418 2683
rect 17372 2611 17378 2645
rect 17412 2611 17418 2645
rect 17372 2573 17418 2611
rect 17372 2539 17378 2573
rect 17412 2539 17418 2573
rect 17372 2524 17418 2539
rect 17468 3509 17514 3524
rect 17468 3475 17474 3509
rect 17508 3475 17514 3509
rect 17468 3437 17514 3475
rect 17468 3403 17474 3437
rect 17508 3403 17514 3437
rect 17468 3365 17514 3403
rect 17468 3331 17474 3365
rect 17508 3331 17514 3365
rect 17468 3293 17514 3331
rect 17468 3259 17474 3293
rect 17508 3259 17514 3293
rect 17468 3221 17514 3259
rect 17468 3187 17474 3221
rect 17508 3187 17514 3221
rect 17468 3149 17514 3187
rect 17468 3115 17474 3149
rect 17508 3115 17514 3149
rect 17468 3077 17514 3115
rect 17468 3043 17474 3077
rect 17508 3043 17514 3077
rect 17468 3005 17514 3043
rect 17468 2971 17474 3005
rect 17508 2971 17514 3005
rect 17468 2933 17514 2971
rect 17468 2899 17474 2933
rect 17508 2899 17514 2933
rect 17468 2861 17514 2899
rect 17468 2827 17474 2861
rect 17508 2827 17514 2861
rect 17468 2789 17514 2827
rect 17468 2755 17474 2789
rect 17508 2755 17514 2789
rect 17468 2717 17514 2755
rect 17468 2683 17474 2717
rect 17508 2683 17514 2717
rect 17468 2645 17514 2683
rect 17468 2611 17474 2645
rect 17508 2611 17514 2645
rect 17468 2573 17514 2611
rect 17468 2539 17474 2573
rect 17508 2539 17514 2573
rect 17468 2524 17514 2539
rect 17564 3509 17610 3524
rect 17564 3475 17570 3509
rect 17604 3475 17610 3509
rect 17564 3437 17610 3475
rect 17564 3403 17570 3437
rect 17604 3403 17610 3437
rect 17564 3365 17610 3403
rect 17564 3331 17570 3365
rect 17604 3331 17610 3365
rect 17564 3293 17610 3331
rect 17564 3259 17570 3293
rect 17604 3259 17610 3293
rect 17564 3221 17610 3259
rect 17564 3187 17570 3221
rect 17604 3187 17610 3221
rect 17564 3149 17610 3187
rect 17564 3115 17570 3149
rect 17604 3115 17610 3149
rect 17564 3077 17610 3115
rect 17564 3043 17570 3077
rect 17604 3043 17610 3077
rect 17564 3005 17610 3043
rect 17564 2971 17570 3005
rect 17604 2971 17610 3005
rect 17564 2933 17610 2971
rect 17564 2899 17570 2933
rect 17604 2899 17610 2933
rect 17564 2861 17610 2899
rect 17564 2827 17570 2861
rect 17604 2827 17610 2861
rect 17564 2789 17610 2827
rect 17564 2755 17570 2789
rect 17604 2755 17610 2789
rect 17564 2717 17610 2755
rect 17564 2683 17570 2717
rect 17604 2683 17610 2717
rect 17564 2645 17610 2683
rect 17564 2611 17570 2645
rect 17604 2611 17610 2645
rect 17564 2573 17610 2611
rect 17564 2539 17570 2573
rect 17604 2539 17610 2573
rect 17564 2524 17610 2539
rect 17660 3509 17706 3524
rect 17660 3475 17666 3509
rect 17700 3475 17706 3509
rect 17660 3437 17706 3475
rect 17660 3403 17666 3437
rect 17700 3403 17706 3437
rect 17660 3365 17706 3403
rect 17660 3331 17666 3365
rect 17700 3331 17706 3365
rect 17660 3293 17706 3331
rect 17660 3259 17666 3293
rect 17700 3259 17706 3293
rect 17660 3221 17706 3259
rect 17660 3187 17666 3221
rect 17700 3187 17706 3221
rect 17660 3149 17706 3187
rect 17660 3115 17666 3149
rect 17700 3115 17706 3149
rect 17660 3077 17706 3115
rect 17660 3043 17666 3077
rect 17700 3043 17706 3077
rect 17660 3005 17706 3043
rect 17660 2971 17666 3005
rect 17700 2971 17706 3005
rect 17660 2933 17706 2971
rect 17660 2899 17666 2933
rect 17700 2899 17706 2933
rect 17660 2861 17706 2899
rect 17660 2827 17666 2861
rect 17700 2827 17706 2861
rect 17660 2789 17706 2827
rect 17660 2755 17666 2789
rect 17700 2755 17706 2789
rect 17660 2717 17706 2755
rect 17660 2683 17666 2717
rect 17700 2683 17706 2717
rect 17660 2645 17706 2683
rect 17660 2611 17666 2645
rect 17700 2611 17706 2645
rect 17660 2573 17706 2611
rect 17660 2539 17666 2573
rect 17700 2539 17706 2573
rect 17660 2524 17706 2539
rect 17756 3509 17802 3524
rect 17756 3475 17762 3509
rect 17796 3475 17802 3509
rect 17756 3437 17802 3475
rect 17756 3403 17762 3437
rect 17796 3403 17802 3437
rect 17756 3365 17802 3403
rect 17756 3331 17762 3365
rect 17796 3331 17802 3365
rect 17756 3293 17802 3331
rect 17756 3259 17762 3293
rect 17796 3259 17802 3293
rect 17756 3221 17802 3259
rect 17756 3187 17762 3221
rect 17796 3187 17802 3221
rect 17756 3149 17802 3187
rect 17756 3115 17762 3149
rect 17796 3115 17802 3149
rect 17756 3077 17802 3115
rect 17756 3043 17762 3077
rect 17796 3043 17802 3077
rect 17756 3005 17802 3043
rect 17756 2971 17762 3005
rect 17796 2971 17802 3005
rect 17756 2933 17802 2971
rect 17756 2899 17762 2933
rect 17796 2899 17802 2933
rect 17756 2861 17802 2899
rect 17756 2827 17762 2861
rect 17796 2827 17802 2861
rect 17756 2789 17802 2827
rect 17756 2755 17762 2789
rect 17796 2755 17802 2789
rect 17756 2717 17802 2755
rect 17756 2683 17762 2717
rect 17796 2683 17802 2717
rect 17756 2645 17802 2683
rect 17756 2611 17762 2645
rect 17796 2611 17802 2645
rect 17756 2573 17802 2611
rect 17756 2539 17762 2573
rect 17796 2539 17802 2573
rect 17756 2524 17802 2539
rect 17852 3509 17898 3524
rect 17852 3475 17858 3509
rect 17892 3475 17898 3509
rect 17852 3437 17898 3475
rect 17852 3403 17858 3437
rect 17892 3403 17898 3437
rect 17852 3365 17898 3403
rect 17852 3331 17858 3365
rect 17892 3331 17898 3365
rect 17852 3293 17898 3331
rect 17852 3259 17858 3293
rect 17892 3259 17898 3293
rect 17852 3221 17898 3259
rect 17852 3187 17858 3221
rect 17892 3187 17898 3221
rect 17852 3149 17898 3187
rect 17852 3115 17858 3149
rect 17892 3115 17898 3149
rect 17852 3077 17898 3115
rect 17852 3043 17858 3077
rect 17892 3043 17898 3077
rect 17852 3005 17898 3043
rect 17852 2971 17858 3005
rect 17892 2971 17898 3005
rect 17852 2933 17898 2971
rect 17852 2899 17858 2933
rect 17892 2899 17898 2933
rect 17852 2861 17898 2899
rect 17852 2827 17858 2861
rect 17892 2827 17898 2861
rect 17852 2789 17898 2827
rect 17852 2755 17858 2789
rect 17892 2755 17898 2789
rect 17852 2717 17898 2755
rect 17852 2683 17858 2717
rect 17892 2683 17898 2717
rect 17852 2645 17898 2683
rect 17852 2611 17858 2645
rect 17892 2611 17898 2645
rect 17852 2573 17898 2611
rect 17852 2539 17858 2573
rect 17892 2539 17898 2573
rect 17852 2524 17898 2539
rect 17948 3509 17994 3524
rect 17948 3475 17954 3509
rect 17988 3475 17994 3509
rect 17948 3437 17994 3475
rect 17948 3403 17954 3437
rect 17988 3403 17994 3437
rect 17948 3365 17994 3403
rect 17948 3331 17954 3365
rect 17988 3331 17994 3365
rect 17948 3293 17994 3331
rect 17948 3259 17954 3293
rect 17988 3259 17994 3293
rect 17948 3221 17994 3259
rect 17948 3187 17954 3221
rect 17988 3187 17994 3221
rect 17948 3149 17994 3187
rect 17948 3115 17954 3149
rect 17988 3115 17994 3149
rect 17948 3077 17994 3115
rect 17948 3043 17954 3077
rect 17988 3043 17994 3077
rect 17948 3005 17994 3043
rect 17948 2971 17954 3005
rect 17988 2971 17994 3005
rect 17948 2933 17994 2971
rect 17948 2899 17954 2933
rect 17988 2899 17994 2933
rect 17948 2861 17994 2899
rect 17948 2827 17954 2861
rect 17988 2827 17994 2861
rect 17948 2789 17994 2827
rect 17948 2755 17954 2789
rect 17988 2755 17994 2789
rect 17948 2717 17994 2755
rect 17948 2683 17954 2717
rect 17988 2683 17994 2717
rect 17948 2645 17994 2683
rect 17948 2611 17954 2645
rect 17988 2611 17994 2645
rect 17948 2573 17994 2611
rect 17948 2539 17954 2573
rect 17988 2539 17994 2573
rect 17948 2524 17994 2539
rect 18044 3509 18090 3524
rect 18044 3475 18050 3509
rect 18084 3475 18090 3509
rect 18044 3437 18090 3475
rect 18044 3403 18050 3437
rect 18084 3403 18090 3437
rect 18044 3365 18090 3403
rect 18044 3331 18050 3365
rect 18084 3331 18090 3365
rect 18044 3293 18090 3331
rect 18044 3259 18050 3293
rect 18084 3259 18090 3293
rect 18044 3221 18090 3259
rect 18044 3187 18050 3221
rect 18084 3187 18090 3221
rect 18044 3149 18090 3187
rect 18044 3115 18050 3149
rect 18084 3115 18090 3149
rect 18044 3077 18090 3115
rect 18044 3043 18050 3077
rect 18084 3043 18090 3077
rect 18044 3005 18090 3043
rect 18044 2971 18050 3005
rect 18084 2971 18090 3005
rect 18044 2933 18090 2971
rect 18044 2899 18050 2933
rect 18084 2899 18090 2933
rect 18044 2861 18090 2899
rect 18044 2827 18050 2861
rect 18084 2827 18090 2861
rect 18044 2789 18090 2827
rect 18044 2755 18050 2789
rect 18084 2755 18090 2789
rect 18044 2717 18090 2755
rect 18044 2683 18050 2717
rect 18084 2683 18090 2717
rect 18044 2645 18090 2683
rect 18044 2611 18050 2645
rect 18084 2611 18090 2645
rect 18044 2573 18090 2611
rect 18044 2539 18050 2573
rect 18084 2539 18090 2573
rect 18044 2524 18090 2539
rect 18140 3509 18186 3524
rect 18140 3475 18146 3509
rect 18180 3475 18186 3509
rect 18140 3437 18186 3475
rect 18140 3403 18146 3437
rect 18180 3403 18186 3437
rect 18140 3365 18186 3403
rect 18140 3331 18146 3365
rect 18180 3331 18186 3365
rect 18140 3293 18186 3331
rect 18140 3259 18146 3293
rect 18180 3259 18186 3293
rect 18140 3221 18186 3259
rect 18140 3187 18146 3221
rect 18180 3187 18186 3221
rect 18140 3149 18186 3187
rect 18140 3115 18146 3149
rect 18180 3115 18186 3149
rect 18140 3077 18186 3115
rect 18140 3043 18146 3077
rect 18180 3043 18186 3077
rect 18140 3005 18186 3043
rect 18140 2971 18146 3005
rect 18180 2971 18186 3005
rect 18140 2933 18186 2971
rect 18140 2899 18146 2933
rect 18180 2899 18186 2933
rect 18140 2861 18186 2899
rect 18140 2827 18146 2861
rect 18180 2827 18186 2861
rect 18140 2789 18186 2827
rect 18140 2755 18146 2789
rect 18180 2755 18186 2789
rect 18140 2717 18186 2755
rect 18140 2683 18146 2717
rect 18180 2683 18186 2717
rect 18140 2645 18186 2683
rect 18140 2611 18146 2645
rect 18180 2611 18186 2645
rect 18140 2573 18186 2611
rect 18140 2539 18146 2573
rect 18180 2539 18186 2573
rect 18140 2524 18186 2539
rect 18236 3509 18282 3524
rect 18236 3475 18242 3509
rect 18276 3475 18282 3509
rect 18236 3437 18282 3475
rect 18236 3403 18242 3437
rect 18276 3403 18282 3437
rect 18236 3365 18282 3403
rect 18236 3331 18242 3365
rect 18276 3331 18282 3365
rect 18236 3293 18282 3331
rect 18236 3259 18242 3293
rect 18276 3259 18282 3293
rect 18236 3221 18282 3259
rect 18236 3187 18242 3221
rect 18276 3187 18282 3221
rect 18236 3149 18282 3187
rect 18236 3115 18242 3149
rect 18276 3115 18282 3149
rect 18236 3077 18282 3115
rect 18236 3043 18242 3077
rect 18276 3043 18282 3077
rect 18236 3005 18282 3043
rect 18236 2971 18242 3005
rect 18276 2971 18282 3005
rect 18236 2933 18282 2971
rect 18236 2899 18242 2933
rect 18276 2899 18282 2933
rect 18236 2861 18282 2899
rect 18236 2827 18242 2861
rect 18276 2827 18282 2861
rect 18236 2789 18282 2827
rect 18236 2755 18242 2789
rect 18276 2755 18282 2789
rect 18236 2717 18282 2755
rect 18236 2683 18242 2717
rect 18276 2683 18282 2717
rect 18236 2645 18282 2683
rect 18236 2611 18242 2645
rect 18276 2611 18282 2645
rect 18236 2573 18282 2611
rect 18236 2539 18242 2573
rect 18276 2539 18282 2573
rect 18236 2524 18282 2539
rect 18332 3509 18378 3524
rect 18332 3475 18338 3509
rect 18372 3475 18378 3509
rect 18332 3437 18378 3475
rect 18332 3403 18338 3437
rect 18372 3403 18378 3437
rect 18332 3365 18378 3403
rect 18332 3331 18338 3365
rect 18372 3331 18378 3365
rect 18332 3293 18378 3331
rect 18332 3259 18338 3293
rect 18372 3259 18378 3293
rect 18332 3221 18378 3259
rect 18332 3187 18338 3221
rect 18372 3187 18378 3221
rect 18332 3149 18378 3187
rect 18332 3115 18338 3149
rect 18372 3115 18378 3149
rect 18332 3077 18378 3115
rect 18332 3043 18338 3077
rect 18372 3043 18378 3077
rect 18332 3005 18378 3043
rect 18332 2971 18338 3005
rect 18372 2971 18378 3005
rect 18332 2933 18378 2971
rect 18332 2899 18338 2933
rect 18372 2899 18378 2933
rect 18332 2861 18378 2899
rect 18332 2827 18338 2861
rect 18372 2827 18378 2861
rect 18332 2789 18378 2827
rect 18332 2755 18338 2789
rect 18372 2755 18378 2789
rect 18332 2717 18378 2755
rect 18332 2683 18338 2717
rect 18372 2683 18378 2717
rect 18332 2645 18378 2683
rect 18332 2611 18338 2645
rect 18372 2611 18378 2645
rect 18332 2573 18378 2611
rect 18332 2539 18338 2573
rect 18372 2539 18378 2573
rect 18332 2524 18378 2539
rect 18570 3505 18616 3520
rect 18570 3471 18576 3505
rect 18610 3471 18616 3505
rect 18570 3433 18616 3471
rect 18570 3399 18576 3433
rect 18610 3399 18616 3433
rect 18570 3361 18616 3399
rect 18570 3327 18576 3361
rect 18610 3327 18616 3361
rect 18570 3289 18616 3327
rect 18570 3255 18576 3289
rect 18610 3255 18616 3289
rect 18570 3217 18616 3255
rect 18570 3183 18576 3217
rect 18610 3183 18616 3217
rect 18570 3145 18616 3183
rect 18570 3111 18576 3145
rect 18610 3111 18616 3145
rect 18570 3073 18616 3111
rect 18570 3039 18576 3073
rect 18610 3039 18616 3073
rect 18570 3001 18616 3039
rect 18570 2967 18576 3001
rect 18610 2967 18616 3001
rect 18570 2929 18616 2967
rect 18570 2895 18576 2929
rect 18610 2895 18616 2929
rect 18570 2857 18616 2895
rect 18570 2823 18576 2857
rect 18610 2823 18616 2857
rect 18570 2785 18616 2823
rect 18570 2751 18576 2785
rect 18610 2751 18616 2785
rect 18570 2713 18616 2751
rect 18570 2679 18576 2713
rect 18610 2679 18616 2713
rect 18570 2641 18616 2679
rect 18570 2607 18576 2641
rect 18610 2607 18616 2641
rect 18570 2569 18616 2607
rect 18570 2535 18576 2569
rect 18610 2535 18616 2569
rect 18570 2520 18616 2535
rect 18666 3505 18712 3520
rect 18666 3471 18672 3505
rect 18706 3471 18712 3505
rect 18666 3433 18712 3471
rect 18666 3399 18672 3433
rect 18706 3399 18712 3433
rect 18666 3361 18712 3399
rect 18666 3327 18672 3361
rect 18706 3327 18712 3361
rect 18666 3289 18712 3327
rect 18666 3255 18672 3289
rect 18706 3255 18712 3289
rect 18666 3217 18712 3255
rect 18666 3183 18672 3217
rect 18706 3183 18712 3217
rect 18666 3145 18712 3183
rect 18666 3111 18672 3145
rect 18706 3111 18712 3145
rect 18666 3073 18712 3111
rect 18666 3039 18672 3073
rect 18706 3039 18712 3073
rect 18666 3001 18712 3039
rect 18666 2967 18672 3001
rect 18706 2967 18712 3001
rect 18666 2929 18712 2967
rect 18666 2895 18672 2929
rect 18706 2895 18712 2929
rect 18666 2857 18712 2895
rect 18666 2823 18672 2857
rect 18706 2823 18712 2857
rect 18666 2785 18712 2823
rect 18666 2751 18672 2785
rect 18706 2751 18712 2785
rect 18666 2713 18712 2751
rect 18666 2679 18672 2713
rect 18706 2679 18712 2713
rect 18666 2641 18712 2679
rect 18666 2607 18672 2641
rect 18706 2607 18712 2641
rect 18666 2569 18712 2607
rect 18666 2535 18672 2569
rect 18706 2535 18712 2569
rect 18666 2520 18712 2535
rect 18762 3505 18808 3520
rect 18762 3471 18768 3505
rect 18802 3471 18808 3505
rect 18762 3433 18808 3471
rect 18762 3399 18768 3433
rect 18802 3399 18808 3433
rect 18762 3361 18808 3399
rect 18762 3327 18768 3361
rect 18802 3327 18808 3361
rect 18762 3289 18808 3327
rect 18762 3255 18768 3289
rect 18802 3255 18808 3289
rect 18762 3217 18808 3255
rect 18762 3183 18768 3217
rect 18802 3183 18808 3217
rect 18762 3145 18808 3183
rect 18762 3111 18768 3145
rect 18802 3111 18808 3145
rect 18762 3073 18808 3111
rect 18762 3039 18768 3073
rect 18802 3039 18808 3073
rect 18762 3001 18808 3039
rect 18762 2967 18768 3001
rect 18802 2967 18808 3001
rect 18762 2929 18808 2967
rect 18762 2895 18768 2929
rect 18802 2895 18808 2929
rect 18762 2857 18808 2895
rect 18762 2823 18768 2857
rect 18802 2823 18808 2857
rect 18762 2785 18808 2823
rect 18762 2751 18768 2785
rect 18802 2751 18808 2785
rect 18762 2713 18808 2751
rect 18762 2679 18768 2713
rect 18802 2679 18808 2713
rect 18762 2641 18808 2679
rect 18762 2607 18768 2641
rect 18802 2607 18808 2641
rect 18762 2569 18808 2607
rect 18762 2535 18768 2569
rect 18802 2535 18808 2569
rect 18762 2520 18808 2535
rect 18858 3505 18904 3520
rect 18858 3471 18864 3505
rect 18898 3471 18904 3505
rect 18858 3433 18904 3471
rect 18858 3399 18864 3433
rect 18898 3399 18904 3433
rect 18858 3361 18904 3399
rect 18858 3327 18864 3361
rect 18898 3327 18904 3361
rect 18858 3289 18904 3327
rect 18858 3255 18864 3289
rect 18898 3255 18904 3289
rect 18858 3217 18904 3255
rect 18858 3183 18864 3217
rect 18898 3183 18904 3217
rect 18858 3145 18904 3183
rect 18858 3111 18864 3145
rect 18898 3111 18904 3145
rect 18858 3073 18904 3111
rect 18858 3039 18864 3073
rect 18898 3039 18904 3073
rect 18858 3001 18904 3039
rect 18858 2967 18864 3001
rect 18898 2967 18904 3001
rect 18858 2929 18904 2967
rect 18858 2895 18864 2929
rect 18898 2895 18904 2929
rect 18858 2857 18904 2895
rect 18858 2823 18864 2857
rect 18898 2823 18904 2857
rect 18858 2785 18904 2823
rect 18858 2751 18864 2785
rect 18898 2751 18904 2785
rect 18858 2713 18904 2751
rect 18858 2679 18864 2713
rect 18898 2679 18904 2713
rect 18858 2641 18904 2679
rect 18858 2607 18864 2641
rect 18898 2607 18904 2641
rect 18858 2569 18904 2607
rect 18858 2535 18864 2569
rect 18898 2535 18904 2569
rect 18858 2520 18904 2535
rect 18954 3505 19000 3520
rect 18954 3471 18960 3505
rect 18994 3471 19000 3505
rect 18954 3433 19000 3471
rect 18954 3399 18960 3433
rect 18994 3399 19000 3433
rect 18954 3361 19000 3399
rect 18954 3327 18960 3361
rect 18994 3327 19000 3361
rect 18954 3289 19000 3327
rect 18954 3255 18960 3289
rect 18994 3255 19000 3289
rect 18954 3217 19000 3255
rect 18954 3183 18960 3217
rect 18994 3183 19000 3217
rect 18954 3145 19000 3183
rect 18954 3111 18960 3145
rect 18994 3111 19000 3145
rect 18954 3073 19000 3111
rect 18954 3039 18960 3073
rect 18994 3039 19000 3073
rect 18954 3001 19000 3039
rect 18954 2967 18960 3001
rect 18994 2967 19000 3001
rect 18954 2929 19000 2967
rect 18954 2895 18960 2929
rect 18994 2895 19000 2929
rect 18954 2857 19000 2895
rect 18954 2823 18960 2857
rect 18994 2823 19000 2857
rect 18954 2785 19000 2823
rect 18954 2751 18960 2785
rect 18994 2751 19000 2785
rect 18954 2713 19000 2751
rect 18954 2679 18960 2713
rect 18994 2679 19000 2713
rect 18954 2641 19000 2679
rect 18954 2607 18960 2641
rect 18994 2607 19000 2641
rect 18954 2569 19000 2607
rect 18954 2535 18960 2569
rect 18994 2535 19000 2569
rect 18954 2520 19000 2535
rect 19050 3505 19096 3520
rect 19050 3471 19056 3505
rect 19090 3471 19096 3505
rect 19050 3433 19096 3471
rect 19050 3399 19056 3433
rect 19090 3399 19096 3433
rect 19050 3361 19096 3399
rect 19050 3327 19056 3361
rect 19090 3327 19096 3361
rect 19050 3289 19096 3327
rect 19050 3255 19056 3289
rect 19090 3255 19096 3289
rect 19050 3217 19096 3255
rect 19050 3183 19056 3217
rect 19090 3183 19096 3217
rect 19050 3145 19096 3183
rect 19050 3111 19056 3145
rect 19090 3111 19096 3145
rect 19050 3073 19096 3111
rect 19050 3039 19056 3073
rect 19090 3039 19096 3073
rect 19050 3001 19096 3039
rect 19050 2967 19056 3001
rect 19090 2967 19096 3001
rect 19050 2929 19096 2967
rect 19050 2895 19056 2929
rect 19090 2895 19096 2929
rect 19050 2857 19096 2895
rect 19050 2823 19056 2857
rect 19090 2823 19096 2857
rect 19050 2785 19096 2823
rect 19050 2751 19056 2785
rect 19090 2751 19096 2785
rect 19050 2713 19096 2751
rect 19050 2679 19056 2713
rect 19090 2679 19096 2713
rect 19050 2641 19096 2679
rect 19050 2607 19056 2641
rect 19090 2607 19096 2641
rect 19050 2569 19096 2607
rect 19050 2535 19056 2569
rect 19090 2535 19096 2569
rect 19050 2520 19096 2535
rect 19146 3505 19192 3520
rect 19146 3471 19152 3505
rect 19186 3471 19192 3505
rect 19146 3433 19192 3471
rect 19146 3399 19152 3433
rect 19186 3399 19192 3433
rect 19146 3361 19192 3399
rect 19146 3327 19152 3361
rect 19186 3327 19192 3361
rect 19146 3289 19192 3327
rect 19146 3255 19152 3289
rect 19186 3255 19192 3289
rect 19146 3217 19192 3255
rect 19146 3183 19152 3217
rect 19186 3183 19192 3217
rect 19146 3145 19192 3183
rect 19146 3111 19152 3145
rect 19186 3111 19192 3145
rect 19146 3073 19192 3111
rect 19146 3039 19152 3073
rect 19186 3039 19192 3073
rect 19146 3001 19192 3039
rect 19146 2967 19152 3001
rect 19186 2967 19192 3001
rect 19146 2929 19192 2967
rect 19146 2895 19152 2929
rect 19186 2895 19192 2929
rect 19146 2857 19192 2895
rect 19146 2823 19152 2857
rect 19186 2823 19192 2857
rect 19146 2785 19192 2823
rect 19146 2751 19152 2785
rect 19186 2751 19192 2785
rect 19146 2713 19192 2751
rect 19146 2679 19152 2713
rect 19186 2679 19192 2713
rect 19146 2641 19192 2679
rect 19146 2607 19152 2641
rect 19186 2607 19192 2641
rect 19146 2569 19192 2607
rect 19146 2535 19152 2569
rect 19186 2535 19192 2569
rect 19146 2520 19192 2535
rect 19242 3505 19288 3520
rect 19242 3471 19248 3505
rect 19282 3471 19288 3505
rect 19242 3433 19288 3471
rect 19242 3399 19248 3433
rect 19282 3399 19288 3433
rect 19242 3361 19288 3399
rect 19242 3327 19248 3361
rect 19282 3327 19288 3361
rect 19242 3289 19288 3327
rect 19242 3255 19248 3289
rect 19282 3255 19288 3289
rect 19242 3217 19288 3255
rect 19242 3183 19248 3217
rect 19282 3183 19288 3217
rect 19242 3145 19288 3183
rect 19242 3111 19248 3145
rect 19282 3111 19288 3145
rect 19242 3073 19288 3111
rect 19242 3039 19248 3073
rect 19282 3039 19288 3073
rect 19242 3001 19288 3039
rect 19242 2967 19248 3001
rect 19282 2967 19288 3001
rect 19242 2929 19288 2967
rect 19242 2895 19248 2929
rect 19282 2895 19288 2929
rect 19242 2857 19288 2895
rect 19242 2823 19248 2857
rect 19282 2823 19288 2857
rect 19242 2785 19288 2823
rect 19242 2751 19248 2785
rect 19282 2751 19288 2785
rect 19242 2713 19288 2751
rect 19242 2679 19248 2713
rect 19282 2679 19288 2713
rect 19242 2641 19288 2679
rect 19242 2607 19248 2641
rect 19282 2607 19288 2641
rect 19242 2569 19288 2607
rect 19242 2535 19248 2569
rect 19282 2535 19288 2569
rect 19242 2520 19288 2535
rect 19338 3505 19384 3520
rect 19338 3471 19344 3505
rect 19378 3471 19384 3505
rect 19338 3433 19384 3471
rect 19338 3399 19344 3433
rect 19378 3399 19384 3433
rect 19338 3361 19384 3399
rect 19338 3327 19344 3361
rect 19378 3327 19384 3361
rect 19338 3289 19384 3327
rect 19338 3255 19344 3289
rect 19378 3255 19384 3289
rect 19338 3217 19384 3255
rect 19338 3183 19344 3217
rect 19378 3183 19384 3217
rect 19338 3145 19384 3183
rect 19338 3111 19344 3145
rect 19378 3111 19384 3145
rect 19338 3073 19384 3111
rect 19338 3039 19344 3073
rect 19378 3039 19384 3073
rect 19338 3001 19384 3039
rect 19338 2967 19344 3001
rect 19378 2967 19384 3001
rect 19338 2929 19384 2967
rect 19338 2895 19344 2929
rect 19378 2895 19384 2929
rect 19338 2857 19384 2895
rect 19338 2823 19344 2857
rect 19378 2823 19384 2857
rect 19338 2785 19384 2823
rect 19338 2751 19344 2785
rect 19378 2751 19384 2785
rect 19338 2713 19384 2751
rect 19338 2679 19344 2713
rect 19378 2679 19384 2713
rect 19338 2641 19384 2679
rect 19338 2607 19344 2641
rect 19378 2607 19384 2641
rect 19338 2569 19384 2607
rect 19338 2535 19344 2569
rect 19378 2535 19384 2569
rect 19338 2520 19384 2535
rect 19434 3505 19480 3520
rect 19434 3471 19440 3505
rect 19474 3471 19480 3505
rect 19434 3433 19480 3471
rect 19434 3399 19440 3433
rect 19474 3399 19480 3433
rect 19434 3361 19480 3399
rect 19434 3327 19440 3361
rect 19474 3327 19480 3361
rect 19434 3289 19480 3327
rect 19434 3255 19440 3289
rect 19474 3255 19480 3289
rect 19434 3217 19480 3255
rect 19434 3183 19440 3217
rect 19474 3183 19480 3217
rect 19434 3145 19480 3183
rect 19434 3111 19440 3145
rect 19474 3111 19480 3145
rect 19434 3073 19480 3111
rect 19434 3039 19440 3073
rect 19474 3039 19480 3073
rect 19434 3001 19480 3039
rect 19434 2967 19440 3001
rect 19474 2967 19480 3001
rect 19434 2929 19480 2967
rect 19434 2895 19440 2929
rect 19474 2895 19480 2929
rect 19434 2857 19480 2895
rect 19434 2823 19440 2857
rect 19474 2823 19480 2857
rect 19434 2785 19480 2823
rect 19434 2751 19440 2785
rect 19474 2751 19480 2785
rect 19434 2713 19480 2751
rect 19434 2679 19440 2713
rect 19474 2679 19480 2713
rect 19434 2641 19480 2679
rect 19434 2607 19440 2641
rect 19474 2607 19480 2641
rect 19434 2569 19480 2607
rect 19434 2535 19440 2569
rect 19474 2535 19480 2569
rect 19434 2520 19480 2535
rect 19530 3505 19576 3520
rect 19530 3471 19536 3505
rect 19570 3471 19576 3505
rect 19530 3433 19576 3471
rect 19530 3399 19536 3433
rect 19570 3399 19576 3433
rect 19530 3361 19576 3399
rect 19530 3327 19536 3361
rect 19570 3327 19576 3361
rect 19530 3289 19576 3327
rect 19530 3255 19536 3289
rect 19570 3255 19576 3289
rect 19530 3217 19576 3255
rect 19530 3183 19536 3217
rect 19570 3183 19576 3217
rect 19530 3145 19576 3183
rect 19530 3111 19536 3145
rect 19570 3111 19576 3145
rect 19530 3073 19576 3111
rect 19530 3039 19536 3073
rect 19570 3039 19576 3073
rect 19530 3001 19576 3039
rect 19530 2967 19536 3001
rect 19570 2967 19576 3001
rect 19530 2929 19576 2967
rect 19530 2895 19536 2929
rect 19570 2895 19576 2929
rect 19530 2857 19576 2895
rect 19530 2823 19536 2857
rect 19570 2823 19576 2857
rect 19530 2785 19576 2823
rect 19530 2751 19536 2785
rect 19570 2751 19576 2785
rect 19530 2713 19576 2751
rect 19530 2679 19536 2713
rect 19570 2679 19576 2713
rect 19530 2641 19576 2679
rect 19530 2607 19536 2641
rect 19570 2607 19576 2641
rect 19530 2569 19576 2607
rect 19530 2535 19536 2569
rect 19570 2535 19576 2569
rect 19530 2520 19576 2535
rect 19626 3505 19672 3520
rect 19626 3471 19632 3505
rect 19666 3471 19672 3505
rect 19626 3433 19672 3471
rect 19626 3399 19632 3433
rect 19666 3399 19672 3433
rect 19626 3361 19672 3399
rect 19626 3327 19632 3361
rect 19666 3327 19672 3361
rect 19626 3289 19672 3327
rect 19626 3255 19632 3289
rect 19666 3255 19672 3289
rect 19626 3217 19672 3255
rect 19626 3183 19632 3217
rect 19666 3183 19672 3217
rect 19626 3145 19672 3183
rect 19626 3111 19632 3145
rect 19666 3111 19672 3145
rect 19626 3073 19672 3111
rect 19626 3039 19632 3073
rect 19666 3039 19672 3073
rect 19626 3001 19672 3039
rect 19626 2967 19632 3001
rect 19666 2967 19672 3001
rect 19626 2929 19672 2967
rect 19626 2895 19632 2929
rect 19666 2895 19672 2929
rect 19626 2857 19672 2895
rect 19626 2823 19632 2857
rect 19666 2823 19672 2857
rect 19626 2785 19672 2823
rect 19626 2751 19632 2785
rect 19666 2751 19672 2785
rect 19626 2713 19672 2751
rect 19626 2679 19632 2713
rect 19666 2679 19672 2713
rect 19626 2641 19672 2679
rect 19626 2607 19632 2641
rect 19666 2607 19672 2641
rect 19626 2569 19672 2607
rect 19626 2535 19632 2569
rect 19666 2535 19672 2569
rect 19626 2520 19672 2535
rect 19722 3505 19768 3520
rect 19722 3471 19728 3505
rect 19762 3471 19768 3505
rect 19722 3433 19768 3471
rect 19722 3399 19728 3433
rect 19762 3399 19768 3433
rect 19722 3361 19768 3399
rect 19722 3327 19728 3361
rect 19762 3327 19768 3361
rect 19722 3289 19768 3327
rect 19722 3255 19728 3289
rect 19762 3255 19768 3289
rect 19722 3217 19768 3255
rect 19722 3183 19728 3217
rect 19762 3183 19768 3217
rect 19722 3145 19768 3183
rect 19722 3111 19728 3145
rect 19762 3111 19768 3145
rect 19722 3073 19768 3111
rect 19722 3039 19728 3073
rect 19762 3039 19768 3073
rect 19722 3001 19768 3039
rect 19722 2967 19728 3001
rect 19762 2967 19768 3001
rect 19722 2929 19768 2967
rect 19722 2895 19728 2929
rect 19762 2895 19768 2929
rect 19722 2857 19768 2895
rect 19722 2823 19728 2857
rect 19762 2823 19768 2857
rect 19722 2785 19768 2823
rect 19722 2751 19728 2785
rect 19762 2751 19768 2785
rect 19722 2713 19768 2751
rect 19722 2679 19728 2713
rect 19762 2679 19768 2713
rect 19722 2641 19768 2679
rect 19722 2607 19728 2641
rect 19762 2607 19768 2641
rect 19722 2569 19768 2607
rect 19722 2535 19728 2569
rect 19762 2535 19768 2569
rect 19722 2520 19768 2535
rect 19818 3505 19864 3520
rect 19818 3471 19824 3505
rect 19858 3471 19864 3505
rect 19818 3433 19864 3471
rect 19818 3399 19824 3433
rect 19858 3399 19864 3433
rect 19818 3361 19864 3399
rect 19818 3327 19824 3361
rect 19858 3327 19864 3361
rect 19818 3289 19864 3327
rect 19818 3255 19824 3289
rect 19858 3255 19864 3289
rect 19818 3217 19864 3255
rect 19818 3183 19824 3217
rect 19858 3183 19864 3217
rect 19818 3145 19864 3183
rect 19818 3111 19824 3145
rect 19858 3111 19864 3145
rect 19818 3073 19864 3111
rect 19818 3039 19824 3073
rect 19858 3039 19864 3073
rect 19818 3001 19864 3039
rect 19818 2967 19824 3001
rect 19858 2967 19864 3001
rect 19818 2929 19864 2967
rect 19818 2895 19824 2929
rect 19858 2895 19864 2929
rect 19818 2857 19864 2895
rect 19818 2823 19824 2857
rect 19858 2823 19864 2857
rect 19818 2785 19864 2823
rect 19818 2751 19824 2785
rect 19858 2751 19864 2785
rect 19818 2713 19864 2751
rect 19818 2679 19824 2713
rect 19858 2679 19864 2713
rect 19818 2641 19864 2679
rect 19818 2607 19824 2641
rect 19858 2607 19864 2641
rect 19818 2569 19864 2607
rect 19818 2535 19824 2569
rect 19858 2535 19864 2569
rect 19818 2520 19864 2535
rect 19914 3505 19960 3520
rect 19914 3471 19920 3505
rect 19954 3471 19960 3505
rect 19914 3433 19960 3471
rect 19914 3399 19920 3433
rect 19954 3399 19960 3433
rect 19914 3361 19960 3399
rect 19914 3327 19920 3361
rect 19954 3327 19960 3361
rect 19914 3289 19960 3327
rect 19914 3255 19920 3289
rect 19954 3255 19960 3289
rect 19914 3217 19960 3255
rect 19914 3183 19920 3217
rect 19954 3183 19960 3217
rect 19914 3145 19960 3183
rect 19914 3111 19920 3145
rect 19954 3111 19960 3145
rect 19914 3073 19960 3111
rect 19914 3039 19920 3073
rect 19954 3039 19960 3073
rect 19914 3001 19960 3039
rect 19914 2967 19920 3001
rect 19954 2967 19960 3001
rect 19914 2929 19960 2967
rect 19914 2895 19920 2929
rect 19954 2895 19960 2929
rect 19914 2857 19960 2895
rect 19914 2823 19920 2857
rect 19954 2823 19960 2857
rect 19914 2785 19960 2823
rect 19914 2751 19920 2785
rect 19954 2751 19960 2785
rect 19914 2713 19960 2751
rect 19914 2679 19920 2713
rect 19954 2679 19960 2713
rect 19914 2641 19960 2679
rect 19914 2607 19920 2641
rect 19954 2607 19960 2641
rect 19914 2569 19960 2607
rect 19914 2535 19920 2569
rect 19954 2535 19960 2569
rect 19914 2520 19960 2535
rect 20010 3505 20056 3520
rect 20010 3471 20016 3505
rect 20050 3471 20056 3505
rect 20010 3433 20056 3471
rect 20010 3399 20016 3433
rect 20050 3399 20056 3433
rect 20010 3361 20056 3399
rect 20010 3327 20016 3361
rect 20050 3327 20056 3361
rect 20010 3289 20056 3327
rect 20010 3255 20016 3289
rect 20050 3255 20056 3289
rect 20010 3217 20056 3255
rect 20010 3183 20016 3217
rect 20050 3183 20056 3217
rect 20010 3145 20056 3183
rect 20010 3111 20016 3145
rect 20050 3111 20056 3145
rect 20010 3073 20056 3111
rect 20010 3039 20016 3073
rect 20050 3039 20056 3073
rect 20010 3001 20056 3039
rect 20010 2967 20016 3001
rect 20050 2967 20056 3001
rect 20010 2929 20056 2967
rect 20010 2895 20016 2929
rect 20050 2895 20056 2929
rect 20010 2857 20056 2895
rect 20010 2823 20016 2857
rect 20050 2823 20056 2857
rect 20010 2785 20056 2823
rect 20010 2751 20016 2785
rect 20050 2751 20056 2785
rect 20010 2713 20056 2751
rect 20010 2679 20016 2713
rect 20050 2679 20056 2713
rect 20010 2641 20056 2679
rect 20010 2607 20016 2641
rect 20050 2607 20056 2641
rect 20010 2569 20056 2607
rect 20010 2535 20016 2569
rect 20050 2535 20056 2569
rect 20010 2520 20056 2535
rect 20238 3513 20284 3528
rect 20238 3479 20244 3513
rect 20278 3479 20284 3513
rect 20238 3441 20284 3479
rect 20238 3407 20244 3441
rect 20278 3407 20284 3441
rect 20238 3369 20284 3407
rect 20238 3335 20244 3369
rect 20278 3335 20284 3369
rect 20238 3297 20284 3335
rect 20238 3263 20244 3297
rect 20278 3263 20284 3297
rect 20238 3225 20284 3263
rect 20238 3191 20244 3225
rect 20278 3191 20284 3225
rect 20238 3153 20284 3191
rect 20238 3119 20244 3153
rect 20278 3119 20284 3153
rect 20238 3081 20284 3119
rect 20238 3047 20244 3081
rect 20278 3047 20284 3081
rect 20238 3009 20284 3047
rect 20238 2975 20244 3009
rect 20278 2975 20284 3009
rect 20238 2937 20284 2975
rect 20238 2903 20244 2937
rect 20278 2903 20284 2937
rect 20238 2865 20284 2903
rect 20238 2831 20244 2865
rect 20278 2831 20284 2865
rect 20238 2793 20284 2831
rect 20238 2759 20244 2793
rect 20278 2759 20284 2793
rect 20238 2721 20284 2759
rect 20238 2687 20244 2721
rect 20278 2687 20284 2721
rect 20238 2649 20284 2687
rect 20238 2615 20244 2649
rect 20278 2615 20284 2649
rect 20238 2577 20284 2615
rect 20238 2543 20244 2577
rect 20278 2543 20284 2577
rect 20238 2528 20284 2543
rect 20334 3513 20380 3528
rect 20334 3479 20340 3513
rect 20374 3479 20380 3513
rect 20334 3441 20380 3479
rect 20334 3407 20340 3441
rect 20374 3407 20380 3441
rect 20334 3369 20380 3407
rect 20334 3335 20340 3369
rect 20374 3335 20380 3369
rect 20334 3297 20380 3335
rect 20334 3263 20340 3297
rect 20374 3263 20380 3297
rect 20334 3225 20380 3263
rect 20334 3191 20340 3225
rect 20374 3191 20380 3225
rect 20334 3153 20380 3191
rect 20334 3119 20340 3153
rect 20374 3119 20380 3153
rect 20334 3081 20380 3119
rect 20334 3047 20340 3081
rect 20374 3047 20380 3081
rect 20334 3009 20380 3047
rect 20334 2975 20340 3009
rect 20374 2975 20380 3009
rect 20334 2937 20380 2975
rect 20334 2903 20340 2937
rect 20374 2903 20380 2937
rect 20334 2865 20380 2903
rect 20334 2831 20340 2865
rect 20374 2831 20380 2865
rect 20334 2793 20380 2831
rect 20334 2759 20340 2793
rect 20374 2759 20380 2793
rect 20334 2721 20380 2759
rect 20334 2687 20340 2721
rect 20374 2687 20380 2721
rect 20334 2649 20380 2687
rect 20334 2615 20340 2649
rect 20374 2615 20380 2649
rect 20334 2577 20380 2615
rect 20334 2543 20340 2577
rect 20374 2543 20380 2577
rect 20334 2528 20380 2543
rect 20430 3513 20476 3528
rect 20430 3479 20436 3513
rect 20470 3479 20476 3513
rect 20430 3441 20476 3479
rect 20430 3407 20436 3441
rect 20470 3407 20476 3441
rect 20430 3369 20476 3407
rect 20430 3335 20436 3369
rect 20470 3335 20476 3369
rect 20430 3297 20476 3335
rect 20430 3263 20436 3297
rect 20470 3263 20476 3297
rect 20430 3225 20476 3263
rect 20430 3191 20436 3225
rect 20470 3191 20476 3225
rect 20430 3153 20476 3191
rect 20430 3119 20436 3153
rect 20470 3119 20476 3153
rect 20430 3081 20476 3119
rect 20430 3047 20436 3081
rect 20470 3047 20476 3081
rect 20430 3009 20476 3047
rect 20430 2975 20436 3009
rect 20470 2975 20476 3009
rect 20430 2937 20476 2975
rect 20430 2903 20436 2937
rect 20470 2903 20476 2937
rect 20430 2865 20476 2903
rect 20430 2831 20436 2865
rect 20470 2831 20476 2865
rect 20430 2793 20476 2831
rect 20430 2759 20436 2793
rect 20470 2759 20476 2793
rect 20430 2721 20476 2759
rect 20430 2687 20436 2721
rect 20470 2687 20476 2721
rect 20430 2649 20476 2687
rect 20430 2615 20436 2649
rect 20470 2615 20476 2649
rect 20430 2577 20476 2615
rect 20430 2543 20436 2577
rect 20470 2543 20476 2577
rect 20430 2528 20476 2543
rect 20526 3513 20572 3528
rect 20526 3479 20532 3513
rect 20566 3479 20572 3513
rect 20526 3441 20572 3479
rect 20526 3407 20532 3441
rect 20566 3407 20572 3441
rect 20526 3369 20572 3407
rect 20526 3335 20532 3369
rect 20566 3335 20572 3369
rect 20526 3297 20572 3335
rect 20526 3263 20532 3297
rect 20566 3263 20572 3297
rect 20526 3225 20572 3263
rect 20526 3191 20532 3225
rect 20566 3191 20572 3225
rect 20526 3153 20572 3191
rect 20526 3119 20532 3153
rect 20566 3119 20572 3153
rect 20526 3081 20572 3119
rect 20526 3047 20532 3081
rect 20566 3047 20572 3081
rect 20526 3009 20572 3047
rect 20526 2975 20532 3009
rect 20566 2975 20572 3009
rect 20526 2937 20572 2975
rect 20526 2903 20532 2937
rect 20566 2903 20572 2937
rect 20526 2865 20572 2903
rect 20526 2831 20532 2865
rect 20566 2831 20572 2865
rect 20526 2793 20572 2831
rect 20526 2759 20532 2793
rect 20566 2759 20572 2793
rect 20526 2721 20572 2759
rect 20526 2687 20532 2721
rect 20566 2687 20572 2721
rect 20526 2649 20572 2687
rect 20526 2615 20532 2649
rect 20566 2615 20572 2649
rect 20526 2577 20572 2615
rect 20526 2543 20532 2577
rect 20566 2543 20572 2577
rect 20526 2528 20572 2543
rect 20622 3513 20668 3528
rect 20622 3479 20628 3513
rect 20662 3479 20668 3513
rect 20622 3441 20668 3479
rect 20622 3407 20628 3441
rect 20662 3407 20668 3441
rect 20622 3369 20668 3407
rect 20622 3335 20628 3369
rect 20662 3335 20668 3369
rect 20622 3297 20668 3335
rect 20622 3263 20628 3297
rect 20662 3263 20668 3297
rect 20622 3225 20668 3263
rect 20622 3191 20628 3225
rect 20662 3191 20668 3225
rect 20622 3153 20668 3191
rect 20622 3119 20628 3153
rect 20662 3119 20668 3153
rect 20622 3081 20668 3119
rect 20622 3047 20628 3081
rect 20662 3047 20668 3081
rect 20622 3009 20668 3047
rect 20622 2975 20628 3009
rect 20662 2975 20668 3009
rect 20622 2937 20668 2975
rect 20622 2903 20628 2937
rect 20662 2903 20668 2937
rect 20622 2865 20668 2903
rect 20622 2831 20628 2865
rect 20662 2831 20668 2865
rect 20622 2793 20668 2831
rect 20622 2759 20628 2793
rect 20662 2759 20668 2793
rect 20622 2721 20668 2759
rect 20622 2687 20628 2721
rect 20662 2687 20668 2721
rect 20622 2649 20668 2687
rect 20622 2615 20628 2649
rect 20662 2615 20668 2649
rect 20622 2577 20668 2615
rect 20622 2543 20628 2577
rect 20662 2543 20668 2577
rect 20622 2528 20668 2543
rect 20718 3513 20764 3528
rect 20718 3479 20724 3513
rect 20758 3479 20764 3513
rect 20718 3441 20764 3479
rect 20718 3407 20724 3441
rect 20758 3407 20764 3441
rect 20718 3369 20764 3407
rect 20718 3335 20724 3369
rect 20758 3335 20764 3369
rect 20718 3297 20764 3335
rect 20718 3263 20724 3297
rect 20758 3263 20764 3297
rect 20718 3225 20764 3263
rect 20718 3191 20724 3225
rect 20758 3191 20764 3225
rect 20718 3153 20764 3191
rect 20718 3119 20724 3153
rect 20758 3119 20764 3153
rect 20718 3081 20764 3119
rect 20718 3047 20724 3081
rect 20758 3047 20764 3081
rect 20718 3009 20764 3047
rect 20718 2975 20724 3009
rect 20758 2975 20764 3009
rect 20718 2937 20764 2975
rect 20718 2903 20724 2937
rect 20758 2903 20764 2937
rect 20718 2865 20764 2903
rect 20718 2831 20724 2865
rect 20758 2831 20764 2865
rect 20718 2793 20764 2831
rect 20718 2759 20724 2793
rect 20758 2759 20764 2793
rect 20718 2721 20764 2759
rect 20718 2687 20724 2721
rect 20758 2687 20764 2721
rect 20718 2649 20764 2687
rect 20718 2615 20724 2649
rect 20758 2615 20764 2649
rect 20718 2577 20764 2615
rect 20718 2543 20724 2577
rect 20758 2543 20764 2577
rect 20718 2528 20764 2543
rect 20814 3513 20860 3528
rect 20814 3479 20820 3513
rect 20854 3479 20860 3513
rect 20814 3441 20860 3479
rect 20814 3407 20820 3441
rect 20854 3407 20860 3441
rect 20814 3369 20860 3407
rect 20814 3335 20820 3369
rect 20854 3335 20860 3369
rect 20814 3297 20860 3335
rect 20814 3263 20820 3297
rect 20854 3263 20860 3297
rect 20814 3225 20860 3263
rect 20814 3191 20820 3225
rect 20854 3191 20860 3225
rect 20814 3153 20860 3191
rect 20814 3119 20820 3153
rect 20854 3119 20860 3153
rect 20814 3081 20860 3119
rect 20814 3047 20820 3081
rect 20854 3047 20860 3081
rect 20814 3009 20860 3047
rect 20814 2975 20820 3009
rect 20854 2975 20860 3009
rect 20814 2937 20860 2975
rect 20814 2903 20820 2937
rect 20854 2903 20860 2937
rect 20814 2865 20860 2903
rect 20814 2831 20820 2865
rect 20854 2831 20860 2865
rect 20814 2793 20860 2831
rect 20814 2759 20820 2793
rect 20854 2759 20860 2793
rect 20814 2721 20860 2759
rect 20814 2687 20820 2721
rect 20854 2687 20860 2721
rect 20814 2649 20860 2687
rect 20814 2615 20820 2649
rect 20854 2615 20860 2649
rect 20814 2577 20860 2615
rect 20814 2543 20820 2577
rect 20854 2543 20860 2577
rect 20814 2528 20860 2543
rect 20910 3513 20956 3528
rect 20910 3479 20916 3513
rect 20950 3479 20956 3513
rect 20910 3441 20956 3479
rect 20910 3407 20916 3441
rect 20950 3407 20956 3441
rect 20910 3369 20956 3407
rect 20910 3335 20916 3369
rect 20950 3335 20956 3369
rect 20910 3297 20956 3335
rect 20910 3263 20916 3297
rect 20950 3263 20956 3297
rect 20910 3225 20956 3263
rect 20910 3191 20916 3225
rect 20950 3191 20956 3225
rect 20910 3153 20956 3191
rect 20910 3119 20916 3153
rect 20950 3119 20956 3153
rect 20910 3081 20956 3119
rect 20910 3047 20916 3081
rect 20950 3047 20956 3081
rect 20910 3009 20956 3047
rect 20910 2975 20916 3009
rect 20950 2975 20956 3009
rect 20910 2937 20956 2975
rect 20910 2903 20916 2937
rect 20950 2903 20956 2937
rect 20910 2865 20956 2903
rect 20910 2831 20916 2865
rect 20950 2831 20956 2865
rect 20910 2793 20956 2831
rect 20910 2759 20916 2793
rect 20950 2759 20956 2793
rect 20910 2721 20956 2759
rect 20910 2687 20916 2721
rect 20950 2687 20956 2721
rect 20910 2649 20956 2687
rect 20910 2615 20916 2649
rect 20950 2615 20956 2649
rect 20910 2577 20956 2615
rect 20910 2543 20916 2577
rect 20950 2543 20956 2577
rect 20910 2528 20956 2543
rect 21006 3513 21052 3528
rect 21006 3479 21012 3513
rect 21046 3479 21052 3513
rect 21006 3441 21052 3479
rect 21006 3407 21012 3441
rect 21046 3407 21052 3441
rect 21006 3369 21052 3407
rect 21006 3335 21012 3369
rect 21046 3335 21052 3369
rect 21006 3297 21052 3335
rect 21006 3263 21012 3297
rect 21046 3263 21052 3297
rect 21006 3225 21052 3263
rect 21006 3191 21012 3225
rect 21046 3191 21052 3225
rect 21006 3153 21052 3191
rect 21006 3119 21012 3153
rect 21046 3119 21052 3153
rect 21006 3081 21052 3119
rect 21006 3047 21012 3081
rect 21046 3047 21052 3081
rect 21006 3009 21052 3047
rect 21006 2975 21012 3009
rect 21046 2975 21052 3009
rect 21006 2937 21052 2975
rect 21006 2903 21012 2937
rect 21046 2903 21052 2937
rect 21006 2865 21052 2903
rect 21006 2831 21012 2865
rect 21046 2831 21052 2865
rect 21006 2793 21052 2831
rect 21006 2759 21012 2793
rect 21046 2759 21052 2793
rect 21006 2721 21052 2759
rect 21006 2687 21012 2721
rect 21046 2687 21052 2721
rect 21006 2649 21052 2687
rect 21006 2615 21012 2649
rect 21046 2615 21052 2649
rect 21006 2577 21052 2615
rect 21006 2543 21012 2577
rect 21046 2543 21052 2577
rect 21006 2528 21052 2543
rect 21102 3513 21148 3528
rect 21102 3479 21108 3513
rect 21142 3479 21148 3513
rect 21102 3441 21148 3479
rect 21102 3407 21108 3441
rect 21142 3407 21148 3441
rect 21102 3369 21148 3407
rect 21102 3335 21108 3369
rect 21142 3335 21148 3369
rect 21102 3297 21148 3335
rect 21102 3263 21108 3297
rect 21142 3263 21148 3297
rect 21102 3225 21148 3263
rect 21102 3191 21108 3225
rect 21142 3191 21148 3225
rect 21102 3153 21148 3191
rect 21102 3119 21108 3153
rect 21142 3119 21148 3153
rect 21102 3081 21148 3119
rect 21102 3047 21108 3081
rect 21142 3047 21148 3081
rect 21102 3009 21148 3047
rect 21102 2975 21108 3009
rect 21142 2975 21148 3009
rect 21102 2937 21148 2975
rect 21102 2903 21108 2937
rect 21142 2903 21148 2937
rect 21102 2865 21148 2903
rect 21102 2831 21108 2865
rect 21142 2831 21148 2865
rect 21102 2793 21148 2831
rect 21102 2759 21108 2793
rect 21142 2759 21148 2793
rect 21102 2721 21148 2759
rect 21102 2687 21108 2721
rect 21142 2687 21148 2721
rect 21102 2649 21148 2687
rect 21102 2615 21108 2649
rect 21142 2615 21148 2649
rect 21102 2577 21148 2615
rect 21102 2543 21108 2577
rect 21142 2543 21148 2577
rect 21102 2528 21148 2543
rect 21198 3513 21244 3528
rect 21198 3479 21204 3513
rect 21238 3479 21244 3513
rect 21198 3441 21244 3479
rect 21198 3407 21204 3441
rect 21238 3407 21244 3441
rect 21198 3369 21244 3407
rect 21198 3335 21204 3369
rect 21238 3335 21244 3369
rect 21198 3297 21244 3335
rect 21198 3263 21204 3297
rect 21238 3263 21244 3297
rect 21198 3225 21244 3263
rect 21198 3191 21204 3225
rect 21238 3191 21244 3225
rect 21198 3153 21244 3191
rect 21198 3119 21204 3153
rect 21238 3119 21244 3153
rect 21198 3081 21244 3119
rect 21198 3047 21204 3081
rect 21238 3047 21244 3081
rect 21198 3009 21244 3047
rect 21198 2975 21204 3009
rect 21238 2975 21244 3009
rect 21198 2937 21244 2975
rect 21198 2903 21204 2937
rect 21238 2903 21244 2937
rect 21198 2865 21244 2903
rect 21198 2831 21204 2865
rect 21238 2831 21244 2865
rect 21198 2793 21244 2831
rect 21198 2759 21204 2793
rect 21238 2759 21244 2793
rect 21198 2721 21244 2759
rect 21198 2687 21204 2721
rect 21238 2687 21244 2721
rect 21198 2649 21244 2687
rect 21198 2615 21204 2649
rect 21238 2615 21244 2649
rect 21198 2577 21244 2615
rect 21198 2543 21204 2577
rect 21238 2543 21244 2577
rect 21198 2528 21244 2543
rect 21294 3513 21340 3528
rect 21294 3479 21300 3513
rect 21334 3479 21340 3513
rect 21294 3441 21340 3479
rect 21294 3407 21300 3441
rect 21334 3407 21340 3441
rect 21294 3369 21340 3407
rect 21294 3335 21300 3369
rect 21334 3335 21340 3369
rect 21294 3297 21340 3335
rect 21294 3263 21300 3297
rect 21334 3263 21340 3297
rect 21294 3225 21340 3263
rect 21294 3191 21300 3225
rect 21334 3191 21340 3225
rect 21294 3153 21340 3191
rect 21294 3119 21300 3153
rect 21334 3119 21340 3153
rect 21294 3081 21340 3119
rect 21294 3047 21300 3081
rect 21334 3047 21340 3081
rect 21294 3009 21340 3047
rect 21294 2975 21300 3009
rect 21334 2975 21340 3009
rect 21294 2937 21340 2975
rect 21294 2903 21300 2937
rect 21334 2903 21340 2937
rect 21294 2865 21340 2903
rect 21294 2831 21300 2865
rect 21334 2831 21340 2865
rect 21294 2793 21340 2831
rect 21294 2759 21300 2793
rect 21334 2759 21340 2793
rect 21294 2721 21340 2759
rect 21294 2687 21300 2721
rect 21334 2687 21340 2721
rect 21294 2649 21340 2687
rect 21294 2615 21300 2649
rect 21334 2615 21340 2649
rect 21294 2577 21340 2615
rect 21294 2543 21300 2577
rect 21334 2543 21340 2577
rect 21294 2528 21340 2543
rect 21390 3513 21436 3528
rect 21390 3479 21396 3513
rect 21430 3479 21436 3513
rect 21390 3441 21436 3479
rect 21390 3407 21396 3441
rect 21430 3407 21436 3441
rect 21390 3369 21436 3407
rect 21390 3335 21396 3369
rect 21430 3335 21436 3369
rect 21390 3297 21436 3335
rect 21390 3263 21396 3297
rect 21430 3263 21436 3297
rect 21390 3225 21436 3263
rect 21390 3191 21396 3225
rect 21430 3191 21436 3225
rect 21390 3153 21436 3191
rect 21390 3119 21396 3153
rect 21430 3119 21436 3153
rect 21390 3081 21436 3119
rect 21390 3047 21396 3081
rect 21430 3047 21436 3081
rect 21390 3009 21436 3047
rect 21390 2975 21396 3009
rect 21430 2975 21436 3009
rect 21390 2937 21436 2975
rect 21390 2903 21396 2937
rect 21430 2903 21436 2937
rect 21390 2865 21436 2903
rect 21390 2831 21396 2865
rect 21430 2831 21436 2865
rect 21390 2793 21436 2831
rect 21390 2759 21396 2793
rect 21430 2759 21436 2793
rect 21390 2721 21436 2759
rect 21390 2687 21396 2721
rect 21430 2687 21436 2721
rect 21390 2649 21436 2687
rect 21390 2615 21396 2649
rect 21430 2615 21436 2649
rect 21390 2577 21436 2615
rect 21390 2543 21396 2577
rect 21430 2543 21436 2577
rect 21390 2528 21436 2543
rect 21486 3513 21532 3528
rect 21486 3479 21492 3513
rect 21526 3479 21532 3513
rect 21486 3441 21532 3479
rect 21486 3407 21492 3441
rect 21526 3407 21532 3441
rect 21486 3369 21532 3407
rect 21486 3335 21492 3369
rect 21526 3335 21532 3369
rect 21486 3297 21532 3335
rect 21486 3263 21492 3297
rect 21526 3263 21532 3297
rect 21486 3225 21532 3263
rect 21486 3191 21492 3225
rect 21526 3191 21532 3225
rect 21486 3153 21532 3191
rect 21486 3119 21492 3153
rect 21526 3119 21532 3153
rect 21486 3081 21532 3119
rect 21486 3047 21492 3081
rect 21526 3047 21532 3081
rect 21486 3009 21532 3047
rect 21486 2975 21492 3009
rect 21526 2975 21532 3009
rect 21486 2937 21532 2975
rect 21486 2903 21492 2937
rect 21526 2903 21532 2937
rect 21486 2865 21532 2903
rect 21486 2831 21492 2865
rect 21526 2831 21532 2865
rect 21486 2793 21532 2831
rect 21486 2759 21492 2793
rect 21526 2759 21532 2793
rect 21486 2721 21532 2759
rect 21486 2687 21492 2721
rect 21526 2687 21532 2721
rect 21486 2649 21532 2687
rect 21486 2615 21492 2649
rect 21526 2615 21532 2649
rect 21486 2577 21532 2615
rect 21486 2543 21492 2577
rect 21526 2543 21532 2577
rect 21486 2528 21532 2543
rect 21582 3513 21628 3528
rect 21582 3479 21588 3513
rect 21622 3479 21628 3513
rect 21582 3441 21628 3479
rect 21582 3407 21588 3441
rect 21622 3407 21628 3441
rect 21582 3369 21628 3407
rect 21582 3335 21588 3369
rect 21622 3335 21628 3369
rect 21582 3297 21628 3335
rect 21582 3263 21588 3297
rect 21622 3263 21628 3297
rect 21582 3225 21628 3263
rect 21582 3191 21588 3225
rect 21622 3191 21628 3225
rect 21582 3153 21628 3191
rect 21582 3119 21588 3153
rect 21622 3119 21628 3153
rect 21582 3081 21628 3119
rect 21582 3047 21588 3081
rect 21622 3047 21628 3081
rect 21582 3009 21628 3047
rect 21582 2975 21588 3009
rect 21622 2975 21628 3009
rect 21582 2937 21628 2975
rect 21582 2903 21588 2937
rect 21622 2903 21628 2937
rect 21582 2865 21628 2903
rect 21582 2831 21588 2865
rect 21622 2831 21628 2865
rect 21582 2793 21628 2831
rect 21582 2759 21588 2793
rect 21622 2759 21628 2793
rect 21582 2721 21628 2759
rect 21582 2687 21588 2721
rect 21622 2687 21628 2721
rect 21582 2649 21628 2687
rect 21582 2615 21588 2649
rect 21622 2615 21628 2649
rect 21582 2577 21628 2615
rect 21582 2543 21588 2577
rect 21622 2543 21628 2577
rect 21582 2528 21628 2543
rect 21678 3513 21724 3528
rect 21678 3479 21684 3513
rect 21718 3479 21724 3513
rect 21678 3441 21724 3479
rect 21678 3407 21684 3441
rect 21718 3407 21724 3441
rect 21678 3369 21724 3407
rect 21678 3335 21684 3369
rect 21718 3335 21724 3369
rect 21678 3297 21724 3335
rect 21678 3263 21684 3297
rect 21718 3263 21724 3297
rect 21678 3225 21724 3263
rect 21678 3191 21684 3225
rect 21718 3191 21724 3225
rect 21678 3153 21724 3191
rect 21678 3119 21684 3153
rect 21718 3119 21724 3153
rect 21678 3081 21724 3119
rect 21678 3047 21684 3081
rect 21718 3047 21724 3081
rect 21678 3009 21724 3047
rect 21678 2975 21684 3009
rect 21718 2975 21724 3009
rect 21678 2937 21724 2975
rect 21678 2903 21684 2937
rect 21718 2903 21724 2937
rect 21678 2865 21724 2903
rect 21678 2831 21684 2865
rect 21718 2831 21724 2865
rect 21678 2793 21724 2831
rect 21678 2759 21684 2793
rect 21718 2759 21724 2793
rect 21678 2721 21724 2759
rect 21678 2687 21684 2721
rect 21718 2687 21724 2721
rect 21678 2649 21724 2687
rect 21678 2615 21684 2649
rect 21718 2615 21724 2649
rect 21678 2577 21724 2615
rect 21678 2543 21684 2577
rect 21718 2543 21724 2577
rect 21678 2528 21724 2543
rect 21774 3513 21820 3528
rect 21774 3479 21780 3513
rect 21814 3479 21820 3513
rect 21774 3441 21820 3479
rect 21774 3407 21780 3441
rect 21814 3407 21820 3441
rect 21774 3369 21820 3407
rect 21774 3335 21780 3369
rect 21814 3335 21820 3369
rect 21774 3297 21820 3335
rect 21774 3263 21780 3297
rect 21814 3263 21820 3297
rect 21774 3225 21820 3263
rect 21774 3191 21780 3225
rect 21814 3191 21820 3225
rect 21774 3153 21820 3191
rect 21774 3119 21780 3153
rect 21814 3119 21820 3153
rect 21774 3081 21820 3119
rect 21774 3047 21780 3081
rect 21814 3047 21820 3081
rect 21774 3009 21820 3047
rect 21774 2975 21780 3009
rect 21814 2975 21820 3009
rect 21774 2937 21820 2975
rect 21774 2903 21780 2937
rect 21814 2903 21820 2937
rect 21774 2865 21820 2903
rect 21774 2831 21780 2865
rect 21814 2831 21820 2865
rect 21774 2793 21820 2831
rect 21774 2759 21780 2793
rect 21814 2759 21820 2793
rect 21774 2721 21820 2759
rect 21774 2687 21780 2721
rect 21814 2687 21820 2721
rect 21774 2649 21820 2687
rect 21774 2615 21780 2649
rect 21814 2615 21820 2649
rect 21774 2577 21820 2615
rect 21774 2543 21780 2577
rect 21814 2543 21820 2577
rect 21774 2528 21820 2543
rect 21870 3513 21916 3528
rect 21870 3479 21876 3513
rect 21910 3479 21916 3513
rect 21870 3441 21916 3479
rect 21870 3407 21876 3441
rect 21910 3407 21916 3441
rect 21870 3369 21916 3407
rect 21870 3335 21876 3369
rect 21910 3335 21916 3369
rect 21870 3297 21916 3335
rect 21870 3263 21876 3297
rect 21910 3263 21916 3297
rect 21870 3225 21916 3263
rect 21870 3191 21876 3225
rect 21910 3191 21916 3225
rect 21870 3153 21916 3191
rect 21870 3119 21876 3153
rect 21910 3119 21916 3153
rect 21870 3081 21916 3119
rect 21870 3047 21876 3081
rect 21910 3047 21916 3081
rect 21870 3009 21916 3047
rect 21870 2975 21876 3009
rect 21910 2975 21916 3009
rect 21870 2937 21916 2975
rect 21870 2903 21876 2937
rect 21910 2903 21916 2937
rect 21870 2865 21916 2903
rect 21870 2831 21876 2865
rect 21910 2831 21916 2865
rect 21870 2793 21916 2831
rect 21870 2759 21876 2793
rect 21910 2759 21916 2793
rect 21870 2721 21916 2759
rect 21870 2687 21876 2721
rect 21910 2687 21916 2721
rect 21870 2649 21916 2687
rect 21870 2615 21876 2649
rect 21910 2615 21916 2649
rect 21870 2577 21916 2615
rect 21870 2543 21876 2577
rect 21910 2543 21916 2577
rect 21870 2528 21916 2543
rect 21966 3513 22012 3528
rect 21966 3479 21972 3513
rect 22006 3479 22012 3513
rect 21966 3441 22012 3479
rect 21966 3407 21972 3441
rect 22006 3407 22012 3441
rect 21966 3369 22012 3407
rect 21966 3335 21972 3369
rect 22006 3335 22012 3369
rect 21966 3297 22012 3335
rect 21966 3263 21972 3297
rect 22006 3263 22012 3297
rect 21966 3225 22012 3263
rect 21966 3191 21972 3225
rect 22006 3191 22012 3225
rect 21966 3153 22012 3191
rect 21966 3119 21972 3153
rect 22006 3119 22012 3153
rect 21966 3081 22012 3119
rect 21966 3047 21972 3081
rect 22006 3047 22012 3081
rect 21966 3009 22012 3047
rect 21966 2975 21972 3009
rect 22006 2975 22012 3009
rect 21966 2937 22012 2975
rect 21966 2903 21972 2937
rect 22006 2903 22012 2937
rect 21966 2865 22012 2903
rect 21966 2831 21972 2865
rect 22006 2831 22012 2865
rect 21966 2793 22012 2831
rect 21966 2759 21972 2793
rect 22006 2759 22012 2793
rect 21966 2721 22012 2759
rect 21966 2687 21972 2721
rect 22006 2687 22012 2721
rect 21966 2649 22012 2687
rect 21966 2615 21972 2649
rect 22006 2615 22012 2649
rect 21966 2577 22012 2615
rect 21966 2543 21972 2577
rect 22006 2543 22012 2577
rect 21966 2528 22012 2543
rect 22062 3513 22108 3528
rect 22062 3479 22068 3513
rect 22102 3479 22108 3513
rect 22062 3441 22108 3479
rect 22062 3407 22068 3441
rect 22102 3407 22108 3441
rect 22062 3369 22108 3407
rect 22062 3335 22068 3369
rect 22102 3335 22108 3369
rect 22062 3297 22108 3335
rect 22062 3263 22068 3297
rect 22102 3263 22108 3297
rect 22062 3225 22108 3263
rect 22062 3191 22068 3225
rect 22102 3191 22108 3225
rect 22062 3153 22108 3191
rect 22062 3119 22068 3153
rect 22102 3119 22108 3153
rect 22062 3081 22108 3119
rect 22062 3047 22068 3081
rect 22102 3047 22108 3081
rect 22062 3009 22108 3047
rect 22062 2975 22068 3009
rect 22102 2975 22108 3009
rect 22062 2937 22108 2975
rect 22062 2903 22068 2937
rect 22102 2903 22108 2937
rect 22062 2865 22108 2903
rect 22062 2831 22068 2865
rect 22102 2831 22108 2865
rect 22062 2793 22108 2831
rect 22062 2759 22068 2793
rect 22102 2759 22108 2793
rect 22062 2721 22108 2759
rect 22062 2687 22068 2721
rect 22102 2687 22108 2721
rect 22062 2649 22108 2687
rect 22062 2615 22068 2649
rect 22102 2615 22108 2649
rect 22062 2577 22108 2615
rect 22062 2543 22068 2577
rect 22102 2543 22108 2577
rect 22062 2528 22108 2543
rect 22158 3513 22204 3528
rect 22158 3479 22164 3513
rect 22198 3479 22204 3513
rect 22158 3441 22204 3479
rect 22158 3407 22164 3441
rect 22198 3407 22204 3441
rect 22158 3369 22204 3407
rect 22158 3335 22164 3369
rect 22198 3335 22204 3369
rect 22158 3297 22204 3335
rect 22158 3263 22164 3297
rect 22198 3263 22204 3297
rect 22158 3225 22204 3263
rect 22158 3191 22164 3225
rect 22198 3191 22204 3225
rect 22158 3153 22204 3191
rect 22158 3119 22164 3153
rect 22198 3119 22204 3153
rect 22158 3081 22204 3119
rect 22158 3047 22164 3081
rect 22198 3047 22204 3081
rect 22158 3009 22204 3047
rect 22158 2975 22164 3009
rect 22198 2975 22204 3009
rect 22158 2937 22204 2975
rect 22158 2903 22164 2937
rect 22198 2903 22204 2937
rect 22158 2865 22204 2903
rect 22158 2831 22164 2865
rect 22198 2831 22204 2865
rect 22158 2793 22204 2831
rect 22158 2759 22164 2793
rect 22198 2759 22204 2793
rect 22158 2721 22204 2759
rect 22158 2687 22164 2721
rect 22198 2687 22204 2721
rect 22158 2649 22204 2687
rect 22158 2615 22164 2649
rect 22198 2615 22204 2649
rect 22158 2577 22204 2615
rect 22158 2543 22164 2577
rect 22198 2543 22204 2577
rect 22158 2528 22204 2543
rect 17892 2339 18190 2342
rect 17892 2159 17919 2339
rect 18163 2159 18190 2339
rect 17892 2156 18190 2159
rect 19892 2339 20190 2342
rect 19892 2159 19919 2339
rect 20163 2159 20190 2339
rect 19892 2156 20190 2159
rect 21890 2339 22190 2342
rect 21890 2159 21918 2339
rect 22162 2159 22190 2339
rect 21890 2156 22190 2159
rect 15320 -320 15760 -258
rect 15320 -400 15384 -320
rect 2794 -446 15384 -400
rect 2794 -460 11751 -446
rect 2794 -462 5639 -460
rect 2794 -514 2889 -462
rect 2941 -512 5639 -462
rect 5691 -512 8677 -460
rect 8729 -498 11751 -460
rect 11803 -498 15384 -446
rect 8729 -512 15384 -498
rect 2941 -514 15384 -512
rect 2794 -570 15384 -514
rect 246 -962 706 -948
rect 246 -1270 258 -962
rect 694 -1270 706 -962
rect 246 -1284 706 -1270
rect 15400 -960 15772 -944
rect 15400 -1268 15432 -960
rect 15740 -1268 15772 -960
rect 15400 -1284 15772 -1268
rect 2218 -1465 2496 -1452
rect 2218 -1468 2269 -1465
rect 2447 -1468 2496 -1465
rect 2218 -1648 2235 -1468
rect 2479 -1648 2496 -1468
rect 2218 -1664 2496 -1648
rect 4218 -1465 4496 -1452
rect 4218 -1468 4269 -1465
rect 4447 -1468 4496 -1465
rect 4218 -1648 4235 -1468
rect 4479 -1648 4496 -1468
rect 4218 -1664 4496 -1648
rect 6218 -1465 6496 -1452
rect 6218 -1468 6269 -1465
rect 6447 -1468 6496 -1465
rect 6218 -1648 6235 -1468
rect 6479 -1648 6496 -1468
rect 6218 -1664 6496 -1648
rect 8436 -1482 8732 -1464
rect 8436 -1493 8493 -1482
rect 8671 -1493 8732 -1482
rect 8436 -1673 8462 -1493
rect 8706 -1673 8732 -1493
rect 10218 -1465 10496 -1452
rect 10218 -1468 10269 -1465
rect 10447 -1468 10496 -1465
rect 10218 -1648 10235 -1468
rect 10479 -1648 10496 -1468
rect 10218 -1664 10496 -1648
rect 12218 -1465 12496 -1452
rect 12218 -1468 12269 -1465
rect 12447 -1468 12496 -1465
rect 12218 -1648 12235 -1468
rect 12479 -1648 12496 -1468
rect 12218 -1664 12496 -1648
rect 14218 -1465 14496 -1452
rect 14218 -1468 14269 -1465
rect 14447 -1468 14496 -1465
rect 14218 -1648 14235 -1468
rect 14479 -1648 14496 -1468
rect 14218 -1664 14496 -1648
rect 8436 -1702 8732 -1673
rect 22450 -5144 22722 3752
rect 22948 3818 23382 3844
rect 23986 3959 24066 3990
rect 23986 3925 24006 3959
rect 24040 3925 24066 3959
rect 23986 3838 24066 3925
rect 25176 3953 25276 3984
rect 25176 3919 25210 3953
rect 25244 3919 25276 3953
rect 25176 3848 25276 3919
rect 24224 3844 25276 3848
rect 22948 3766 22981 3818
rect 23033 3766 23382 3818
rect 23434 3819 24066 3838
rect 23434 3785 23462 3819
rect 23496 3785 24066 3819
rect 23434 3768 24066 3785
rect 22948 3740 23382 3766
rect 23284 3704 23382 3740
rect 23284 3670 23318 3704
rect 23352 3670 23382 3704
rect 23986 3734 24066 3768
rect 24138 3817 25276 3844
rect 26836 3947 26948 3992
rect 26836 3913 26874 3947
rect 26908 3913 26948 3947
rect 26836 3830 26948 3913
rect 24138 3783 24278 3817
rect 24312 3783 25276 3817
rect 24138 3752 25276 3783
rect 24138 3740 24252 3752
rect 23986 3700 24010 3734
rect 24044 3700 24066 3734
rect 23986 3678 24066 3700
rect 25176 3690 25276 3752
rect 25878 3804 26948 3830
rect 25878 3770 25931 3804
rect 25965 3770 26948 3804
rect 25878 3746 26948 3770
rect 28078 3802 29438 3822
rect 28078 3768 28134 3802
rect 28168 3768 29438 3802
rect 28078 3750 29438 3768
rect 23284 3644 23382 3670
rect 25176 3656 25208 3690
rect 25242 3656 25276 3690
rect 25176 3630 25276 3656
rect 26836 3688 26948 3746
rect 26836 3654 26876 3688
rect 26910 3654 26948 3688
rect 26836 3614 26948 3654
rect 23168 3517 23214 3532
rect 23168 3483 23174 3517
rect 23208 3483 23214 3517
rect 23168 3445 23214 3483
rect 23168 3411 23174 3445
rect 23208 3411 23214 3445
rect 23168 3373 23214 3411
rect 23168 3339 23174 3373
rect 23208 3339 23214 3373
rect 23168 3301 23214 3339
rect 23168 3267 23174 3301
rect 23208 3267 23214 3301
rect 23168 3229 23214 3267
rect 23168 3195 23174 3229
rect 23208 3195 23214 3229
rect 23168 3157 23214 3195
rect 23168 3123 23174 3157
rect 23208 3123 23214 3157
rect 23168 3085 23214 3123
rect 23168 3051 23174 3085
rect 23208 3051 23214 3085
rect 23168 3013 23214 3051
rect 23168 2979 23174 3013
rect 23208 2979 23214 3013
rect 23168 2941 23214 2979
rect 23168 2907 23174 2941
rect 23208 2907 23214 2941
rect 23168 2869 23214 2907
rect 23168 2835 23174 2869
rect 23208 2835 23214 2869
rect 23168 2797 23214 2835
rect 23168 2763 23174 2797
rect 23208 2763 23214 2797
rect 23168 2725 23214 2763
rect 23168 2691 23174 2725
rect 23208 2691 23214 2725
rect 23168 2653 23214 2691
rect 23168 2619 23174 2653
rect 23208 2619 23214 2653
rect 23168 2581 23214 2619
rect 23168 2547 23174 2581
rect 23208 2547 23214 2581
rect 23168 2532 23214 2547
rect 23264 3517 23310 3532
rect 23264 3483 23270 3517
rect 23304 3483 23310 3517
rect 23264 3445 23310 3483
rect 23264 3411 23270 3445
rect 23304 3411 23310 3445
rect 23264 3373 23310 3411
rect 23264 3339 23270 3373
rect 23304 3339 23310 3373
rect 23264 3301 23310 3339
rect 23264 3267 23270 3301
rect 23304 3267 23310 3301
rect 23264 3229 23310 3267
rect 23264 3195 23270 3229
rect 23304 3195 23310 3229
rect 23264 3157 23310 3195
rect 23264 3123 23270 3157
rect 23304 3123 23310 3157
rect 23264 3085 23310 3123
rect 23264 3051 23270 3085
rect 23304 3051 23310 3085
rect 23264 3013 23310 3051
rect 23264 2979 23270 3013
rect 23304 2979 23310 3013
rect 23264 2941 23310 2979
rect 23264 2907 23270 2941
rect 23304 2907 23310 2941
rect 23264 2869 23310 2907
rect 23264 2835 23270 2869
rect 23304 2835 23310 2869
rect 23264 2797 23310 2835
rect 23264 2763 23270 2797
rect 23304 2763 23310 2797
rect 23264 2725 23310 2763
rect 23264 2691 23270 2725
rect 23304 2691 23310 2725
rect 23264 2653 23310 2691
rect 23264 2619 23270 2653
rect 23304 2619 23310 2653
rect 23264 2581 23310 2619
rect 23264 2547 23270 2581
rect 23304 2547 23310 2581
rect 23264 2532 23310 2547
rect 23360 3517 23406 3532
rect 23360 3483 23366 3517
rect 23400 3483 23406 3517
rect 23360 3445 23406 3483
rect 23360 3411 23366 3445
rect 23400 3411 23406 3445
rect 23360 3373 23406 3411
rect 23360 3339 23366 3373
rect 23400 3339 23406 3373
rect 23360 3301 23406 3339
rect 23360 3267 23366 3301
rect 23400 3267 23406 3301
rect 23360 3229 23406 3267
rect 23360 3195 23366 3229
rect 23400 3195 23406 3229
rect 23360 3157 23406 3195
rect 23360 3123 23366 3157
rect 23400 3123 23406 3157
rect 23360 3085 23406 3123
rect 23360 3051 23366 3085
rect 23400 3051 23406 3085
rect 23360 3013 23406 3051
rect 23360 2979 23366 3013
rect 23400 2979 23406 3013
rect 23360 2941 23406 2979
rect 23360 2907 23366 2941
rect 23400 2907 23406 2941
rect 23360 2869 23406 2907
rect 23360 2835 23366 2869
rect 23400 2835 23406 2869
rect 23360 2797 23406 2835
rect 23360 2763 23366 2797
rect 23400 2763 23406 2797
rect 23360 2725 23406 2763
rect 23360 2691 23366 2725
rect 23400 2691 23406 2725
rect 23360 2653 23406 2691
rect 23360 2619 23366 2653
rect 23400 2619 23406 2653
rect 23360 2581 23406 2619
rect 23360 2547 23366 2581
rect 23400 2547 23406 2581
rect 23360 2532 23406 2547
rect 23456 3517 23502 3532
rect 23456 3483 23462 3517
rect 23496 3483 23502 3517
rect 23456 3445 23502 3483
rect 23456 3411 23462 3445
rect 23496 3411 23502 3445
rect 23456 3373 23502 3411
rect 23456 3339 23462 3373
rect 23496 3339 23502 3373
rect 23456 3301 23502 3339
rect 23456 3267 23462 3301
rect 23496 3267 23502 3301
rect 23456 3229 23502 3267
rect 23456 3195 23462 3229
rect 23496 3195 23502 3229
rect 23456 3157 23502 3195
rect 23456 3123 23462 3157
rect 23496 3123 23502 3157
rect 23456 3085 23502 3123
rect 23456 3051 23462 3085
rect 23496 3051 23502 3085
rect 23456 3013 23502 3051
rect 23456 2979 23462 3013
rect 23496 2979 23502 3013
rect 23456 2941 23502 2979
rect 23456 2907 23462 2941
rect 23496 2907 23502 2941
rect 23456 2869 23502 2907
rect 23456 2835 23462 2869
rect 23496 2835 23502 2869
rect 23456 2797 23502 2835
rect 23456 2763 23462 2797
rect 23496 2763 23502 2797
rect 23456 2725 23502 2763
rect 23456 2691 23462 2725
rect 23496 2691 23502 2725
rect 23456 2653 23502 2691
rect 23456 2619 23462 2653
rect 23496 2619 23502 2653
rect 23456 2581 23502 2619
rect 23456 2547 23462 2581
rect 23496 2547 23502 2581
rect 23456 2532 23502 2547
rect 23552 3517 23598 3532
rect 23552 3483 23558 3517
rect 23592 3483 23598 3517
rect 23552 3445 23598 3483
rect 23552 3411 23558 3445
rect 23592 3411 23598 3445
rect 23552 3373 23598 3411
rect 23552 3339 23558 3373
rect 23592 3339 23598 3373
rect 23552 3301 23598 3339
rect 23552 3267 23558 3301
rect 23592 3267 23598 3301
rect 23552 3229 23598 3267
rect 23552 3195 23558 3229
rect 23592 3195 23598 3229
rect 23552 3157 23598 3195
rect 23552 3123 23558 3157
rect 23592 3123 23598 3157
rect 23552 3085 23598 3123
rect 23552 3051 23558 3085
rect 23592 3051 23598 3085
rect 23552 3013 23598 3051
rect 23552 2979 23558 3013
rect 23592 2979 23598 3013
rect 23552 2941 23598 2979
rect 23552 2907 23558 2941
rect 23592 2907 23598 2941
rect 23552 2869 23598 2907
rect 23552 2835 23558 2869
rect 23592 2835 23598 2869
rect 23552 2797 23598 2835
rect 23552 2763 23558 2797
rect 23592 2763 23598 2797
rect 23552 2725 23598 2763
rect 23552 2691 23558 2725
rect 23592 2691 23598 2725
rect 23552 2653 23598 2691
rect 23552 2619 23558 2653
rect 23592 2619 23598 2653
rect 23552 2581 23598 2619
rect 23552 2547 23558 2581
rect 23592 2547 23598 2581
rect 23552 2532 23598 2547
rect 23648 3517 23694 3532
rect 23648 3483 23654 3517
rect 23688 3483 23694 3517
rect 23648 3445 23694 3483
rect 23648 3411 23654 3445
rect 23688 3411 23694 3445
rect 23648 3373 23694 3411
rect 23648 3339 23654 3373
rect 23688 3339 23694 3373
rect 23648 3301 23694 3339
rect 23648 3267 23654 3301
rect 23688 3267 23694 3301
rect 23648 3229 23694 3267
rect 23648 3195 23654 3229
rect 23688 3195 23694 3229
rect 23648 3157 23694 3195
rect 23648 3123 23654 3157
rect 23688 3123 23694 3157
rect 23648 3085 23694 3123
rect 23648 3051 23654 3085
rect 23688 3051 23694 3085
rect 23648 3013 23694 3051
rect 23648 2979 23654 3013
rect 23688 2979 23694 3013
rect 23648 2941 23694 2979
rect 23648 2907 23654 2941
rect 23688 2907 23694 2941
rect 23648 2869 23694 2907
rect 23648 2835 23654 2869
rect 23688 2835 23694 2869
rect 23648 2797 23694 2835
rect 23648 2763 23654 2797
rect 23688 2763 23694 2797
rect 23648 2725 23694 2763
rect 23648 2691 23654 2725
rect 23688 2691 23694 2725
rect 23648 2653 23694 2691
rect 23648 2619 23654 2653
rect 23688 2619 23694 2653
rect 23648 2581 23694 2619
rect 23648 2547 23654 2581
rect 23688 2547 23694 2581
rect 23648 2532 23694 2547
rect 23860 3507 23906 3522
rect 23860 3473 23866 3507
rect 23900 3473 23906 3507
rect 23860 3435 23906 3473
rect 23860 3401 23866 3435
rect 23900 3401 23906 3435
rect 23860 3363 23906 3401
rect 23860 3329 23866 3363
rect 23900 3329 23906 3363
rect 23860 3291 23906 3329
rect 23860 3257 23866 3291
rect 23900 3257 23906 3291
rect 23860 3219 23906 3257
rect 23860 3185 23866 3219
rect 23900 3185 23906 3219
rect 23860 3147 23906 3185
rect 23860 3113 23866 3147
rect 23900 3113 23906 3147
rect 23860 3075 23906 3113
rect 23860 3041 23866 3075
rect 23900 3041 23906 3075
rect 23860 3003 23906 3041
rect 23860 2969 23866 3003
rect 23900 2969 23906 3003
rect 23860 2931 23906 2969
rect 23860 2897 23866 2931
rect 23900 2897 23906 2931
rect 23860 2859 23906 2897
rect 23860 2825 23866 2859
rect 23900 2825 23906 2859
rect 23860 2787 23906 2825
rect 23860 2753 23866 2787
rect 23900 2753 23906 2787
rect 23860 2715 23906 2753
rect 23860 2681 23866 2715
rect 23900 2681 23906 2715
rect 23860 2643 23906 2681
rect 23860 2609 23866 2643
rect 23900 2609 23906 2643
rect 23860 2571 23906 2609
rect 23860 2537 23866 2571
rect 23900 2537 23906 2571
rect 23860 2522 23906 2537
rect 23956 3507 24002 3522
rect 23956 3473 23962 3507
rect 23996 3473 24002 3507
rect 23956 3435 24002 3473
rect 23956 3401 23962 3435
rect 23996 3401 24002 3435
rect 23956 3363 24002 3401
rect 23956 3329 23962 3363
rect 23996 3329 24002 3363
rect 23956 3291 24002 3329
rect 23956 3257 23962 3291
rect 23996 3257 24002 3291
rect 23956 3219 24002 3257
rect 23956 3185 23962 3219
rect 23996 3185 24002 3219
rect 23956 3147 24002 3185
rect 23956 3113 23962 3147
rect 23996 3113 24002 3147
rect 23956 3075 24002 3113
rect 23956 3041 23962 3075
rect 23996 3041 24002 3075
rect 23956 3003 24002 3041
rect 23956 2969 23962 3003
rect 23996 2969 24002 3003
rect 23956 2931 24002 2969
rect 23956 2897 23962 2931
rect 23996 2897 24002 2931
rect 23956 2859 24002 2897
rect 23956 2825 23962 2859
rect 23996 2825 24002 2859
rect 23956 2787 24002 2825
rect 23956 2753 23962 2787
rect 23996 2753 24002 2787
rect 23956 2715 24002 2753
rect 23956 2681 23962 2715
rect 23996 2681 24002 2715
rect 23956 2643 24002 2681
rect 23956 2609 23962 2643
rect 23996 2609 24002 2643
rect 23956 2571 24002 2609
rect 23956 2537 23962 2571
rect 23996 2537 24002 2571
rect 23956 2522 24002 2537
rect 24052 3507 24098 3522
rect 24052 3473 24058 3507
rect 24092 3473 24098 3507
rect 24052 3435 24098 3473
rect 24052 3401 24058 3435
rect 24092 3401 24098 3435
rect 24052 3363 24098 3401
rect 24052 3329 24058 3363
rect 24092 3329 24098 3363
rect 24052 3291 24098 3329
rect 24052 3257 24058 3291
rect 24092 3257 24098 3291
rect 24052 3219 24098 3257
rect 24052 3185 24058 3219
rect 24092 3185 24098 3219
rect 24052 3147 24098 3185
rect 24052 3113 24058 3147
rect 24092 3113 24098 3147
rect 24052 3075 24098 3113
rect 24052 3041 24058 3075
rect 24092 3041 24098 3075
rect 24052 3003 24098 3041
rect 24052 2969 24058 3003
rect 24092 2969 24098 3003
rect 24052 2931 24098 2969
rect 24052 2897 24058 2931
rect 24092 2897 24098 2931
rect 24052 2859 24098 2897
rect 24052 2825 24058 2859
rect 24092 2825 24098 2859
rect 24052 2787 24098 2825
rect 24052 2753 24058 2787
rect 24092 2753 24098 2787
rect 24052 2715 24098 2753
rect 24052 2681 24058 2715
rect 24092 2681 24098 2715
rect 24052 2643 24098 2681
rect 24052 2609 24058 2643
rect 24092 2609 24098 2643
rect 24052 2571 24098 2609
rect 24052 2537 24058 2571
rect 24092 2537 24098 2571
rect 24052 2522 24098 2537
rect 24148 3507 24194 3522
rect 24148 3473 24154 3507
rect 24188 3473 24194 3507
rect 24148 3435 24194 3473
rect 24148 3401 24154 3435
rect 24188 3401 24194 3435
rect 24148 3363 24194 3401
rect 24148 3329 24154 3363
rect 24188 3329 24194 3363
rect 24148 3291 24194 3329
rect 24148 3257 24154 3291
rect 24188 3257 24194 3291
rect 24148 3219 24194 3257
rect 24148 3185 24154 3219
rect 24188 3185 24194 3219
rect 24148 3147 24194 3185
rect 24148 3113 24154 3147
rect 24188 3113 24194 3147
rect 24148 3075 24194 3113
rect 24148 3041 24154 3075
rect 24188 3041 24194 3075
rect 24148 3003 24194 3041
rect 24148 2969 24154 3003
rect 24188 2969 24194 3003
rect 24148 2931 24194 2969
rect 24148 2897 24154 2931
rect 24188 2897 24194 2931
rect 24148 2859 24194 2897
rect 24148 2825 24154 2859
rect 24188 2825 24194 2859
rect 24148 2787 24194 2825
rect 24148 2753 24154 2787
rect 24188 2753 24194 2787
rect 24148 2715 24194 2753
rect 24148 2681 24154 2715
rect 24188 2681 24194 2715
rect 24148 2643 24194 2681
rect 24148 2609 24154 2643
rect 24188 2609 24194 2643
rect 24148 2571 24194 2609
rect 24148 2537 24154 2571
rect 24188 2537 24194 2571
rect 24148 2522 24194 2537
rect 24244 3507 24290 3522
rect 24244 3473 24250 3507
rect 24284 3473 24290 3507
rect 24244 3435 24290 3473
rect 24244 3401 24250 3435
rect 24284 3401 24290 3435
rect 24244 3363 24290 3401
rect 24244 3329 24250 3363
rect 24284 3329 24290 3363
rect 24244 3291 24290 3329
rect 24244 3257 24250 3291
rect 24284 3257 24290 3291
rect 24244 3219 24290 3257
rect 24244 3185 24250 3219
rect 24284 3185 24290 3219
rect 24244 3147 24290 3185
rect 24244 3113 24250 3147
rect 24284 3113 24290 3147
rect 24244 3075 24290 3113
rect 24244 3041 24250 3075
rect 24284 3041 24290 3075
rect 24244 3003 24290 3041
rect 24244 2969 24250 3003
rect 24284 2969 24290 3003
rect 24244 2931 24290 2969
rect 24244 2897 24250 2931
rect 24284 2897 24290 2931
rect 24244 2859 24290 2897
rect 24244 2825 24250 2859
rect 24284 2825 24290 2859
rect 24244 2787 24290 2825
rect 24244 2753 24250 2787
rect 24284 2753 24290 2787
rect 24244 2715 24290 2753
rect 24244 2681 24250 2715
rect 24284 2681 24290 2715
rect 24244 2643 24290 2681
rect 24244 2609 24250 2643
rect 24284 2609 24290 2643
rect 24244 2571 24290 2609
rect 24244 2537 24250 2571
rect 24284 2537 24290 2571
rect 24244 2522 24290 2537
rect 24340 3507 24386 3522
rect 24340 3473 24346 3507
rect 24380 3473 24386 3507
rect 24340 3435 24386 3473
rect 24340 3401 24346 3435
rect 24380 3401 24386 3435
rect 24340 3363 24386 3401
rect 24340 3329 24346 3363
rect 24380 3329 24386 3363
rect 24340 3291 24386 3329
rect 24340 3257 24346 3291
rect 24380 3257 24386 3291
rect 24340 3219 24386 3257
rect 24340 3185 24346 3219
rect 24380 3185 24386 3219
rect 24340 3147 24386 3185
rect 24340 3113 24346 3147
rect 24380 3113 24386 3147
rect 24340 3075 24386 3113
rect 24340 3041 24346 3075
rect 24380 3041 24386 3075
rect 24340 3003 24386 3041
rect 24340 2969 24346 3003
rect 24380 2969 24386 3003
rect 24340 2931 24386 2969
rect 24340 2897 24346 2931
rect 24380 2897 24386 2931
rect 24340 2859 24386 2897
rect 24340 2825 24346 2859
rect 24380 2825 24386 2859
rect 24340 2787 24386 2825
rect 24340 2753 24346 2787
rect 24380 2753 24386 2787
rect 24340 2715 24386 2753
rect 24340 2681 24346 2715
rect 24380 2681 24386 2715
rect 24340 2643 24386 2681
rect 24340 2609 24346 2643
rect 24380 2609 24386 2643
rect 24340 2571 24386 2609
rect 24340 2537 24346 2571
rect 24380 2537 24386 2571
rect 24340 2522 24386 2537
rect 24436 3507 24482 3522
rect 24436 3473 24442 3507
rect 24476 3473 24482 3507
rect 24436 3435 24482 3473
rect 24436 3401 24442 3435
rect 24476 3401 24482 3435
rect 24436 3363 24482 3401
rect 24436 3329 24442 3363
rect 24476 3329 24482 3363
rect 24436 3291 24482 3329
rect 24436 3257 24442 3291
rect 24476 3257 24482 3291
rect 24436 3219 24482 3257
rect 24436 3185 24442 3219
rect 24476 3185 24482 3219
rect 24436 3147 24482 3185
rect 24436 3113 24442 3147
rect 24476 3113 24482 3147
rect 24436 3075 24482 3113
rect 24436 3041 24442 3075
rect 24476 3041 24482 3075
rect 24436 3003 24482 3041
rect 24436 2969 24442 3003
rect 24476 2969 24482 3003
rect 24436 2931 24482 2969
rect 24436 2897 24442 2931
rect 24476 2897 24482 2931
rect 24436 2859 24482 2897
rect 24436 2825 24442 2859
rect 24476 2825 24482 2859
rect 24436 2787 24482 2825
rect 24436 2753 24442 2787
rect 24476 2753 24482 2787
rect 24436 2715 24482 2753
rect 24436 2681 24442 2715
rect 24476 2681 24482 2715
rect 24436 2643 24482 2681
rect 24436 2609 24442 2643
rect 24476 2609 24482 2643
rect 24436 2571 24482 2609
rect 24436 2537 24442 2571
rect 24476 2537 24482 2571
rect 24436 2522 24482 2537
rect 24532 3507 24578 3522
rect 24532 3473 24538 3507
rect 24572 3473 24578 3507
rect 24532 3435 24578 3473
rect 24532 3401 24538 3435
rect 24572 3401 24578 3435
rect 24532 3363 24578 3401
rect 24532 3329 24538 3363
rect 24572 3329 24578 3363
rect 24532 3291 24578 3329
rect 24532 3257 24538 3291
rect 24572 3257 24578 3291
rect 24532 3219 24578 3257
rect 24532 3185 24538 3219
rect 24572 3185 24578 3219
rect 24532 3147 24578 3185
rect 24532 3113 24538 3147
rect 24572 3113 24578 3147
rect 24532 3075 24578 3113
rect 24532 3041 24538 3075
rect 24572 3041 24578 3075
rect 24532 3003 24578 3041
rect 24532 2969 24538 3003
rect 24572 2969 24578 3003
rect 24532 2931 24578 2969
rect 24532 2897 24538 2931
rect 24572 2897 24578 2931
rect 24532 2859 24578 2897
rect 24532 2825 24538 2859
rect 24572 2825 24578 2859
rect 24532 2787 24578 2825
rect 24532 2753 24538 2787
rect 24572 2753 24578 2787
rect 24532 2715 24578 2753
rect 24532 2681 24538 2715
rect 24572 2681 24578 2715
rect 24532 2643 24578 2681
rect 24532 2609 24538 2643
rect 24572 2609 24578 2643
rect 24532 2571 24578 2609
rect 24532 2537 24538 2571
rect 24572 2537 24578 2571
rect 24532 2522 24578 2537
rect 24628 3507 24674 3522
rect 24628 3473 24634 3507
rect 24668 3473 24674 3507
rect 24628 3435 24674 3473
rect 24628 3401 24634 3435
rect 24668 3401 24674 3435
rect 24628 3363 24674 3401
rect 24628 3329 24634 3363
rect 24668 3329 24674 3363
rect 24628 3291 24674 3329
rect 24628 3257 24634 3291
rect 24668 3257 24674 3291
rect 24628 3219 24674 3257
rect 24628 3185 24634 3219
rect 24668 3185 24674 3219
rect 24628 3147 24674 3185
rect 24628 3113 24634 3147
rect 24668 3113 24674 3147
rect 24628 3075 24674 3113
rect 24628 3041 24634 3075
rect 24668 3041 24674 3075
rect 24628 3003 24674 3041
rect 24628 2969 24634 3003
rect 24668 2969 24674 3003
rect 24628 2931 24674 2969
rect 24628 2897 24634 2931
rect 24668 2897 24674 2931
rect 24628 2859 24674 2897
rect 24628 2825 24634 2859
rect 24668 2825 24674 2859
rect 24628 2787 24674 2825
rect 24628 2753 24634 2787
rect 24668 2753 24674 2787
rect 24628 2715 24674 2753
rect 24628 2681 24634 2715
rect 24668 2681 24674 2715
rect 24628 2643 24674 2681
rect 24628 2609 24634 2643
rect 24668 2609 24674 2643
rect 24628 2571 24674 2609
rect 24628 2537 24634 2571
rect 24668 2537 24674 2571
rect 24628 2522 24674 2537
rect 24724 3507 24770 3522
rect 24724 3473 24730 3507
rect 24764 3473 24770 3507
rect 24724 3435 24770 3473
rect 24724 3401 24730 3435
rect 24764 3401 24770 3435
rect 24724 3363 24770 3401
rect 24724 3329 24730 3363
rect 24764 3329 24770 3363
rect 24724 3291 24770 3329
rect 24724 3257 24730 3291
rect 24764 3257 24770 3291
rect 24724 3219 24770 3257
rect 24724 3185 24730 3219
rect 24764 3185 24770 3219
rect 24724 3147 24770 3185
rect 24724 3113 24730 3147
rect 24764 3113 24770 3147
rect 24724 3075 24770 3113
rect 24724 3041 24730 3075
rect 24764 3041 24770 3075
rect 24724 3003 24770 3041
rect 24724 2969 24730 3003
rect 24764 2969 24770 3003
rect 24724 2931 24770 2969
rect 24724 2897 24730 2931
rect 24764 2897 24770 2931
rect 24724 2859 24770 2897
rect 24724 2825 24730 2859
rect 24764 2825 24770 2859
rect 24724 2787 24770 2825
rect 24724 2753 24730 2787
rect 24764 2753 24770 2787
rect 24724 2715 24770 2753
rect 24724 2681 24730 2715
rect 24764 2681 24770 2715
rect 24724 2643 24770 2681
rect 24724 2609 24730 2643
rect 24764 2609 24770 2643
rect 24724 2571 24770 2609
rect 24724 2537 24730 2571
rect 24764 2537 24770 2571
rect 24724 2522 24770 2537
rect 24820 3507 24866 3522
rect 24820 3473 24826 3507
rect 24860 3473 24866 3507
rect 24820 3435 24866 3473
rect 24820 3401 24826 3435
rect 24860 3401 24866 3435
rect 24820 3363 24866 3401
rect 24820 3329 24826 3363
rect 24860 3329 24866 3363
rect 24820 3291 24866 3329
rect 24820 3257 24826 3291
rect 24860 3257 24866 3291
rect 24820 3219 24866 3257
rect 24820 3185 24826 3219
rect 24860 3185 24866 3219
rect 24820 3147 24866 3185
rect 24820 3113 24826 3147
rect 24860 3113 24866 3147
rect 24820 3075 24866 3113
rect 24820 3041 24826 3075
rect 24860 3041 24866 3075
rect 24820 3003 24866 3041
rect 24820 2969 24826 3003
rect 24860 2969 24866 3003
rect 24820 2931 24866 2969
rect 24820 2897 24826 2931
rect 24860 2897 24866 2931
rect 24820 2859 24866 2897
rect 24820 2825 24826 2859
rect 24860 2825 24866 2859
rect 24820 2787 24866 2825
rect 24820 2753 24826 2787
rect 24860 2753 24866 2787
rect 24820 2715 24866 2753
rect 24820 2681 24826 2715
rect 24860 2681 24866 2715
rect 24820 2643 24866 2681
rect 24820 2609 24826 2643
rect 24860 2609 24866 2643
rect 24820 2571 24866 2609
rect 24820 2537 24826 2571
rect 24860 2537 24866 2571
rect 24820 2522 24866 2537
rect 25058 3503 25104 3518
rect 25058 3469 25064 3503
rect 25098 3469 25104 3503
rect 25058 3431 25104 3469
rect 25058 3397 25064 3431
rect 25098 3397 25104 3431
rect 25058 3359 25104 3397
rect 25058 3325 25064 3359
rect 25098 3325 25104 3359
rect 25058 3287 25104 3325
rect 25058 3253 25064 3287
rect 25098 3253 25104 3287
rect 25058 3215 25104 3253
rect 25058 3181 25064 3215
rect 25098 3181 25104 3215
rect 25058 3143 25104 3181
rect 25058 3109 25064 3143
rect 25098 3109 25104 3143
rect 25058 3071 25104 3109
rect 25058 3037 25064 3071
rect 25098 3037 25104 3071
rect 25058 2999 25104 3037
rect 25058 2965 25064 2999
rect 25098 2965 25104 2999
rect 25058 2927 25104 2965
rect 25058 2893 25064 2927
rect 25098 2893 25104 2927
rect 25058 2855 25104 2893
rect 25058 2821 25064 2855
rect 25098 2821 25104 2855
rect 25058 2783 25104 2821
rect 25058 2749 25064 2783
rect 25098 2749 25104 2783
rect 25058 2711 25104 2749
rect 25058 2677 25064 2711
rect 25098 2677 25104 2711
rect 25058 2639 25104 2677
rect 25058 2605 25064 2639
rect 25098 2605 25104 2639
rect 25058 2567 25104 2605
rect 25058 2533 25064 2567
rect 25098 2533 25104 2567
rect 25058 2518 25104 2533
rect 25154 3503 25200 3518
rect 25154 3469 25160 3503
rect 25194 3469 25200 3503
rect 25154 3431 25200 3469
rect 25154 3397 25160 3431
rect 25194 3397 25200 3431
rect 25154 3359 25200 3397
rect 25154 3325 25160 3359
rect 25194 3325 25200 3359
rect 25154 3287 25200 3325
rect 25154 3253 25160 3287
rect 25194 3253 25200 3287
rect 25154 3215 25200 3253
rect 25154 3181 25160 3215
rect 25194 3181 25200 3215
rect 25154 3143 25200 3181
rect 25154 3109 25160 3143
rect 25194 3109 25200 3143
rect 25154 3071 25200 3109
rect 25154 3037 25160 3071
rect 25194 3037 25200 3071
rect 25154 2999 25200 3037
rect 25154 2965 25160 2999
rect 25194 2965 25200 2999
rect 25154 2927 25200 2965
rect 25154 2893 25160 2927
rect 25194 2893 25200 2927
rect 25154 2855 25200 2893
rect 25154 2821 25160 2855
rect 25194 2821 25200 2855
rect 25154 2783 25200 2821
rect 25154 2749 25160 2783
rect 25194 2749 25200 2783
rect 25154 2711 25200 2749
rect 25154 2677 25160 2711
rect 25194 2677 25200 2711
rect 25154 2639 25200 2677
rect 25154 2605 25160 2639
rect 25194 2605 25200 2639
rect 25154 2567 25200 2605
rect 25154 2533 25160 2567
rect 25194 2533 25200 2567
rect 25154 2518 25200 2533
rect 25250 3503 25296 3518
rect 25250 3469 25256 3503
rect 25290 3469 25296 3503
rect 25250 3431 25296 3469
rect 25250 3397 25256 3431
rect 25290 3397 25296 3431
rect 25250 3359 25296 3397
rect 25250 3325 25256 3359
rect 25290 3325 25296 3359
rect 25250 3287 25296 3325
rect 25250 3253 25256 3287
rect 25290 3253 25296 3287
rect 25250 3215 25296 3253
rect 25250 3181 25256 3215
rect 25290 3181 25296 3215
rect 25250 3143 25296 3181
rect 25250 3109 25256 3143
rect 25290 3109 25296 3143
rect 25250 3071 25296 3109
rect 25250 3037 25256 3071
rect 25290 3037 25296 3071
rect 25250 2999 25296 3037
rect 25250 2965 25256 2999
rect 25290 2965 25296 2999
rect 25250 2927 25296 2965
rect 25250 2893 25256 2927
rect 25290 2893 25296 2927
rect 25250 2855 25296 2893
rect 25250 2821 25256 2855
rect 25290 2821 25296 2855
rect 25250 2783 25296 2821
rect 25250 2749 25256 2783
rect 25290 2749 25296 2783
rect 25250 2711 25296 2749
rect 25250 2677 25256 2711
rect 25290 2677 25296 2711
rect 25250 2639 25296 2677
rect 25250 2605 25256 2639
rect 25290 2605 25296 2639
rect 25250 2567 25296 2605
rect 25250 2533 25256 2567
rect 25290 2533 25296 2567
rect 25250 2518 25296 2533
rect 25346 3503 25392 3518
rect 25346 3469 25352 3503
rect 25386 3469 25392 3503
rect 25346 3431 25392 3469
rect 25346 3397 25352 3431
rect 25386 3397 25392 3431
rect 25346 3359 25392 3397
rect 25346 3325 25352 3359
rect 25386 3325 25392 3359
rect 25346 3287 25392 3325
rect 25346 3253 25352 3287
rect 25386 3253 25392 3287
rect 25346 3215 25392 3253
rect 25346 3181 25352 3215
rect 25386 3181 25392 3215
rect 25346 3143 25392 3181
rect 25346 3109 25352 3143
rect 25386 3109 25392 3143
rect 25346 3071 25392 3109
rect 25346 3037 25352 3071
rect 25386 3037 25392 3071
rect 25346 2999 25392 3037
rect 25346 2965 25352 2999
rect 25386 2965 25392 2999
rect 25346 2927 25392 2965
rect 25346 2893 25352 2927
rect 25386 2893 25392 2927
rect 25346 2855 25392 2893
rect 25346 2821 25352 2855
rect 25386 2821 25392 2855
rect 25346 2783 25392 2821
rect 25346 2749 25352 2783
rect 25386 2749 25392 2783
rect 25346 2711 25392 2749
rect 25346 2677 25352 2711
rect 25386 2677 25392 2711
rect 25346 2639 25392 2677
rect 25346 2605 25352 2639
rect 25386 2605 25392 2639
rect 25346 2567 25392 2605
rect 25346 2533 25352 2567
rect 25386 2533 25392 2567
rect 25346 2518 25392 2533
rect 25442 3503 25488 3518
rect 25442 3469 25448 3503
rect 25482 3469 25488 3503
rect 25442 3431 25488 3469
rect 25442 3397 25448 3431
rect 25482 3397 25488 3431
rect 25442 3359 25488 3397
rect 25442 3325 25448 3359
rect 25482 3325 25488 3359
rect 25442 3287 25488 3325
rect 25442 3253 25448 3287
rect 25482 3253 25488 3287
rect 25442 3215 25488 3253
rect 25442 3181 25448 3215
rect 25482 3181 25488 3215
rect 25442 3143 25488 3181
rect 25442 3109 25448 3143
rect 25482 3109 25488 3143
rect 25442 3071 25488 3109
rect 25442 3037 25448 3071
rect 25482 3037 25488 3071
rect 25442 2999 25488 3037
rect 25442 2965 25448 2999
rect 25482 2965 25488 2999
rect 25442 2927 25488 2965
rect 25442 2893 25448 2927
rect 25482 2893 25488 2927
rect 25442 2855 25488 2893
rect 25442 2821 25448 2855
rect 25482 2821 25488 2855
rect 25442 2783 25488 2821
rect 25442 2749 25448 2783
rect 25482 2749 25488 2783
rect 25442 2711 25488 2749
rect 25442 2677 25448 2711
rect 25482 2677 25488 2711
rect 25442 2639 25488 2677
rect 25442 2605 25448 2639
rect 25482 2605 25488 2639
rect 25442 2567 25488 2605
rect 25442 2533 25448 2567
rect 25482 2533 25488 2567
rect 25442 2518 25488 2533
rect 25538 3503 25584 3518
rect 25538 3469 25544 3503
rect 25578 3469 25584 3503
rect 25538 3431 25584 3469
rect 25538 3397 25544 3431
rect 25578 3397 25584 3431
rect 25538 3359 25584 3397
rect 25538 3325 25544 3359
rect 25578 3325 25584 3359
rect 25538 3287 25584 3325
rect 25538 3253 25544 3287
rect 25578 3253 25584 3287
rect 25538 3215 25584 3253
rect 25538 3181 25544 3215
rect 25578 3181 25584 3215
rect 25538 3143 25584 3181
rect 25538 3109 25544 3143
rect 25578 3109 25584 3143
rect 25538 3071 25584 3109
rect 25538 3037 25544 3071
rect 25578 3037 25584 3071
rect 25538 2999 25584 3037
rect 25538 2965 25544 2999
rect 25578 2965 25584 2999
rect 25538 2927 25584 2965
rect 25538 2893 25544 2927
rect 25578 2893 25584 2927
rect 25538 2855 25584 2893
rect 25538 2821 25544 2855
rect 25578 2821 25584 2855
rect 25538 2783 25584 2821
rect 25538 2749 25544 2783
rect 25578 2749 25584 2783
rect 25538 2711 25584 2749
rect 25538 2677 25544 2711
rect 25578 2677 25584 2711
rect 25538 2639 25584 2677
rect 25538 2605 25544 2639
rect 25578 2605 25584 2639
rect 25538 2567 25584 2605
rect 25538 2533 25544 2567
rect 25578 2533 25584 2567
rect 25538 2518 25584 2533
rect 25634 3503 25680 3518
rect 25634 3469 25640 3503
rect 25674 3469 25680 3503
rect 25634 3431 25680 3469
rect 25634 3397 25640 3431
rect 25674 3397 25680 3431
rect 25634 3359 25680 3397
rect 25634 3325 25640 3359
rect 25674 3325 25680 3359
rect 25634 3287 25680 3325
rect 25634 3253 25640 3287
rect 25674 3253 25680 3287
rect 25634 3215 25680 3253
rect 25634 3181 25640 3215
rect 25674 3181 25680 3215
rect 25634 3143 25680 3181
rect 25634 3109 25640 3143
rect 25674 3109 25680 3143
rect 25634 3071 25680 3109
rect 25634 3037 25640 3071
rect 25674 3037 25680 3071
rect 25634 2999 25680 3037
rect 25634 2965 25640 2999
rect 25674 2965 25680 2999
rect 25634 2927 25680 2965
rect 25634 2893 25640 2927
rect 25674 2893 25680 2927
rect 25634 2855 25680 2893
rect 25634 2821 25640 2855
rect 25674 2821 25680 2855
rect 25634 2783 25680 2821
rect 25634 2749 25640 2783
rect 25674 2749 25680 2783
rect 25634 2711 25680 2749
rect 25634 2677 25640 2711
rect 25674 2677 25680 2711
rect 25634 2639 25680 2677
rect 25634 2605 25640 2639
rect 25674 2605 25680 2639
rect 25634 2567 25680 2605
rect 25634 2533 25640 2567
rect 25674 2533 25680 2567
rect 25634 2518 25680 2533
rect 25730 3503 25776 3518
rect 25730 3469 25736 3503
rect 25770 3469 25776 3503
rect 25730 3431 25776 3469
rect 25730 3397 25736 3431
rect 25770 3397 25776 3431
rect 25730 3359 25776 3397
rect 25730 3325 25736 3359
rect 25770 3325 25776 3359
rect 25730 3287 25776 3325
rect 25730 3253 25736 3287
rect 25770 3253 25776 3287
rect 25730 3215 25776 3253
rect 25730 3181 25736 3215
rect 25770 3181 25776 3215
rect 25730 3143 25776 3181
rect 25730 3109 25736 3143
rect 25770 3109 25776 3143
rect 25730 3071 25776 3109
rect 25730 3037 25736 3071
rect 25770 3037 25776 3071
rect 25730 2999 25776 3037
rect 25730 2965 25736 2999
rect 25770 2965 25776 2999
rect 25730 2927 25776 2965
rect 25730 2893 25736 2927
rect 25770 2893 25776 2927
rect 25730 2855 25776 2893
rect 25730 2821 25736 2855
rect 25770 2821 25776 2855
rect 25730 2783 25776 2821
rect 25730 2749 25736 2783
rect 25770 2749 25776 2783
rect 25730 2711 25776 2749
rect 25730 2677 25736 2711
rect 25770 2677 25776 2711
rect 25730 2639 25776 2677
rect 25730 2605 25736 2639
rect 25770 2605 25776 2639
rect 25730 2567 25776 2605
rect 25730 2533 25736 2567
rect 25770 2533 25776 2567
rect 25730 2518 25776 2533
rect 25826 3503 25872 3518
rect 25826 3469 25832 3503
rect 25866 3469 25872 3503
rect 25826 3431 25872 3469
rect 25826 3397 25832 3431
rect 25866 3397 25872 3431
rect 25826 3359 25872 3397
rect 25826 3325 25832 3359
rect 25866 3325 25872 3359
rect 25826 3287 25872 3325
rect 25826 3253 25832 3287
rect 25866 3253 25872 3287
rect 25826 3215 25872 3253
rect 25826 3181 25832 3215
rect 25866 3181 25872 3215
rect 25826 3143 25872 3181
rect 25826 3109 25832 3143
rect 25866 3109 25872 3143
rect 25826 3071 25872 3109
rect 25826 3037 25832 3071
rect 25866 3037 25872 3071
rect 25826 2999 25872 3037
rect 25826 2965 25832 2999
rect 25866 2965 25872 2999
rect 25826 2927 25872 2965
rect 25826 2893 25832 2927
rect 25866 2893 25872 2927
rect 25826 2855 25872 2893
rect 25826 2821 25832 2855
rect 25866 2821 25872 2855
rect 25826 2783 25872 2821
rect 25826 2749 25832 2783
rect 25866 2749 25872 2783
rect 25826 2711 25872 2749
rect 25826 2677 25832 2711
rect 25866 2677 25872 2711
rect 25826 2639 25872 2677
rect 25826 2605 25832 2639
rect 25866 2605 25872 2639
rect 25826 2567 25872 2605
rect 25826 2533 25832 2567
rect 25866 2533 25872 2567
rect 25826 2518 25872 2533
rect 25922 3503 25968 3518
rect 25922 3469 25928 3503
rect 25962 3469 25968 3503
rect 25922 3431 25968 3469
rect 25922 3397 25928 3431
rect 25962 3397 25968 3431
rect 25922 3359 25968 3397
rect 25922 3325 25928 3359
rect 25962 3325 25968 3359
rect 25922 3287 25968 3325
rect 25922 3253 25928 3287
rect 25962 3253 25968 3287
rect 25922 3215 25968 3253
rect 25922 3181 25928 3215
rect 25962 3181 25968 3215
rect 25922 3143 25968 3181
rect 25922 3109 25928 3143
rect 25962 3109 25968 3143
rect 25922 3071 25968 3109
rect 25922 3037 25928 3071
rect 25962 3037 25968 3071
rect 25922 2999 25968 3037
rect 25922 2965 25928 2999
rect 25962 2965 25968 2999
rect 25922 2927 25968 2965
rect 25922 2893 25928 2927
rect 25962 2893 25968 2927
rect 25922 2855 25968 2893
rect 25922 2821 25928 2855
rect 25962 2821 25968 2855
rect 25922 2783 25968 2821
rect 25922 2749 25928 2783
rect 25962 2749 25968 2783
rect 25922 2711 25968 2749
rect 25922 2677 25928 2711
rect 25962 2677 25968 2711
rect 25922 2639 25968 2677
rect 25922 2605 25928 2639
rect 25962 2605 25968 2639
rect 25922 2567 25968 2605
rect 25922 2533 25928 2567
rect 25962 2533 25968 2567
rect 25922 2518 25968 2533
rect 26018 3503 26064 3518
rect 26018 3469 26024 3503
rect 26058 3469 26064 3503
rect 26018 3431 26064 3469
rect 26018 3397 26024 3431
rect 26058 3397 26064 3431
rect 26018 3359 26064 3397
rect 26018 3325 26024 3359
rect 26058 3325 26064 3359
rect 26018 3287 26064 3325
rect 26018 3253 26024 3287
rect 26058 3253 26064 3287
rect 26018 3215 26064 3253
rect 26018 3181 26024 3215
rect 26058 3181 26064 3215
rect 26018 3143 26064 3181
rect 26018 3109 26024 3143
rect 26058 3109 26064 3143
rect 26018 3071 26064 3109
rect 26018 3037 26024 3071
rect 26058 3037 26064 3071
rect 26018 2999 26064 3037
rect 26018 2965 26024 2999
rect 26058 2965 26064 2999
rect 26018 2927 26064 2965
rect 26018 2893 26024 2927
rect 26058 2893 26064 2927
rect 26018 2855 26064 2893
rect 26018 2821 26024 2855
rect 26058 2821 26064 2855
rect 26018 2783 26064 2821
rect 26018 2749 26024 2783
rect 26058 2749 26064 2783
rect 26018 2711 26064 2749
rect 26018 2677 26024 2711
rect 26058 2677 26064 2711
rect 26018 2639 26064 2677
rect 26018 2605 26024 2639
rect 26058 2605 26064 2639
rect 26018 2567 26064 2605
rect 26018 2533 26024 2567
rect 26058 2533 26064 2567
rect 26018 2518 26064 2533
rect 26114 3503 26160 3518
rect 26114 3469 26120 3503
rect 26154 3469 26160 3503
rect 26114 3431 26160 3469
rect 26114 3397 26120 3431
rect 26154 3397 26160 3431
rect 26114 3359 26160 3397
rect 26114 3325 26120 3359
rect 26154 3325 26160 3359
rect 26114 3287 26160 3325
rect 26114 3253 26120 3287
rect 26154 3253 26160 3287
rect 26114 3215 26160 3253
rect 26114 3181 26120 3215
rect 26154 3181 26160 3215
rect 26114 3143 26160 3181
rect 26114 3109 26120 3143
rect 26154 3109 26160 3143
rect 26114 3071 26160 3109
rect 26114 3037 26120 3071
rect 26154 3037 26160 3071
rect 26114 2999 26160 3037
rect 26114 2965 26120 2999
rect 26154 2965 26160 2999
rect 26114 2927 26160 2965
rect 26114 2893 26120 2927
rect 26154 2893 26160 2927
rect 26114 2855 26160 2893
rect 26114 2821 26120 2855
rect 26154 2821 26160 2855
rect 26114 2783 26160 2821
rect 26114 2749 26120 2783
rect 26154 2749 26160 2783
rect 26114 2711 26160 2749
rect 26114 2677 26120 2711
rect 26154 2677 26160 2711
rect 26114 2639 26160 2677
rect 26114 2605 26120 2639
rect 26154 2605 26160 2639
rect 26114 2567 26160 2605
rect 26114 2533 26120 2567
rect 26154 2533 26160 2567
rect 26114 2518 26160 2533
rect 26210 3503 26256 3518
rect 26210 3469 26216 3503
rect 26250 3469 26256 3503
rect 26210 3431 26256 3469
rect 26210 3397 26216 3431
rect 26250 3397 26256 3431
rect 26210 3359 26256 3397
rect 26210 3325 26216 3359
rect 26250 3325 26256 3359
rect 26210 3287 26256 3325
rect 26210 3253 26216 3287
rect 26250 3253 26256 3287
rect 26210 3215 26256 3253
rect 26210 3181 26216 3215
rect 26250 3181 26256 3215
rect 26210 3143 26256 3181
rect 26210 3109 26216 3143
rect 26250 3109 26256 3143
rect 26210 3071 26256 3109
rect 26210 3037 26216 3071
rect 26250 3037 26256 3071
rect 26210 2999 26256 3037
rect 26210 2965 26216 2999
rect 26250 2965 26256 2999
rect 26210 2927 26256 2965
rect 26210 2893 26216 2927
rect 26250 2893 26256 2927
rect 26210 2855 26256 2893
rect 26210 2821 26216 2855
rect 26250 2821 26256 2855
rect 26210 2783 26256 2821
rect 26210 2749 26216 2783
rect 26250 2749 26256 2783
rect 26210 2711 26256 2749
rect 26210 2677 26216 2711
rect 26250 2677 26256 2711
rect 26210 2639 26256 2677
rect 26210 2605 26216 2639
rect 26250 2605 26256 2639
rect 26210 2567 26256 2605
rect 26210 2533 26216 2567
rect 26250 2533 26256 2567
rect 26210 2518 26256 2533
rect 26306 3503 26352 3518
rect 26306 3469 26312 3503
rect 26346 3469 26352 3503
rect 26306 3431 26352 3469
rect 26306 3397 26312 3431
rect 26346 3397 26352 3431
rect 26306 3359 26352 3397
rect 26306 3325 26312 3359
rect 26346 3325 26352 3359
rect 26306 3287 26352 3325
rect 26306 3253 26312 3287
rect 26346 3253 26352 3287
rect 26306 3215 26352 3253
rect 26306 3181 26312 3215
rect 26346 3181 26352 3215
rect 26306 3143 26352 3181
rect 26306 3109 26312 3143
rect 26346 3109 26352 3143
rect 26306 3071 26352 3109
rect 26306 3037 26312 3071
rect 26346 3037 26352 3071
rect 26306 2999 26352 3037
rect 26306 2965 26312 2999
rect 26346 2965 26352 2999
rect 26306 2927 26352 2965
rect 26306 2893 26312 2927
rect 26346 2893 26352 2927
rect 26306 2855 26352 2893
rect 26306 2821 26312 2855
rect 26346 2821 26352 2855
rect 26306 2783 26352 2821
rect 26306 2749 26312 2783
rect 26346 2749 26352 2783
rect 26306 2711 26352 2749
rect 26306 2677 26312 2711
rect 26346 2677 26352 2711
rect 26306 2639 26352 2677
rect 26306 2605 26312 2639
rect 26346 2605 26352 2639
rect 26306 2567 26352 2605
rect 26306 2533 26312 2567
rect 26346 2533 26352 2567
rect 26306 2518 26352 2533
rect 26402 3503 26448 3518
rect 26402 3469 26408 3503
rect 26442 3469 26448 3503
rect 26402 3431 26448 3469
rect 26402 3397 26408 3431
rect 26442 3397 26448 3431
rect 26402 3359 26448 3397
rect 26402 3325 26408 3359
rect 26442 3325 26448 3359
rect 26402 3287 26448 3325
rect 26402 3253 26408 3287
rect 26442 3253 26448 3287
rect 26402 3215 26448 3253
rect 26402 3181 26408 3215
rect 26442 3181 26448 3215
rect 26402 3143 26448 3181
rect 26402 3109 26408 3143
rect 26442 3109 26448 3143
rect 26402 3071 26448 3109
rect 26402 3037 26408 3071
rect 26442 3037 26448 3071
rect 26402 2999 26448 3037
rect 26402 2965 26408 2999
rect 26442 2965 26448 2999
rect 26402 2927 26448 2965
rect 26402 2893 26408 2927
rect 26442 2893 26448 2927
rect 26402 2855 26448 2893
rect 26402 2821 26408 2855
rect 26442 2821 26448 2855
rect 26402 2783 26448 2821
rect 26402 2749 26408 2783
rect 26442 2749 26448 2783
rect 26402 2711 26448 2749
rect 26402 2677 26408 2711
rect 26442 2677 26448 2711
rect 26402 2639 26448 2677
rect 26402 2605 26408 2639
rect 26442 2605 26448 2639
rect 26402 2567 26448 2605
rect 26402 2533 26408 2567
rect 26442 2533 26448 2567
rect 26402 2518 26448 2533
rect 26498 3503 26544 3518
rect 26498 3469 26504 3503
rect 26538 3469 26544 3503
rect 26498 3431 26544 3469
rect 26498 3397 26504 3431
rect 26538 3397 26544 3431
rect 26498 3359 26544 3397
rect 26498 3325 26504 3359
rect 26538 3325 26544 3359
rect 26498 3287 26544 3325
rect 26498 3253 26504 3287
rect 26538 3253 26544 3287
rect 26498 3215 26544 3253
rect 26498 3181 26504 3215
rect 26538 3181 26544 3215
rect 26498 3143 26544 3181
rect 26498 3109 26504 3143
rect 26538 3109 26544 3143
rect 26498 3071 26544 3109
rect 26498 3037 26504 3071
rect 26538 3037 26544 3071
rect 26498 2999 26544 3037
rect 26498 2965 26504 2999
rect 26538 2965 26544 2999
rect 26498 2927 26544 2965
rect 26498 2893 26504 2927
rect 26538 2893 26544 2927
rect 26498 2855 26544 2893
rect 26498 2821 26504 2855
rect 26538 2821 26544 2855
rect 26498 2783 26544 2821
rect 26498 2749 26504 2783
rect 26538 2749 26544 2783
rect 26498 2711 26544 2749
rect 26498 2677 26504 2711
rect 26538 2677 26544 2711
rect 26498 2639 26544 2677
rect 26498 2605 26504 2639
rect 26538 2605 26544 2639
rect 26498 2567 26544 2605
rect 26498 2533 26504 2567
rect 26538 2533 26544 2567
rect 26498 2518 26544 2533
rect 26726 3511 26772 3526
rect 26726 3477 26732 3511
rect 26766 3477 26772 3511
rect 26726 3439 26772 3477
rect 26726 3405 26732 3439
rect 26766 3405 26772 3439
rect 26726 3367 26772 3405
rect 26726 3333 26732 3367
rect 26766 3333 26772 3367
rect 26726 3295 26772 3333
rect 26726 3261 26732 3295
rect 26766 3261 26772 3295
rect 26726 3223 26772 3261
rect 26726 3189 26732 3223
rect 26766 3189 26772 3223
rect 26726 3151 26772 3189
rect 26726 3117 26732 3151
rect 26766 3117 26772 3151
rect 26726 3079 26772 3117
rect 26726 3045 26732 3079
rect 26766 3045 26772 3079
rect 26726 3007 26772 3045
rect 26726 2973 26732 3007
rect 26766 2973 26772 3007
rect 26726 2935 26772 2973
rect 26726 2901 26732 2935
rect 26766 2901 26772 2935
rect 26726 2863 26772 2901
rect 26726 2829 26732 2863
rect 26766 2829 26772 2863
rect 26726 2791 26772 2829
rect 26726 2757 26732 2791
rect 26766 2757 26772 2791
rect 26726 2719 26772 2757
rect 26726 2685 26732 2719
rect 26766 2685 26772 2719
rect 26726 2647 26772 2685
rect 26726 2613 26732 2647
rect 26766 2613 26772 2647
rect 26726 2575 26772 2613
rect 26726 2541 26732 2575
rect 26766 2541 26772 2575
rect 26726 2526 26772 2541
rect 26822 3511 26868 3526
rect 26822 3477 26828 3511
rect 26862 3477 26868 3511
rect 26822 3439 26868 3477
rect 26822 3405 26828 3439
rect 26862 3405 26868 3439
rect 26822 3367 26868 3405
rect 26822 3333 26828 3367
rect 26862 3333 26868 3367
rect 26822 3295 26868 3333
rect 26822 3261 26828 3295
rect 26862 3261 26868 3295
rect 26822 3223 26868 3261
rect 26822 3189 26828 3223
rect 26862 3189 26868 3223
rect 26822 3151 26868 3189
rect 26822 3117 26828 3151
rect 26862 3117 26868 3151
rect 26822 3079 26868 3117
rect 26822 3045 26828 3079
rect 26862 3045 26868 3079
rect 26822 3007 26868 3045
rect 26822 2973 26828 3007
rect 26862 2973 26868 3007
rect 26822 2935 26868 2973
rect 26822 2901 26828 2935
rect 26862 2901 26868 2935
rect 26822 2863 26868 2901
rect 26822 2829 26828 2863
rect 26862 2829 26868 2863
rect 26822 2791 26868 2829
rect 26822 2757 26828 2791
rect 26862 2757 26868 2791
rect 26822 2719 26868 2757
rect 26822 2685 26828 2719
rect 26862 2685 26868 2719
rect 26822 2647 26868 2685
rect 26822 2613 26828 2647
rect 26862 2613 26868 2647
rect 26822 2575 26868 2613
rect 26822 2541 26828 2575
rect 26862 2541 26868 2575
rect 26822 2526 26868 2541
rect 26918 3511 26964 3526
rect 26918 3477 26924 3511
rect 26958 3477 26964 3511
rect 26918 3439 26964 3477
rect 26918 3405 26924 3439
rect 26958 3405 26964 3439
rect 26918 3367 26964 3405
rect 26918 3333 26924 3367
rect 26958 3333 26964 3367
rect 26918 3295 26964 3333
rect 26918 3261 26924 3295
rect 26958 3261 26964 3295
rect 26918 3223 26964 3261
rect 26918 3189 26924 3223
rect 26958 3189 26964 3223
rect 26918 3151 26964 3189
rect 26918 3117 26924 3151
rect 26958 3117 26964 3151
rect 26918 3079 26964 3117
rect 26918 3045 26924 3079
rect 26958 3045 26964 3079
rect 26918 3007 26964 3045
rect 26918 2973 26924 3007
rect 26958 2973 26964 3007
rect 26918 2935 26964 2973
rect 26918 2901 26924 2935
rect 26958 2901 26964 2935
rect 26918 2863 26964 2901
rect 26918 2829 26924 2863
rect 26958 2829 26964 2863
rect 26918 2791 26964 2829
rect 26918 2757 26924 2791
rect 26958 2757 26964 2791
rect 26918 2719 26964 2757
rect 26918 2685 26924 2719
rect 26958 2685 26964 2719
rect 26918 2647 26964 2685
rect 26918 2613 26924 2647
rect 26958 2613 26964 2647
rect 26918 2575 26964 2613
rect 26918 2541 26924 2575
rect 26958 2541 26964 2575
rect 26918 2526 26964 2541
rect 27014 3511 27060 3526
rect 27014 3477 27020 3511
rect 27054 3477 27060 3511
rect 27014 3439 27060 3477
rect 27014 3405 27020 3439
rect 27054 3405 27060 3439
rect 27014 3367 27060 3405
rect 27014 3333 27020 3367
rect 27054 3333 27060 3367
rect 27014 3295 27060 3333
rect 27014 3261 27020 3295
rect 27054 3261 27060 3295
rect 27014 3223 27060 3261
rect 27014 3189 27020 3223
rect 27054 3189 27060 3223
rect 27014 3151 27060 3189
rect 27014 3117 27020 3151
rect 27054 3117 27060 3151
rect 27014 3079 27060 3117
rect 27014 3045 27020 3079
rect 27054 3045 27060 3079
rect 27014 3007 27060 3045
rect 27014 2973 27020 3007
rect 27054 2973 27060 3007
rect 27014 2935 27060 2973
rect 27014 2901 27020 2935
rect 27054 2901 27060 2935
rect 27014 2863 27060 2901
rect 27014 2829 27020 2863
rect 27054 2829 27060 2863
rect 27014 2791 27060 2829
rect 27014 2757 27020 2791
rect 27054 2757 27060 2791
rect 27014 2719 27060 2757
rect 27014 2685 27020 2719
rect 27054 2685 27060 2719
rect 27014 2647 27060 2685
rect 27014 2613 27020 2647
rect 27054 2613 27060 2647
rect 27014 2575 27060 2613
rect 27014 2541 27020 2575
rect 27054 2541 27060 2575
rect 27014 2526 27060 2541
rect 27110 3511 27156 3526
rect 27110 3477 27116 3511
rect 27150 3477 27156 3511
rect 27110 3439 27156 3477
rect 27110 3405 27116 3439
rect 27150 3405 27156 3439
rect 27110 3367 27156 3405
rect 27110 3333 27116 3367
rect 27150 3333 27156 3367
rect 27110 3295 27156 3333
rect 27110 3261 27116 3295
rect 27150 3261 27156 3295
rect 27110 3223 27156 3261
rect 27110 3189 27116 3223
rect 27150 3189 27156 3223
rect 27110 3151 27156 3189
rect 27110 3117 27116 3151
rect 27150 3117 27156 3151
rect 27110 3079 27156 3117
rect 27110 3045 27116 3079
rect 27150 3045 27156 3079
rect 27110 3007 27156 3045
rect 27110 2973 27116 3007
rect 27150 2973 27156 3007
rect 27110 2935 27156 2973
rect 27110 2901 27116 2935
rect 27150 2901 27156 2935
rect 27110 2863 27156 2901
rect 27110 2829 27116 2863
rect 27150 2829 27156 2863
rect 27110 2791 27156 2829
rect 27110 2757 27116 2791
rect 27150 2757 27156 2791
rect 27110 2719 27156 2757
rect 27110 2685 27116 2719
rect 27150 2685 27156 2719
rect 27110 2647 27156 2685
rect 27110 2613 27116 2647
rect 27150 2613 27156 2647
rect 27110 2575 27156 2613
rect 27110 2541 27116 2575
rect 27150 2541 27156 2575
rect 27110 2526 27156 2541
rect 27206 3511 27252 3526
rect 27206 3477 27212 3511
rect 27246 3477 27252 3511
rect 27206 3439 27252 3477
rect 27206 3405 27212 3439
rect 27246 3405 27252 3439
rect 27206 3367 27252 3405
rect 27206 3333 27212 3367
rect 27246 3333 27252 3367
rect 27206 3295 27252 3333
rect 27206 3261 27212 3295
rect 27246 3261 27252 3295
rect 27206 3223 27252 3261
rect 27206 3189 27212 3223
rect 27246 3189 27252 3223
rect 27206 3151 27252 3189
rect 27206 3117 27212 3151
rect 27246 3117 27252 3151
rect 27206 3079 27252 3117
rect 27206 3045 27212 3079
rect 27246 3045 27252 3079
rect 27206 3007 27252 3045
rect 27206 2973 27212 3007
rect 27246 2973 27252 3007
rect 27206 2935 27252 2973
rect 27206 2901 27212 2935
rect 27246 2901 27252 2935
rect 27206 2863 27252 2901
rect 27206 2829 27212 2863
rect 27246 2829 27252 2863
rect 27206 2791 27252 2829
rect 27206 2757 27212 2791
rect 27246 2757 27252 2791
rect 27206 2719 27252 2757
rect 27206 2685 27212 2719
rect 27246 2685 27252 2719
rect 27206 2647 27252 2685
rect 27206 2613 27212 2647
rect 27246 2613 27252 2647
rect 27206 2575 27252 2613
rect 27206 2541 27212 2575
rect 27246 2541 27252 2575
rect 27206 2526 27252 2541
rect 27302 3511 27348 3526
rect 27302 3477 27308 3511
rect 27342 3477 27348 3511
rect 27302 3439 27348 3477
rect 27302 3405 27308 3439
rect 27342 3405 27348 3439
rect 27302 3367 27348 3405
rect 27302 3333 27308 3367
rect 27342 3333 27348 3367
rect 27302 3295 27348 3333
rect 27302 3261 27308 3295
rect 27342 3261 27348 3295
rect 27302 3223 27348 3261
rect 27302 3189 27308 3223
rect 27342 3189 27348 3223
rect 27302 3151 27348 3189
rect 27302 3117 27308 3151
rect 27342 3117 27348 3151
rect 27302 3079 27348 3117
rect 27302 3045 27308 3079
rect 27342 3045 27348 3079
rect 27302 3007 27348 3045
rect 27302 2973 27308 3007
rect 27342 2973 27348 3007
rect 27302 2935 27348 2973
rect 27302 2901 27308 2935
rect 27342 2901 27348 2935
rect 27302 2863 27348 2901
rect 27302 2829 27308 2863
rect 27342 2829 27348 2863
rect 27302 2791 27348 2829
rect 27302 2757 27308 2791
rect 27342 2757 27348 2791
rect 27302 2719 27348 2757
rect 27302 2685 27308 2719
rect 27342 2685 27348 2719
rect 27302 2647 27348 2685
rect 27302 2613 27308 2647
rect 27342 2613 27348 2647
rect 27302 2575 27348 2613
rect 27302 2541 27308 2575
rect 27342 2541 27348 2575
rect 27302 2526 27348 2541
rect 27398 3511 27444 3526
rect 27398 3477 27404 3511
rect 27438 3477 27444 3511
rect 27398 3439 27444 3477
rect 27398 3405 27404 3439
rect 27438 3405 27444 3439
rect 27398 3367 27444 3405
rect 27398 3333 27404 3367
rect 27438 3333 27444 3367
rect 27398 3295 27444 3333
rect 27398 3261 27404 3295
rect 27438 3261 27444 3295
rect 27398 3223 27444 3261
rect 27398 3189 27404 3223
rect 27438 3189 27444 3223
rect 27398 3151 27444 3189
rect 27398 3117 27404 3151
rect 27438 3117 27444 3151
rect 27398 3079 27444 3117
rect 27398 3045 27404 3079
rect 27438 3045 27444 3079
rect 27398 3007 27444 3045
rect 27398 2973 27404 3007
rect 27438 2973 27444 3007
rect 27398 2935 27444 2973
rect 27398 2901 27404 2935
rect 27438 2901 27444 2935
rect 27398 2863 27444 2901
rect 27398 2829 27404 2863
rect 27438 2829 27444 2863
rect 27398 2791 27444 2829
rect 27398 2757 27404 2791
rect 27438 2757 27444 2791
rect 27398 2719 27444 2757
rect 27398 2685 27404 2719
rect 27438 2685 27444 2719
rect 27398 2647 27444 2685
rect 27398 2613 27404 2647
rect 27438 2613 27444 2647
rect 27398 2575 27444 2613
rect 27398 2541 27404 2575
rect 27438 2541 27444 2575
rect 27398 2526 27444 2541
rect 27494 3511 27540 3526
rect 27494 3477 27500 3511
rect 27534 3477 27540 3511
rect 27494 3439 27540 3477
rect 27494 3405 27500 3439
rect 27534 3405 27540 3439
rect 27494 3367 27540 3405
rect 27494 3333 27500 3367
rect 27534 3333 27540 3367
rect 27494 3295 27540 3333
rect 27494 3261 27500 3295
rect 27534 3261 27540 3295
rect 27494 3223 27540 3261
rect 27494 3189 27500 3223
rect 27534 3189 27540 3223
rect 27494 3151 27540 3189
rect 27494 3117 27500 3151
rect 27534 3117 27540 3151
rect 27494 3079 27540 3117
rect 27494 3045 27500 3079
rect 27534 3045 27540 3079
rect 27494 3007 27540 3045
rect 27494 2973 27500 3007
rect 27534 2973 27540 3007
rect 27494 2935 27540 2973
rect 27494 2901 27500 2935
rect 27534 2901 27540 2935
rect 27494 2863 27540 2901
rect 27494 2829 27500 2863
rect 27534 2829 27540 2863
rect 27494 2791 27540 2829
rect 27494 2757 27500 2791
rect 27534 2757 27540 2791
rect 27494 2719 27540 2757
rect 27494 2685 27500 2719
rect 27534 2685 27540 2719
rect 27494 2647 27540 2685
rect 27494 2613 27500 2647
rect 27534 2613 27540 2647
rect 27494 2575 27540 2613
rect 27494 2541 27500 2575
rect 27534 2541 27540 2575
rect 27494 2526 27540 2541
rect 27590 3511 27636 3526
rect 27590 3477 27596 3511
rect 27630 3477 27636 3511
rect 27590 3439 27636 3477
rect 27590 3405 27596 3439
rect 27630 3405 27636 3439
rect 27590 3367 27636 3405
rect 27590 3333 27596 3367
rect 27630 3333 27636 3367
rect 27590 3295 27636 3333
rect 27590 3261 27596 3295
rect 27630 3261 27636 3295
rect 27590 3223 27636 3261
rect 27590 3189 27596 3223
rect 27630 3189 27636 3223
rect 27590 3151 27636 3189
rect 27590 3117 27596 3151
rect 27630 3117 27636 3151
rect 27590 3079 27636 3117
rect 27590 3045 27596 3079
rect 27630 3045 27636 3079
rect 27590 3007 27636 3045
rect 27590 2973 27596 3007
rect 27630 2973 27636 3007
rect 27590 2935 27636 2973
rect 27590 2901 27596 2935
rect 27630 2901 27636 2935
rect 27590 2863 27636 2901
rect 27590 2829 27596 2863
rect 27630 2829 27636 2863
rect 27590 2791 27636 2829
rect 27590 2757 27596 2791
rect 27630 2757 27636 2791
rect 27590 2719 27636 2757
rect 27590 2685 27596 2719
rect 27630 2685 27636 2719
rect 27590 2647 27636 2685
rect 27590 2613 27596 2647
rect 27630 2613 27636 2647
rect 27590 2575 27636 2613
rect 27590 2541 27596 2575
rect 27630 2541 27636 2575
rect 27590 2526 27636 2541
rect 27686 3511 27732 3526
rect 27686 3477 27692 3511
rect 27726 3477 27732 3511
rect 27686 3439 27732 3477
rect 27686 3405 27692 3439
rect 27726 3405 27732 3439
rect 27686 3367 27732 3405
rect 27686 3333 27692 3367
rect 27726 3333 27732 3367
rect 27686 3295 27732 3333
rect 27686 3261 27692 3295
rect 27726 3261 27732 3295
rect 27686 3223 27732 3261
rect 27686 3189 27692 3223
rect 27726 3189 27732 3223
rect 27686 3151 27732 3189
rect 27686 3117 27692 3151
rect 27726 3117 27732 3151
rect 27686 3079 27732 3117
rect 27686 3045 27692 3079
rect 27726 3045 27732 3079
rect 27686 3007 27732 3045
rect 27686 2973 27692 3007
rect 27726 2973 27732 3007
rect 27686 2935 27732 2973
rect 27686 2901 27692 2935
rect 27726 2901 27732 2935
rect 27686 2863 27732 2901
rect 27686 2829 27692 2863
rect 27726 2829 27732 2863
rect 27686 2791 27732 2829
rect 27686 2757 27692 2791
rect 27726 2757 27732 2791
rect 27686 2719 27732 2757
rect 27686 2685 27692 2719
rect 27726 2685 27732 2719
rect 27686 2647 27732 2685
rect 27686 2613 27692 2647
rect 27726 2613 27732 2647
rect 27686 2575 27732 2613
rect 27686 2541 27692 2575
rect 27726 2541 27732 2575
rect 27686 2526 27732 2541
rect 27782 3511 27828 3526
rect 27782 3477 27788 3511
rect 27822 3477 27828 3511
rect 27782 3439 27828 3477
rect 27782 3405 27788 3439
rect 27822 3405 27828 3439
rect 27782 3367 27828 3405
rect 27782 3333 27788 3367
rect 27822 3333 27828 3367
rect 27782 3295 27828 3333
rect 27782 3261 27788 3295
rect 27822 3261 27828 3295
rect 27782 3223 27828 3261
rect 27782 3189 27788 3223
rect 27822 3189 27828 3223
rect 27782 3151 27828 3189
rect 27782 3117 27788 3151
rect 27822 3117 27828 3151
rect 27782 3079 27828 3117
rect 27782 3045 27788 3079
rect 27822 3045 27828 3079
rect 27782 3007 27828 3045
rect 27782 2973 27788 3007
rect 27822 2973 27828 3007
rect 27782 2935 27828 2973
rect 27782 2901 27788 2935
rect 27822 2901 27828 2935
rect 27782 2863 27828 2901
rect 27782 2829 27788 2863
rect 27822 2829 27828 2863
rect 27782 2791 27828 2829
rect 27782 2757 27788 2791
rect 27822 2757 27828 2791
rect 27782 2719 27828 2757
rect 27782 2685 27788 2719
rect 27822 2685 27828 2719
rect 27782 2647 27828 2685
rect 27782 2613 27788 2647
rect 27822 2613 27828 2647
rect 27782 2575 27828 2613
rect 27782 2541 27788 2575
rect 27822 2541 27828 2575
rect 27782 2526 27828 2541
rect 27878 3511 27924 3526
rect 27878 3477 27884 3511
rect 27918 3477 27924 3511
rect 27878 3439 27924 3477
rect 27878 3405 27884 3439
rect 27918 3405 27924 3439
rect 27878 3367 27924 3405
rect 27878 3333 27884 3367
rect 27918 3333 27924 3367
rect 27878 3295 27924 3333
rect 27878 3261 27884 3295
rect 27918 3261 27924 3295
rect 27878 3223 27924 3261
rect 27878 3189 27884 3223
rect 27918 3189 27924 3223
rect 27878 3151 27924 3189
rect 27878 3117 27884 3151
rect 27918 3117 27924 3151
rect 27878 3079 27924 3117
rect 27878 3045 27884 3079
rect 27918 3045 27924 3079
rect 27878 3007 27924 3045
rect 27878 2973 27884 3007
rect 27918 2973 27924 3007
rect 27878 2935 27924 2973
rect 27878 2901 27884 2935
rect 27918 2901 27924 2935
rect 27878 2863 27924 2901
rect 27878 2829 27884 2863
rect 27918 2829 27924 2863
rect 27878 2791 27924 2829
rect 27878 2757 27884 2791
rect 27918 2757 27924 2791
rect 27878 2719 27924 2757
rect 27878 2685 27884 2719
rect 27918 2685 27924 2719
rect 27878 2647 27924 2685
rect 27878 2613 27884 2647
rect 27918 2613 27924 2647
rect 27878 2575 27924 2613
rect 27878 2541 27884 2575
rect 27918 2541 27924 2575
rect 27878 2526 27924 2541
rect 27974 3511 28020 3526
rect 27974 3477 27980 3511
rect 28014 3477 28020 3511
rect 27974 3439 28020 3477
rect 27974 3405 27980 3439
rect 28014 3405 28020 3439
rect 27974 3367 28020 3405
rect 27974 3333 27980 3367
rect 28014 3333 28020 3367
rect 27974 3295 28020 3333
rect 27974 3261 27980 3295
rect 28014 3261 28020 3295
rect 27974 3223 28020 3261
rect 27974 3189 27980 3223
rect 28014 3189 28020 3223
rect 27974 3151 28020 3189
rect 27974 3117 27980 3151
rect 28014 3117 28020 3151
rect 27974 3079 28020 3117
rect 27974 3045 27980 3079
rect 28014 3045 28020 3079
rect 27974 3007 28020 3045
rect 27974 2973 27980 3007
rect 28014 2973 28020 3007
rect 27974 2935 28020 2973
rect 27974 2901 27980 2935
rect 28014 2901 28020 2935
rect 27974 2863 28020 2901
rect 27974 2829 27980 2863
rect 28014 2829 28020 2863
rect 27974 2791 28020 2829
rect 27974 2757 27980 2791
rect 28014 2757 28020 2791
rect 27974 2719 28020 2757
rect 27974 2685 27980 2719
rect 28014 2685 28020 2719
rect 27974 2647 28020 2685
rect 27974 2613 27980 2647
rect 28014 2613 28020 2647
rect 27974 2575 28020 2613
rect 27974 2541 27980 2575
rect 28014 2541 28020 2575
rect 27974 2526 28020 2541
rect 28070 3511 28116 3526
rect 28070 3477 28076 3511
rect 28110 3477 28116 3511
rect 28070 3439 28116 3477
rect 28070 3405 28076 3439
rect 28110 3405 28116 3439
rect 28070 3367 28116 3405
rect 28070 3333 28076 3367
rect 28110 3333 28116 3367
rect 28070 3295 28116 3333
rect 28070 3261 28076 3295
rect 28110 3261 28116 3295
rect 28070 3223 28116 3261
rect 28070 3189 28076 3223
rect 28110 3189 28116 3223
rect 28070 3151 28116 3189
rect 28070 3117 28076 3151
rect 28110 3117 28116 3151
rect 28070 3079 28116 3117
rect 28070 3045 28076 3079
rect 28110 3045 28116 3079
rect 28070 3007 28116 3045
rect 28070 2973 28076 3007
rect 28110 2973 28116 3007
rect 28070 2935 28116 2973
rect 28070 2901 28076 2935
rect 28110 2901 28116 2935
rect 28070 2863 28116 2901
rect 28070 2829 28076 2863
rect 28110 2829 28116 2863
rect 28070 2791 28116 2829
rect 28070 2757 28076 2791
rect 28110 2757 28116 2791
rect 28070 2719 28116 2757
rect 28070 2685 28076 2719
rect 28110 2685 28116 2719
rect 28070 2647 28116 2685
rect 28070 2613 28076 2647
rect 28110 2613 28116 2647
rect 28070 2575 28116 2613
rect 28070 2541 28076 2575
rect 28110 2541 28116 2575
rect 28070 2526 28116 2541
rect 28166 3511 28212 3526
rect 28166 3477 28172 3511
rect 28206 3477 28212 3511
rect 28166 3439 28212 3477
rect 28166 3405 28172 3439
rect 28206 3405 28212 3439
rect 28166 3367 28212 3405
rect 28166 3333 28172 3367
rect 28206 3333 28212 3367
rect 28166 3295 28212 3333
rect 28166 3261 28172 3295
rect 28206 3261 28212 3295
rect 28166 3223 28212 3261
rect 28166 3189 28172 3223
rect 28206 3189 28212 3223
rect 28166 3151 28212 3189
rect 28166 3117 28172 3151
rect 28206 3117 28212 3151
rect 28166 3079 28212 3117
rect 28166 3045 28172 3079
rect 28206 3045 28212 3079
rect 28166 3007 28212 3045
rect 28166 2973 28172 3007
rect 28206 2973 28212 3007
rect 28166 2935 28212 2973
rect 28166 2901 28172 2935
rect 28206 2901 28212 2935
rect 28166 2863 28212 2901
rect 28166 2829 28172 2863
rect 28206 2829 28212 2863
rect 28166 2791 28212 2829
rect 28166 2757 28172 2791
rect 28206 2757 28212 2791
rect 28166 2719 28212 2757
rect 28166 2685 28172 2719
rect 28206 2685 28212 2719
rect 28166 2647 28212 2685
rect 28166 2613 28172 2647
rect 28206 2613 28212 2647
rect 28166 2575 28212 2613
rect 28166 2541 28172 2575
rect 28206 2541 28212 2575
rect 28166 2526 28212 2541
rect 28262 3511 28308 3526
rect 28262 3477 28268 3511
rect 28302 3477 28308 3511
rect 28262 3439 28308 3477
rect 28262 3405 28268 3439
rect 28302 3405 28308 3439
rect 28262 3367 28308 3405
rect 28262 3333 28268 3367
rect 28302 3333 28308 3367
rect 28262 3295 28308 3333
rect 28262 3261 28268 3295
rect 28302 3261 28308 3295
rect 28262 3223 28308 3261
rect 28262 3189 28268 3223
rect 28302 3189 28308 3223
rect 28262 3151 28308 3189
rect 28262 3117 28268 3151
rect 28302 3117 28308 3151
rect 28262 3079 28308 3117
rect 28262 3045 28268 3079
rect 28302 3045 28308 3079
rect 28262 3007 28308 3045
rect 28262 2973 28268 3007
rect 28302 2973 28308 3007
rect 28262 2935 28308 2973
rect 28262 2901 28268 2935
rect 28302 2901 28308 2935
rect 28262 2863 28308 2901
rect 28262 2829 28268 2863
rect 28302 2829 28308 2863
rect 28262 2791 28308 2829
rect 28262 2757 28268 2791
rect 28302 2757 28308 2791
rect 28262 2719 28308 2757
rect 28262 2685 28268 2719
rect 28302 2685 28308 2719
rect 28262 2647 28308 2685
rect 28262 2613 28268 2647
rect 28302 2613 28308 2647
rect 28262 2575 28308 2613
rect 28262 2541 28268 2575
rect 28302 2541 28308 2575
rect 28262 2526 28308 2541
rect 28358 3511 28404 3526
rect 28358 3477 28364 3511
rect 28398 3477 28404 3511
rect 28358 3439 28404 3477
rect 28358 3405 28364 3439
rect 28398 3405 28404 3439
rect 28358 3367 28404 3405
rect 28358 3333 28364 3367
rect 28398 3333 28404 3367
rect 28358 3295 28404 3333
rect 28358 3261 28364 3295
rect 28398 3261 28404 3295
rect 28358 3223 28404 3261
rect 28358 3189 28364 3223
rect 28398 3189 28404 3223
rect 28358 3151 28404 3189
rect 28358 3117 28364 3151
rect 28398 3117 28404 3151
rect 28358 3079 28404 3117
rect 28358 3045 28364 3079
rect 28398 3045 28404 3079
rect 28358 3007 28404 3045
rect 28358 2973 28364 3007
rect 28398 2973 28404 3007
rect 28358 2935 28404 2973
rect 28358 2901 28364 2935
rect 28398 2901 28404 2935
rect 28358 2863 28404 2901
rect 28358 2829 28364 2863
rect 28398 2829 28404 2863
rect 28358 2791 28404 2829
rect 28358 2757 28364 2791
rect 28398 2757 28404 2791
rect 28358 2719 28404 2757
rect 28358 2685 28364 2719
rect 28398 2685 28404 2719
rect 28358 2647 28404 2685
rect 28358 2613 28364 2647
rect 28398 2613 28404 2647
rect 28358 2575 28404 2613
rect 28358 2541 28364 2575
rect 28398 2541 28404 2575
rect 28358 2526 28404 2541
rect 28454 3511 28500 3526
rect 28454 3477 28460 3511
rect 28494 3477 28500 3511
rect 28454 3439 28500 3477
rect 28454 3405 28460 3439
rect 28494 3405 28500 3439
rect 28454 3367 28500 3405
rect 28454 3333 28460 3367
rect 28494 3333 28500 3367
rect 28454 3295 28500 3333
rect 28454 3261 28460 3295
rect 28494 3261 28500 3295
rect 28454 3223 28500 3261
rect 28454 3189 28460 3223
rect 28494 3189 28500 3223
rect 28454 3151 28500 3189
rect 28454 3117 28460 3151
rect 28494 3117 28500 3151
rect 28454 3079 28500 3117
rect 28454 3045 28460 3079
rect 28494 3045 28500 3079
rect 28454 3007 28500 3045
rect 28454 2973 28460 3007
rect 28494 2973 28500 3007
rect 28454 2935 28500 2973
rect 28454 2901 28460 2935
rect 28494 2901 28500 2935
rect 28454 2863 28500 2901
rect 28454 2829 28460 2863
rect 28494 2829 28500 2863
rect 28454 2791 28500 2829
rect 28454 2757 28460 2791
rect 28494 2757 28500 2791
rect 28454 2719 28500 2757
rect 28454 2685 28460 2719
rect 28494 2685 28500 2719
rect 28454 2647 28500 2685
rect 28454 2613 28460 2647
rect 28494 2613 28500 2647
rect 28454 2575 28500 2613
rect 28454 2541 28460 2575
rect 28494 2541 28500 2575
rect 28454 2526 28500 2541
rect 28550 3511 28596 3526
rect 28550 3477 28556 3511
rect 28590 3477 28596 3511
rect 28550 3439 28596 3477
rect 28550 3405 28556 3439
rect 28590 3405 28596 3439
rect 28550 3367 28596 3405
rect 28550 3333 28556 3367
rect 28590 3333 28596 3367
rect 28550 3295 28596 3333
rect 28550 3261 28556 3295
rect 28590 3261 28596 3295
rect 28550 3223 28596 3261
rect 28550 3189 28556 3223
rect 28590 3189 28596 3223
rect 28550 3151 28596 3189
rect 28550 3117 28556 3151
rect 28590 3117 28596 3151
rect 28550 3079 28596 3117
rect 28550 3045 28556 3079
rect 28590 3045 28596 3079
rect 28550 3007 28596 3045
rect 28550 2973 28556 3007
rect 28590 2973 28596 3007
rect 28550 2935 28596 2973
rect 28550 2901 28556 2935
rect 28590 2901 28596 2935
rect 28550 2863 28596 2901
rect 28550 2829 28556 2863
rect 28590 2829 28596 2863
rect 28550 2791 28596 2829
rect 28550 2757 28556 2791
rect 28590 2757 28596 2791
rect 28550 2719 28596 2757
rect 28550 2685 28556 2719
rect 28590 2685 28596 2719
rect 28550 2647 28596 2685
rect 28550 2613 28556 2647
rect 28590 2613 28596 2647
rect 28550 2575 28596 2613
rect 28550 2541 28556 2575
rect 28590 2541 28596 2575
rect 28550 2526 28596 2541
rect 28646 3511 28692 3526
rect 28646 3477 28652 3511
rect 28686 3477 28692 3511
rect 28646 3439 28692 3477
rect 28646 3405 28652 3439
rect 28686 3405 28692 3439
rect 28646 3367 28692 3405
rect 28646 3333 28652 3367
rect 28686 3333 28692 3367
rect 28646 3295 28692 3333
rect 28646 3261 28652 3295
rect 28686 3261 28692 3295
rect 28646 3223 28692 3261
rect 28646 3189 28652 3223
rect 28686 3189 28692 3223
rect 28646 3151 28692 3189
rect 28646 3117 28652 3151
rect 28686 3117 28692 3151
rect 28646 3079 28692 3117
rect 28646 3045 28652 3079
rect 28686 3045 28692 3079
rect 28646 3007 28692 3045
rect 28646 2973 28652 3007
rect 28686 2973 28692 3007
rect 28646 2935 28692 2973
rect 28646 2901 28652 2935
rect 28686 2901 28692 2935
rect 28646 2863 28692 2901
rect 28646 2829 28652 2863
rect 28686 2829 28692 2863
rect 28646 2791 28692 2829
rect 28646 2757 28652 2791
rect 28686 2757 28692 2791
rect 28646 2719 28692 2757
rect 28646 2685 28652 2719
rect 28686 2685 28692 2719
rect 28646 2647 28692 2685
rect 28646 2613 28652 2647
rect 28686 2613 28692 2647
rect 28646 2575 28692 2613
rect 28646 2541 28652 2575
rect 28686 2541 28692 2575
rect 28646 2526 28692 2541
rect 23244 2336 23546 2338
rect 23244 2156 23273 2336
rect 23517 2156 23546 2336
rect 23244 2154 23546 2156
rect 25244 2337 25542 2340
rect 25244 2157 25271 2337
rect 25515 2157 25542 2337
rect 25244 2154 25542 2157
rect 29162 -5146 29438 3750
<< via1 >>
rect -374 9022 -130 9061
rect -374 8844 -344 9022
rect -344 8844 -166 9022
rect -166 8844 -130 9022
rect -374 8817 -130 8844
rect 1626 9022 1870 9061
rect 1626 8844 1656 9022
rect 1656 8844 1834 9022
rect 1834 8844 1870 9022
rect 1626 8817 1870 8844
rect 3626 9022 3870 9061
rect 3626 8844 3656 9022
rect 3656 8844 3834 9022
rect 3834 8844 3870 9022
rect 3626 8817 3870 8844
rect 5626 9022 5870 9061
rect 5626 8844 5656 9022
rect 5656 8844 5834 9022
rect 5834 8844 5870 9022
rect 5626 8817 5870 8844
rect 7626 9022 7870 9061
rect 7626 8844 7656 9022
rect 7656 8844 7834 9022
rect 7834 8844 7870 9022
rect 7626 8817 7870 8844
rect 9626 9022 9870 9061
rect 9626 8844 9656 9022
rect 9656 8844 9834 9022
rect 9834 8844 9870 9022
rect 9626 8817 9870 8844
rect 11626 9022 11870 9061
rect 11626 8844 11656 9022
rect 11656 8844 11834 9022
rect 11834 8844 11870 9022
rect 11626 8817 11870 8844
rect 13626 9022 13870 9061
rect 13626 8844 13656 9022
rect 13656 8844 13834 9022
rect 13834 8844 13870 9022
rect 13626 8817 13870 8844
rect 15421 9057 15665 9066
rect 15421 8886 15454 9057
rect 15454 8886 15632 9057
rect 15632 8886 15665 9057
rect -1343 8099 -779 8166
rect -1343 7921 -1251 8099
rect -1251 7921 -857 8099
rect -857 7921 -779 8099
rect -1343 7858 -779 7921
rect 15427 8106 15799 8159
rect 15427 7928 15491 8106
rect 15491 7928 15741 8106
rect 15741 7928 15799 8106
rect 15427 7851 15799 7928
rect -23006 4779 -22698 4812
rect -23006 4673 -22950 4779
rect -22950 4673 -22772 4779
rect -22772 4673 -22698 4779
rect -23006 4632 -22698 4673
rect -21002 4771 -20694 4813
rect -21002 4665 -20936 4771
rect -20936 4665 -20758 4771
rect -20758 4665 -20694 4771
rect -21002 4633 -20694 4665
rect -19004 4772 -18696 4811
rect -19004 4666 -18939 4772
rect -18939 4666 -18761 4772
rect -18761 4666 -18696 4772
rect -19004 4631 -18696 4666
rect -16386 4789 -16078 4824
rect -16386 4683 -16317 4789
rect -16317 4683 -16139 4789
rect -16139 4683 -16078 4789
rect -16386 4644 -16078 4683
rect -14382 4778 -14074 4825
rect -14382 4672 -14320 4778
rect -14320 4672 -14142 4778
rect -14142 4672 -14074 4778
rect -14382 4645 -14074 4672
rect -12384 4782 -12076 4827
rect -12384 4676 -12320 4782
rect -12320 4676 -12142 4782
rect -12142 4676 -12076 4782
rect -12384 4647 -12076 4676
rect -10036 4785 -9728 4822
rect -10036 4679 -9969 4785
rect -9969 4679 -9791 4785
rect -9791 4679 -9728 4785
rect -10036 4642 -9728 4679
rect -8037 4777 -7729 4820
rect -8037 4671 -7976 4777
rect -7976 4671 -7798 4777
rect -7798 4671 -7729 4777
rect -8037 4640 -7729 4671
rect -6036 4778 -5728 4820
rect -6036 4672 -5972 4778
rect -5972 4672 -5794 4778
rect -5794 4672 -5728 4778
rect -6036 4640 -5728 4672
rect 2893 6757 2945 6809
rect 5923 6751 5975 6803
rect 8905 6747 8957 6799
rect 12055 6749 12107 6801
rect 14855 6717 14907 6769
rect -17870 3088 -17818 3140
rect -17806 3088 -17754 3140
rect -23091 1628 -22783 1665
rect -23091 1522 -23029 1628
rect -23029 1522 -22851 1628
rect -22851 1522 -22783 1628
rect -23091 1485 -22783 1522
rect -21091 1622 -20783 1664
rect -21091 1516 -21034 1622
rect -21034 1516 -20856 1622
rect -20856 1516 -20783 1622
rect -21091 1484 -20783 1516
rect -19091 1631 -18783 1666
rect -19091 1525 -19026 1631
rect -19026 1525 -18848 1631
rect -18848 1525 -18783 1631
rect -19091 1486 -18783 1525
rect -11002 3106 -10950 3158
rect -16609 1639 -16301 1677
rect -16609 1533 -16546 1639
rect -16546 1533 -16368 1639
rect -16368 1533 -16301 1639
rect -16609 1497 -16301 1533
rect -14409 1636 -14101 1678
rect -14409 1530 -14350 1636
rect -14350 1530 -14172 1636
rect -14172 1530 -14101 1636
rect -14409 1498 -14101 1530
rect -12007 1641 -11699 1677
rect -12007 1535 -11944 1641
rect -11944 1535 -11766 1641
rect -11766 1535 -11699 1641
rect -12007 1497 -11699 1535
rect -4538 3099 -4486 3151
rect -2396 2506 -2244 2668
rect 16985 5450 17229 5487
rect 16985 5344 17019 5450
rect 17019 5344 17197 5450
rect 17197 5344 17229 5450
rect 16985 5307 17229 5344
rect 18984 5442 19228 5484
rect 18984 5336 19014 5442
rect 19014 5336 19192 5442
rect 19192 5336 19228 5442
rect 18984 5304 19228 5336
rect 20985 5444 21229 5484
rect 20985 5338 21017 5444
rect 21017 5338 21195 5444
rect 21195 5338 21229 5444
rect 20985 5304 21229 5338
rect 23530 5447 23774 5483
rect 23530 5341 23566 5447
rect 23566 5341 23744 5447
rect 23744 5341 23774 5447
rect 23530 5303 23774 5341
rect 25531 5446 25775 5484
rect 25531 5340 25603 5446
rect 25603 5340 25709 5446
rect 25709 5340 25775 5446
rect 25531 5304 25775 5340
rect 27531 5441 27775 5483
rect 27531 5335 27563 5441
rect 27563 5335 27741 5441
rect 27741 5335 27775 5441
rect 27531 5303 27775 5335
rect 2101 3735 2153 3787
rect 4933 3717 4985 3769
rect 4602 3568 4696 3662
rect 1642 3358 1744 3472
rect 3663 3253 3715 3305
rect 1409 2961 1461 3013
rect -9408 1637 -9100 1675
rect -9408 1531 -9379 1637
rect -9379 1531 -9129 1637
rect -9129 1531 -9100 1637
rect -9408 1495 -9100 1531
rect -7408 1636 -7100 1675
rect -7408 1530 -7345 1636
rect -7345 1530 -7167 1636
rect -7167 1530 -7100 1636
rect -7408 1495 -7100 1530
rect -5409 1638 -5101 1675
rect -5409 1532 -5345 1638
rect -5345 1532 -5167 1638
rect -5167 1532 -5101 1638
rect -5409 1495 -5101 1532
rect 10023 3715 10075 3767
rect 7127 3427 7179 3479
rect 5605 3163 5657 3215
rect 7304 3099 7356 3151
rect 2570 2540 2622 2592
rect 11081 3717 11133 3769
rect 8691 3608 8743 3660
rect 10409 3419 10461 3471
rect 8772 3354 8824 3406
rect 13081 3419 13133 3471
rect 13441 3412 13493 3464
rect 13901 3429 13953 3481
rect 5570 2540 5622 2592
rect 8571 2545 8623 2597
rect 13578 2915 13630 2967
rect 11570 2516 11622 2568
rect 16487 3768 16539 3820
rect 15324 1856 15408 1948
rect 15471 1618 15523 1670
rect 2779 -67 2831 -15
rect 5735 -63 5787 -11
rect 8765 -77 8817 -25
rect 11853 -77 11905 -25
rect 17919 2299 18163 2339
rect 17919 2193 17947 2299
rect 17947 2193 18125 2299
rect 18125 2193 18163 2299
rect 17919 2159 18163 2193
rect 19919 2299 20163 2339
rect 19919 2193 19954 2299
rect 19954 2193 20132 2299
rect 20132 2193 20163 2299
rect 19919 2159 20163 2193
rect 21918 2302 22162 2339
rect 21918 2196 21949 2302
rect 21949 2196 22127 2302
rect 22127 2196 22162 2302
rect 21918 2159 22162 2196
rect 2889 -514 2941 -462
rect 5639 -512 5691 -460
rect 8677 -512 8729 -460
rect 11751 -498 11803 -446
rect 258 -1038 694 -962
rect 258 -1216 346 -1038
rect 346 -1216 596 -1038
rect 596 -1216 694 -1038
rect 258 -1270 694 -1216
rect 15432 -1019 15740 -960
rect 15432 -1197 15498 -1019
rect 15498 -1197 15676 -1019
rect 15676 -1197 15740 -1019
rect 15432 -1268 15740 -1197
rect 2235 -1643 2269 -1468
rect 2269 -1643 2447 -1468
rect 2447 -1643 2479 -1468
rect 2235 -1648 2479 -1643
rect 4235 -1643 4269 -1468
rect 4269 -1643 4447 -1468
rect 4447 -1643 4479 -1468
rect 4235 -1648 4479 -1643
rect 6235 -1643 6269 -1468
rect 6269 -1643 6447 -1468
rect 6447 -1643 6479 -1468
rect 6235 -1648 6479 -1643
rect 8462 -1660 8493 -1493
rect 8493 -1660 8671 -1493
rect 8671 -1660 8706 -1493
rect 8462 -1673 8706 -1660
rect 10235 -1643 10269 -1468
rect 10269 -1643 10447 -1468
rect 10447 -1643 10479 -1468
rect 10235 -1648 10479 -1643
rect 12235 -1643 12269 -1468
rect 12269 -1643 12447 -1468
rect 12447 -1643 12479 -1468
rect 12235 -1648 12479 -1643
rect 14235 -1643 14269 -1468
rect 14269 -1643 14447 -1468
rect 14447 -1643 14479 -1468
rect 14235 -1648 14479 -1643
rect 22981 3766 23033 3818
rect 23273 2297 23517 2336
rect 23273 2191 23302 2297
rect 23302 2191 23480 2297
rect 23480 2191 23517 2297
rect 23273 2156 23517 2191
rect 25271 2296 25515 2337
rect 25271 2190 25305 2296
rect 25305 2190 25483 2296
rect 25483 2190 25515 2296
rect 25271 2157 25515 2190
<< metal2 >>
rect 15414 9084 15672 9100
rect -382 9061 -122 9084
rect -382 8817 -374 9061
rect -130 8817 -122 9061
rect -382 8794 -122 8817
rect 1618 9061 1878 9084
rect 1618 8817 1626 9061
rect 1870 8817 1878 9061
rect 1618 8794 1878 8817
rect 3618 9061 3878 9084
rect 3618 8817 3626 9061
rect 3870 8817 3878 9061
rect 3618 8794 3878 8817
rect 5618 9061 5878 9084
rect 5618 8817 5626 9061
rect 5870 8817 5878 9061
rect 5618 8794 5878 8817
rect 7618 9061 7878 9084
rect 7618 8817 7626 9061
rect 7870 8817 7878 9061
rect 7618 8794 7878 8817
rect 9618 9061 9878 9084
rect 9618 8817 9626 9061
rect 9870 8817 9878 9061
rect 9618 8794 9878 8817
rect 11618 9061 11878 9084
rect 11618 8817 11626 9061
rect 11870 8817 11878 9061
rect 11618 8794 11878 8817
rect 13618 9061 13878 9084
rect 13618 8817 13626 9061
rect 13870 8817 13878 9061
rect 15414 9066 15435 9084
rect 15651 9066 15672 9084
rect 15414 8886 15421 9066
rect 15665 8886 15672 9066
rect 15414 8868 15435 8886
rect 15651 8868 15672 8886
rect 15414 8852 15672 8868
rect 13618 8794 13878 8817
rect -1350 8166 -772 8192
rect -1350 7858 -1343 8166
rect -779 7858 -772 8166
rect -1350 7832 -772 7858
rect 15404 8159 15822 8188
rect 15404 8153 15427 8159
rect 15799 8153 15822 8159
rect 15404 7857 15425 8153
rect 15801 7857 15822 8153
rect 15404 7851 15427 7857
rect 15799 7851 15822 7857
rect 15404 7822 15822 7851
rect 2814 7344 15236 7564
rect 2888 6809 2950 7344
rect 2888 6757 2893 6809
rect 2945 6757 2950 6809
rect 2888 6742 2950 6757
rect 5918 6803 5980 7344
rect 5918 6751 5923 6803
rect 5975 6751 5980 6803
rect 5918 6738 5980 6751
rect 8900 6799 8962 7344
rect 8900 6747 8905 6799
rect 8957 6747 8962 6799
rect 8900 6732 8962 6747
rect 12050 6801 12112 7344
rect 12050 6749 12055 6801
rect 12107 6749 12112 6801
rect 12050 6734 12112 6749
rect 14850 6769 14912 7344
rect 14850 6717 14855 6769
rect 14907 6717 14912 6769
rect 14850 6702 14912 6717
rect -23006 4812 -22698 4822
rect -23006 4622 -22698 4632
rect -21010 4813 -20686 4836
rect -21010 4633 -21002 4813
rect -20694 4633 -20686 4813
rect -21010 4610 -20686 4633
rect -19010 4811 -18690 4836
rect -19010 4631 -19004 4811
rect -18696 4631 -18690 4811
rect -19010 4606 -18690 4631
rect -16390 4824 -16074 4844
rect -16390 4644 -16386 4824
rect -16078 4644 -16074 4824
rect -16390 4624 -16074 4644
rect -14392 4825 -14064 4848
rect -14392 4645 -14382 4825
rect -14074 4645 -14064 4825
rect -14392 4622 -14064 4645
rect -12392 4827 -12068 4848
rect -12392 4647 -12384 4827
rect -12076 4647 -12068 4827
rect -12392 4626 -12068 4647
rect -10042 4822 -9722 4846
rect -10042 4642 -10036 4822
rect -9728 4642 -9722 4822
rect -10042 4618 -9722 4642
rect -8042 4820 -7724 4846
rect -8042 4640 -8037 4820
rect -7729 4640 -7724 4820
rect -8042 4614 -7724 4640
rect -6042 4820 -5722 4846
rect -6042 4640 -6036 4820
rect -5728 4640 -5722 4820
rect -6042 4614 -5722 4640
rect 2096 3787 2158 3802
rect 2096 3735 2101 3787
rect 2153 3735 2158 3787
rect 2096 3484 2158 3735
rect 4928 3769 4990 3784
rect 4928 3717 4933 3769
rect 4985 3717 4990 3769
rect 4602 3662 4696 3672
rect 4928 3666 4990 3717
rect 10018 3767 10080 3782
rect 10018 3715 10023 3767
rect 10075 3715 10080 3767
rect 8682 3666 8752 3686
rect 4928 3664 5082 3666
rect 5484 3664 8752 3666
rect 4928 3660 8752 3664
rect 4928 3634 8691 3660
rect 4928 3604 5383 3634
rect 4602 3558 4696 3568
rect 5364 3578 5383 3604
rect 5439 3608 8691 3634
rect 8743 3608 8752 3660
rect 5439 3604 8752 3608
rect 5439 3578 5458 3604
rect 8682 3582 8752 3604
rect 5364 3556 5458 3578
rect 2720 3484 2824 3500
rect 2096 3482 7194 3484
rect 1642 3472 1744 3482
rect 2096 3426 2744 3482
rect 2800 3479 7194 3482
rect 2800 3427 7127 3479
rect 7179 3427 7194 3479
rect 2800 3426 7194 3427
rect 2096 3422 7194 3426
rect 2720 3408 2824 3422
rect 8746 3408 8850 3418
rect 1642 3348 1744 3358
rect 8746 3352 8770 3408
rect 8826 3352 8850 3408
rect 8746 3342 8850 3352
rect 10018 3310 10080 3715
rect 11064 3771 11150 3790
rect 11064 3715 11079 3771
rect 11135 3715 11150 3771
rect 11064 3696 11150 3715
rect 13892 3483 13962 3500
rect 10394 3471 13148 3476
rect 10394 3419 10409 3471
rect 10461 3419 13081 3471
rect 13133 3419 13148 3471
rect 10394 3414 13148 3419
rect 13436 3464 13498 3474
rect 3648 3305 10080 3310
rect 3648 3253 3663 3305
rect 3715 3253 10080 3305
rect 3648 3248 10080 3253
rect 13436 3412 13441 3464
rect 13493 3412 13498 3464
rect 1404 3215 5680 3220
rect -11028 3160 -10924 3194
rect -17870 3142 -17754 3160
rect -17870 3140 -17840 3142
rect -17784 3140 -17754 3142
rect -17870 3086 -17840 3088
rect -17784 3086 -17754 3088
rect -17870 3068 -17754 3086
rect -11028 3104 -11004 3160
rect -10948 3104 -10924 3160
rect -11028 3070 -10924 3104
rect -4566 3153 -4458 3192
rect -4566 3097 -4540 3153
rect -4484 3097 -4458 3153
rect -4566 3058 -4458 3097
rect -4288 3174 -4078 3184
rect -4288 3074 -4280 3174
rect -4088 3074 -4078 3174
rect -4288 1808 -4078 3074
rect 1404 3163 5605 3215
rect 5657 3163 5680 3215
rect 1404 3158 5680 3163
rect 1404 3013 1466 3158
rect 7286 3156 7374 3168
rect 13436 3156 13498 3412
rect 13892 3427 13899 3483
rect 13955 3427 13962 3483
rect 13892 3410 13962 3427
rect 7286 3151 13498 3156
rect 7286 3099 7304 3151
rect 7356 3099 13498 3151
rect 7286 3094 13498 3099
rect 7286 3082 7374 3094
rect 1404 2961 1409 3013
rect 1461 2961 1466 3013
rect 1404 2946 1466 2961
rect 13576 2969 13632 2982
rect 13576 2900 13632 2913
rect -2396 2668 -2244 2678
rect 2540 2594 2828 2612
rect 2540 2592 2744 2594
rect 2540 2540 2570 2592
rect 2622 2540 2744 2592
rect 2540 2538 2744 2540
rect 2800 2538 2828 2594
rect 2540 2520 2828 2538
rect 5356 2594 5652 2612
rect 5356 2538 5384 2594
rect 5440 2592 5652 2594
rect 5440 2540 5570 2592
rect 5622 2540 5652 2592
rect 5440 2538 5652 2540
rect 5356 2520 5652 2538
rect 8540 2599 8856 2618
rect 8540 2597 8771 2599
rect 8540 2545 8571 2597
rect 8623 2545 8771 2597
rect 8540 2543 8771 2545
rect 8827 2543 8856 2599
rect 8540 2524 8856 2543
rect 11540 2570 11836 2588
rect 11540 2568 11752 2570
rect -2396 2496 -2244 2506
rect 11540 2516 11570 2568
rect 11622 2516 11752 2568
rect 11540 2514 11752 2516
rect 11808 2514 11836 2570
rect 11540 2496 11836 2514
rect -4288 1784 -2702 1808
rect -23116 1665 -22758 1678
rect -23116 1485 -23091 1665
rect -22783 1485 -22758 1665
rect -23116 1472 -22758 1485
rect -21116 1664 -20758 1676
rect -21116 1484 -21091 1664
rect -20783 1484 -20758 1664
rect -21116 1472 -20758 1484
rect -19116 1666 -18758 1678
rect -19116 1486 -19091 1666
rect -18783 1486 -18758 1666
rect -19116 1474 -18758 1486
rect -16634 1677 -16276 1690
rect -16634 1497 -16609 1677
rect -16301 1497 -16276 1677
rect -16634 1484 -16276 1497
rect -14432 1678 -14078 1690
rect -14432 1498 -14409 1678
rect -14101 1498 -14078 1678
rect -14432 1486 -14078 1498
rect -12032 1677 -11674 1690
rect -12032 1497 -12007 1677
rect -11699 1497 -11674 1677
rect -12032 1484 -11674 1497
rect -9432 1675 -9076 1688
rect -9432 1495 -9408 1675
rect -9100 1495 -9076 1675
rect -9432 1482 -9076 1495
rect -7432 1675 -7076 1688
rect -7432 1495 -7408 1675
rect -7100 1495 -7076 1675
rect -7432 1482 -7076 1495
rect -5434 1675 -5076 1688
rect -5434 1495 -5409 1675
rect -5101 1495 -5076 1675
rect -4288 1588 -2902 1784
rect -2708 1588 -2702 1784
rect -4288 1556 -2702 1588
rect 15056 1746 15236 7344
rect 16972 5487 17242 5510
rect 16972 5307 16985 5487
rect 17229 5307 17242 5487
rect 16972 5284 17242 5307
rect 18970 5484 19242 5510
rect 18970 5304 18984 5484
rect 19228 5304 19242 5484
rect 18970 5278 19242 5304
rect 20972 5484 21242 5510
rect 20972 5304 20985 5484
rect 21229 5304 21242 5484
rect 20972 5278 21242 5304
rect 23518 5483 23786 5508
rect 23518 5303 23530 5483
rect 23774 5303 23786 5483
rect 23518 5278 23786 5303
rect 25518 5484 25788 5510
rect 25518 5304 25531 5484
rect 25775 5304 25788 5484
rect 25518 5278 25788 5304
rect 27518 5483 27788 5508
rect 27518 5303 27531 5483
rect 27775 5303 27788 5483
rect 27518 5278 27788 5303
rect 16466 3822 16560 3856
rect 16466 3766 16485 3822
rect 16541 3766 16560 3822
rect 16466 3732 16560 3766
rect 22962 3820 23052 3854
rect 22962 3764 22979 3820
rect 23035 3764 23052 3820
rect 22962 3730 23052 3764
rect 17902 2339 18180 2352
rect 17902 2159 17919 2339
rect 18163 2159 18180 2339
rect 17902 2146 18180 2159
rect 19902 2339 20180 2352
rect 19902 2159 19919 2339
rect 20163 2159 20180 2339
rect 19902 2146 20180 2159
rect 21900 2339 22180 2352
rect 21900 2159 21918 2339
rect 22162 2159 22180 2339
rect 21900 2146 22180 2159
rect 23254 2336 23536 2348
rect 23254 2156 23273 2336
rect 23517 2156 23536 2336
rect 23254 2144 23536 2156
rect 25254 2337 25532 2350
rect 25254 2157 25271 2337
rect 25515 2157 25532 2337
rect 25254 2144 25532 2157
rect 15312 1948 16000 1966
rect 15312 1856 15324 1948
rect 15408 1856 16000 1948
rect 15312 1836 16000 1856
rect 15056 1672 15548 1746
rect 15056 1616 15469 1672
rect 15525 1616 15548 1672
rect 15056 1574 15548 1616
rect -4288 1554 -3222 1556
rect -5434 1482 -5076 1495
rect 2764 -15 2946 -10
rect 2764 -67 2779 -15
rect 2831 -67 2946 -15
rect 2764 -72 2946 -67
rect 2884 -462 2946 -72
rect 2884 -514 2889 -462
rect 2941 -514 2946 -462
rect 2884 -528 2946 -514
rect 5634 -11 5802 -6
rect 5634 -63 5735 -11
rect 5787 -63 5802 -11
rect 5634 -68 5802 -63
rect 8672 -25 8832 -20
rect 5634 -460 5696 -68
rect 5634 -512 5639 -460
rect 5691 -512 5696 -460
rect 5634 -526 5696 -512
rect 8672 -77 8765 -25
rect 8817 -77 8832 -25
rect 8672 -82 8832 -77
rect 11746 -25 11920 -20
rect 11746 -77 11853 -25
rect 11905 -77 11920 -25
rect 11746 -82 11920 -77
rect 8672 -460 8734 -82
rect 8672 -512 8677 -460
rect 8729 -512 8734 -460
rect 11746 -446 11808 -82
rect 11746 -498 11751 -446
rect 11803 -498 11808 -446
rect 11746 -512 11808 -498
rect 8672 -522 8734 -512
rect 15882 -528 16000 1836
rect 15622 -626 16000 -528
rect 15622 -934 15724 -626
rect 256 -962 696 -938
rect 256 -1270 258 -962
rect 694 -1270 696 -962
rect 256 -1294 696 -1270
rect 15410 -960 15762 -934
rect 15410 -1268 15432 -960
rect 15740 -1268 15762 -960
rect 15410 -1294 15762 -1268
rect 2228 -1468 2486 -1442
rect 2228 -1648 2235 -1468
rect 2479 -1648 2486 -1468
rect 2228 -1674 2486 -1648
rect 4228 -1468 4486 -1442
rect 4228 -1648 4235 -1468
rect 4479 -1648 4486 -1468
rect 4228 -1674 4486 -1648
rect 6228 -1468 6486 -1442
rect 6228 -1648 6235 -1468
rect 6479 -1648 6486 -1468
rect 6228 -1674 6486 -1648
rect 8446 -1475 8722 -1454
rect 8446 -1493 8476 -1475
rect 8692 -1493 8722 -1475
rect 8446 -1673 8462 -1493
rect 8706 -1673 8722 -1493
rect 8446 -1691 8476 -1673
rect 8692 -1691 8722 -1673
rect 10228 -1468 10486 -1442
rect 10228 -1648 10235 -1468
rect 10479 -1648 10486 -1468
rect 10228 -1674 10486 -1648
rect 12228 -1468 12486 -1442
rect 12228 -1648 12235 -1468
rect 12479 -1648 12486 -1468
rect 12228 -1674 12486 -1648
rect 14228 -1468 14486 -1442
rect 14228 -1648 14235 -1468
rect 14479 -1648 14486 -1468
rect 14228 -1674 14486 -1648
rect 8446 -1712 8722 -1691
<< via2 >>
rect -360 8831 -144 9047
rect 1640 8831 1856 9047
rect 3640 8831 3856 9047
rect 5640 8831 5856 9047
rect 7640 8831 7856 9047
rect 9640 8831 9856 9047
rect 11640 8831 11856 9047
rect 13640 8831 13856 9047
rect 15435 9066 15651 9084
rect 15435 8886 15651 9066
rect 15435 8868 15651 8886
rect -1329 7864 -793 8160
rect 15425 7857 15427 8153
rect 15427 7857 15799 8153
rect 15799 7857 15801 8153
rect -23000 4654 -22704 4790
rect -20996 4655 -20700 4791
rect -18998 4653 -18702 4789
rect -16380 4666 -16084 4802
rect -14376 4667 -14080 4803
rect -12378 4669 -12082 4805
rect -10030 4664 -9734 4800
rect -8031 4662 -7735 4798
rect -6030 4662 -5734 4798
rect 4602 3568 4696 3662
rect 5383 3578 5439 3634
rect 1642 3358 1744 3472
rect 2744 3426 2800 3482
rect 8770 3406 8826 3408
rect 8770 3354 8772 3406
rect 8772 3354 8824 3406
rect 8824 3354 8826 3406
rect 8770 3352 8826 3354
rect 11079 3769 11135 3771
rect 11079 3717 11081 3769
rect 11081 3717 11133 3769
rect 11133 3717 11135 3769
rect 11079 3715 11135 3717
rect -17840 3140 -17784 3142
rect -17840 3088 -17818 3140
rect -17818 3088 -17806 3140
rect -17806 3088 -17784 3140
rect -17840 3086 -17784 3088
rect -11004 3158 -10948 3160
rect -11004 3106 -11002 3158
rect -11002 3106 -10950 3158
rect -10950 3106 -10948 3158
rect -11004 3104 -10948 3106
rect -4540 3151 -4484 3153
rect -4540 3099 -4538 3151
rect -4538 3099 -4486 3151
rect -4486 3099 -4484 3151
rect -4540 3097 -4484 3099
rect -4280 3074 -4088 3174
rect 13899 3481 13955 3483
rect 13899 3429 13901 3481
rect 13901 3429 13953 3481
rect 13953 3429 13955 3481
rect 13899 3427 13955 3429
rect 13576 2967 13632 2969
rect 13576 2915 13578 2967
rect 13578 2915 13630 2967
rect 13630 2915 13632 2967
rect 13576 2913 13632 2915
rect -2396 2506 -2244 2668
rect 2744 2538 2800 2594
rect 5384 2538 5440 2594
rect 8771 2543 8827 2599
rect 11752 2514 11808 2570
rect -23085 1507 -22789 1643
rect -21085 1506 -20789 1642
rect -19085 1508 -18789 1644
rect -16603 1519 -16307 1655
rect -14403 1520 -14107 1656
rect -12001 1519 -11705 1655
rect -9402 1517 -9106 1653
rect -7402 1517 -7106 1653
rect -5403 1517 -5107 1653
rect -2902 1588 -2708 1784
rect 16999 5329 17215 5465
rect 18998 5326 19214 5462
rect 20999 5326 21215 5462
rect 23544 5325 23760 5461
rect 25545 5326 25761 5462
rect 27545 5325 27761 5461
rect 16485 3820 16541 3822
rect 16485 3768 16487 3820
rect 16487 3768 16539 3820
rect 16539 3768 16541 3820
rect 16485 3766 16541 3768
rect 22979 3818 23035 3820
rect 22979 3766 22981 3818
rect 22981 3766 23033 3818
rect 23033 3766 23035 3818
rect 22979 3764 23035 3766
rect 17933 2181 18149 2317
rect 19933 2181 20149 2317
rect 21932 2181 22148 2317
rect 23287 2178 23503 2314
rect 25285 2179 25501 2315
rect 15469 1670 15525 1672
rect 15469 1618 15471 1670
rect 15471 1618 15523 1670
rect 15523 1618 15525 1670
rect 15469 1616 15525 1618
rect 288 -1264 664 -968
rect 15438 -1262 15734 -966
rect 2249 -1626 2465 -1490
rect 4249 -1626 4465 -1490
rect 6249 -1626 6465 -1490
rect 8476 -1493 8692 -1475
rect 8476 -1673 8692 -1493
rect 8476 -1691 8692 -1673
rect 10249 -1626 10465 -1490
rect 12249 -1626 12465 -1490
rect 14249 -1626 14465 -1490
<< metal3 >>
rect 15404 9088 15682 9095
rect -392 9051 -112 9079
rect -392 8827 -364 9051
rect -140 8827 -112 9051
rect -392 8799 -112 8827
rect 1608 9051 1888 9079
rect 1608 8827 1636 9051
rect 1860 8827 1888 9051
rect 1608 8799 1888 8827
rect 3608 9051 3888 9079
rect 3608 8827 3636 9051
rect 3860 8827 3888 9051
rect 3608 8799 3888 8827
rect 5608 9051 5888 9079
rect 5608 8827 5636 9051
rect 5860 8827 5888 9051
rect 5608 8799 5888 8827
rect 7608 9051 7888 9079
rect 7608 8827 7636 9051
rect 7860 8827 7888 9051
rect 7608 8799 7888 8827
rect 9608 9051 9888 9079
rect 9608 8827 9636 9051
rect 9860 8827 9888 9051
rect 9608 8799 9888 8827
rect 11608 9051 11888 9079
rect 11608 8827 11636 9051
rect 11860 8827 11888 9051
rect 11608 8799 11888 8827
rect 13608 9051 13888 9079
rect 13608 8827 13636 9051
rect 13860 8827 13888 9051
rect 15404 8864 15431 9088
rect 15655 8864 15682 9088
rect 15404 8857 15682 8864
rect 13608 8799 13888 8827
rect -1360 8164 -762 8187
rect -1360 7860 -1333 8164
rect -789 7860 -762 8164
rect -1360 7837 -762 7860
rect 15394 8157 15832 8183
rect 15394 7853 15421 8157
rect 15805 7853 15832 8157
rect 15394 7827 15832 7853
rect -11014 6072 -3734 6138
rect -23016 4794 -22688 4817
rect -23016 4650 -23004 4794
rect -22700 4650 -22688 4794
rect -23016 4627 -22688 4650
rect -21020 4795 -20676 4831
rect -21020 4651 -21000 4795
rect -20696 4651 -20676 4795
rect -21020 4615 -20676 4651
rect -19020 4793 -18680 4831
rect -19020 4649 -19002 4793
rect -18698 4649 -18680 4793
rect -19020 4611 -18680 4649
rect -16400 4806 -16064 4839
rect -16400 4662 -16384 4806
rect -16080 4662 -16064 4806
rect -16400 4629 -16064 4662
rect -14402 4807 -14054 4843
rect -14402 4663 -14380 4807
rect -14076 4663 -14054 4807
rect -14402 4627 -14054 4663
rect -12402 4809 -12058 4843
rect -12402 4665 -12382 4809
rect -12078 4665 -12058 4809
rect -12402 4631 -12058 4665
rect -11014 3189 -10892 6072
rect -10052 4804 -9712 4841
rect -10052 4660 -10034 4804
rect -9730 4660 -9712 4804
rect -10052 4623 -9712 4660
rect -8052 4802 -7714 4841
rect -8052 4658 -8035 4802
rect -7731 4658 -7714 4802
rect -8052 4619 -7714 4658
rect -6052 4802 -5712 4841
rect -6052 4658 -6034 4802
rect -5730 4658 -5712 4802
rect -6052 4619 -5712 4658
rect -3806 3650 -3734 6072
rect 16962 5469 17252 5505
rect 16962 5325 16995 5469
rect 17219 5325 17252 5469
rect 16962 5289 17252 5325
rect 18960 5466 19252 5505
rect 18960 5322 18994 5466
rect 19218 5322 19252 5466
rect 18960 5283 19252 5322
rect 20962 5466 21252 5505
rect 20962 5322 20995 5466
rect 21219 5322 21252 5466
rect 20962 5283 21252 5322
rect 23508 5465 23796 5503
rect 23508 5321 23540 5465
rect 23764 5321 23796 5465
rect 23508 5283 23796 5321
rect 25508 5466 25798 5505
rect 25508 5322 25541 5466
rect 25765 5322 25798 5466
rect 25508 5283 25798 5322
rect 27508 5465 27798 5503
rect 27508 5321 27541 5465
rect 27765 5321 27798 5465
rect 27508 5283 27798 5321
rect 16248 3846 16314 3848
rect 16456 3846 16570 3851
rect 16248 3822 16570 3846
rect 11054 3780 11160 3785
rect 11726 3780 11832 3782
rect 11054 3771 11832 3780
rect 11054 3715 11079 3771
rect 11135 3715 11832 3771
rect 11054 3706 11832 3715
rect 11054 3701 11160 3706
rect 4592 3662 4706 3667
rect 4592 3650 4602 3662
rect -3806 3584 4602 3650
rect 4592 3568 4602 3584
rect 4696 3568 4706 3662
rect 5360 3651 5464 3672
rect 4592 3563 4706 3568
rect 5354 3634 5468 3651
rect 5354 3578 5383 3634
rect 5439 3578 5468 3634
rect 5354 3561 5468 3578
rect 2710 3482 2834 3495
rect 1632 3472 1754 3477
rect -11038 3160 -10892 3189
rect -17880 3142 -17744 3155
rect -17880 3086 -17840 3142
rect -17784 3086 -17744 3142
rect -17880 3073 -17744 3086
rect -11038 3104 -11004 3160
rect -10948 3104 -10892 3160
rect -11038 3082 -10892 3104
rect -10706 3358 1642 3472
rect 1744 3358 1754 3472
rect 2710 3426 2744 3482
rect 2800 3426 2834 3482
rect 2710 3413 2834 3426
rect -11038 3075 -10914 3082
rect -17870 2926 -17754 3073
rect -10706 2926 -10576 3358
rect 1632 3353 1754 3358
rect -4576 3182 -4448 3187
rect -4576 3180 -4274 3182
rect -102 3180 150 3184
rect 2720 3180 2824 3413
rect -4576 3174 -4032 3180
rect -4576 3153 -4280 3174
rect -4576 3097 -4540 3153
rect -4484 3097 -4280 3153
rect -4576 3074 -4280 3097
rect -4088 3074 -4032 3174
rect -4576 3068 -4032 3074
rect -102 3068 2824 3180
rect -4576 3063 -4448 3068
rect -17870 2798 -10576 2926
rect -3674 2668 -2176 2704
rect -3674 2506 -2396 2668
rect -2244 2506 -2176 2668
rect -3674 2474 -2176 2506
rect -23126 1647 -22748 1673
rect -23126 1503 -23089 1647
rect -22785 1503 -22748 1647
rect -23126 1477 -22748 1503
rect -21126 1646 -20748 1671
rect -21126 1502 -21089 1646
rect -20785 1502 -20748 1646
rect -21126 1477 -20748 1502
rect -19126 1648 -18748 1673
rect -19126 1504 -19089 1648
rect -18785 1504 -18748 1648
rect -19126 1479 -18748 1504
rect -16644 1659 -16266 1685
rect -16644 1515 -16607 1659
rect -16303 1515 -16266 1659
rect -16644 1489 -16266 1515
rect -14442 1660 -14068 1685
rect -14442 1516 -14407 1660
rect -14103 1516 -14068 1660
rect -14442 1491 -14068 1516
rect -12042 1659 -11664 1685
rect -12042 1515 -12005 1659
rect -11701 1515 -11664 1659
rect -12042 1489 -11664 1515
rect -9442 1657 -9066 1683
rect -9442 1513 -9406 1657
rect -9102 1513 -9066 1657
rect -9442 1487 -9066 1513
rect -7442 1657 -7066 1683
rect -7442 1513 -7406 1657
rect -7102 1513 -7066 1657
rect -7442 1487 -7066 1513
rect -5444 1657 -5066 1683
rect -5444 1513 -5407 1657
rect -5103 1513 -5066 1657
rect -5444 1487 -5066 1513
rect -3654 -5908 -3374 2474
rect -2912 1784 -2698 1789
rect -2912 1588 -2902 1784
rect -2708 1780 -2698 1784
rect -102 1780 150 3068
rect 2720 2616 2824 3068
rect 2721 2594 2823 2616
rect 2721 2538 2744 2594
rect 2800 2538 2823 2594
rect 5360 2594 5464 3561
rect 8746 3413 8852 3414
rect 8736 3408 8860 3413
rect 8736 3352 8770 3408
rect 8826 3352 8860 3408
rect 8736 3347 8860 3352
rect 8746 2624 8852 3347
rect 5360 2582 5384 2594
rect 2721 2510 2823 2538
rect 5361 2538 5384 2582
rect 5440 2582 5464 2594
rect 8747 2599 8851 2624
rect 5440 2538 5463 2582
rect 5361 2510 5463 2538
rect 8747 2543 8771 2599
rect 8827 2543 8851 2599
rect 11728 2590 11832 3706
rect 16248 3766 16485 3822
rect 16541 3766 16570 3822
rect 16248 3742 16570 3766
rect 13882 3490 13972 3495
rect 16248 3490 16314 3742
rect 16456 3737 16570 3742
rect 22900 3849 23054 3862
rect 22900 3820 23062 3849
rect 22900 3764 22979 3820
rect 23035 3764 23062 3820
rect 13882 3483 16314 3490
rect 13882 3427 13899 3483
rect 13955 3427 16314 3483
rect 13882 3420 16314 3427
rect 22900 3735 23062 3764
rect 13882 3415 13972 3420
rect 16186 3076 16320 3078
rect 22900 3076 23054 3735
rect 13560 3000 16320 3076
rect 22892 3000 23054 3076
rect 13560 2969 13648 3000
rect 13560 2913 13576 2969
rect 13632 2913 13648 2969
rect 13560 2890 13648 2913
rect 8747 2514 8851 2543
rect 11729 2570 11831 2590
rect 11729 2514 11752 2570
rect 11808 2514 11831 2570
rect 11729 2486 11831 2514
rect 16186 2088 16320 3000
rect 17892 2321 18190 2347
rect 17892 2177 17929 2321
rect 18153 2177 18190 2321
rect 17892 2151 18190 2177
rect 19892 2321 20190 2347
rect 19892 2177 19929 2321
rect 20153 2177 20190 2321
rect 19892 2151 20190 2177
rect 21890 2321 22190 2347
rect 21890 2177 21928 2321
rect 22152 2177 22190 2321
rect 21890 2151 22190 2177
rect 22900 2088 23054 3000
rect 23244 2318 23546 2343
rect 23244 2174 23283 2318
rect 23507 2174 23546 2318
rect 23244 2149 23546 2174
rect 25244 2319 25542 2345
rect 25244 2175 25281 2319
rect 25505 2175 25542 2319
rect 25244 2149 25542 2175
rect 16186 1968 23054 2088
rect 16186 1966 23016 1968
rect -2708 1592 150 1780
rect 16674 1746 16684 1788
rect 15442 1672 16684 1746
rect 15442 1616 15469 1672
rect 15525 1616 16684 1672
rect -2708 1588 76 1592
rect -2912 1583 -2698 1588
rect 15442 1574 16684 1616
rect 15446 1572 16684 1574
rect 16674 1514 16684 1572
rect 16968 1514 16978 1788
rect 246 -964 706 -943
rect 246 -1268 284 -964
rect 668 -1268 706 -964
rect 246 -1289 706 -1268
rect 15400 -962 15772 -939
rect 15400 -1266 15434 -962
rect 15738 -1266 15772 -962
rect 15400 -1289 15772 -1266
rect 2218 -1486 2496 -1447
rect 2218 -1630 2245 -1486
rect 2469 -1630 2496 -1486
rect 2218 -1669 2496 -1630
rect 4218 -1486 4496 -1447
rect 4218 -1630 4245 -1486
rect 4469 -1630 4496 -1486
rect 4218 -1669 4496 -1630
rect 6218 -1486 6496 -1447
rect 6218 -1630 6245 -1486
rect 6469 -1630 6496 -1486
rect 6218 -1669 6496 -1630
rect 8436 -1471 8732 -1459
rect 8436 -1695 8472 -1471
rect 8696 -1695 8732 -1471
rect 10218 -1486 10496 -1447
rect 10218 -1630 10245 -1486
rect 10469 -1630 10496 -1486
rect 10218 -1669 10496 -1630
rect 12218 -1486 12496 -1447
rect 12218 -1630 12245 -1486
rect 12469 -1630 12496 -1486
rect 12218 -1669 12496 -1630
rect 14218 -1486 14496 -1447
rect 14218 -1630 14245 -1486
rect 14469 -1630 14496 -1486
rect 14218 -1669 14496 -1630
rect 8436 -1707 8732 -1695
<< via3 >>
rect -364 9047 -140 9051
rect -364 8831 -360 9047
rect -360 8831 -144 9047
rect -144 8831 -140 9047
rect -364 8827 -140 8831
rect 1636 9047 1860 9051
rect 1636 8831 1640 9047
rect 1640 8831 1856 9047
rect 1856 8831 1860 9047
rect 1636 8827 1860 8831
rect 3636 9047 3860 9051
rect 3636 8831 3640 9047
rect 3640 8831 3856 9047
rect 3856 8831 3860 9047
rect 3636 8827 3860 8831
rect 5636 9047 5860 9051
rect 5636 8831 5640 9047
rect 5640 8831 5856 9047
rect 5856 8831 5860 9047
rect 5636 8827 5860 8831
rect 7636 9047 7860 9051
rect 7636 8831 7640 9047
rect 7640 8831 7856 9047
rect 7856 8831 7860 9047
rect 7636 8827 7860 8831
rect 9636 9047 9860 9051
rect 9636 8831 9640 9047
rect 9640 8831 9856 9047
rect 9856 8831 9860 9047
rect 9636 8827 9860 8831
rect 11636 9047 11860 9051
rect 11636 8831 11640 9047
rect 11640 8831 11856 9047
rect 11856 8831 11860 9047
rect 11636 8827 11860 8831
rect 13636 9047 13860 9051
rect 13636 8831 13640 9047
rect 13640 8831 13856 9047
rect 13856 8831 13860 9047
rect 13636 8827 13860 8831
rect 15431 9084 15655 9088
rect 15431 8868 15435 9084
rect 15435 8868 15651 9084
rect 15651 8868 15655 9084
rect 15431 8864 15655 8868
rect -1333 8160 -789 8164
rect -1333 7864 -1329 8160
rect -1329 7864 -793 8160
rect -793 7864 -789 8160
rect -1333 7860 -789 7864
rect 15421 8153 15805 8157
rect 15421 7857 15425 8153
rect 15425 7857 15801 8153
rect 15801 7857 15805 8153
rect 15421 7853 15805 7857
rect -23004 4790 -22700 4794
rect -23004 4654 -23000 4790
rect -23000 4654 -22704 4790
rect -22704 4654 -22700 4790
rect -23004 4650 -22700 4654
rect -21000 4791 -20696 4795
rect -21000 4655 -20996 4791
rect -20996 4655 -20700 4791
rect -20700 4655 -20696 4791
rect -21000 4651 -20696 4655
rect -19002 4789 -18698 4793
rect -19002 4653 -18998 4789
rect -18998 4653 -18702 4789
rect -18702 4653 -18698 4789
rect -19002 4649 -18698 4653
rect -16384 4802 -16080 4806
rect -16384 4666 -16380 4802
rect -16380 4666 -16084 4802
rect -16084 4666 -16080 4802
rect -16384 4662 -16080 4666
rect -14380 4803 -14076 4807
rect -14380 4667 -14376 4803
rect -14376 4667 -14080 4803
rect -14080 4667 -14076 4803
rect -14380 4663 -14076 4667
rect -12382 4805 -12078 4809
rect -12382 4669 -12378 4805
rect -12378 4669 -12082 4805
rect -12082 4669 -12078 4805
rect -12382 4665 -12078 4669
rect -10034 4800 -9730 4804
rect -10034 4664 -10030 4800
rect -10030 4664 -9734 4800
rect -9734 4664 -9730 4800
rect -10034 4660 -9730 4664
rect -8035 4798 -7731 4802
rect -8035 4662 -8031 4798
rect -8031 4662 -7735 4798
rect -7735 4662 -7731 4798
rect -8035 4658 -7731 4662
rect -6034 4798 -5730 4802
rect -6034 4662 -6030 4798
rect -6030 4662 -5734 4798
rect -5734 4662 -5730 4798
rect -6034 4658 -5730 4662
rect 16995 5465 17219 5469
rect 16995 5329 16999 5465
rect 16999 5329 17215 5465
rect 17215 5329 17219 5465
rect 16995 5325 17219 5329
rect 18994 5462 19218 5466
rect 18994 5326 18998 5462
rect 18998 5326 19214 5462
rect 19214 5326 19218 5462
rect 18994 5322 19218 5326
rect 20995 5462 21219 5466
rect 20995 5326 20999 5462
rect 20999 5326 21215 5462
rect 21215 5326 21219 5462
rect 20995 5322 21219 5326
rect 23540 5461 23764 5465
rect 23540 5325 23544 5461
rect 23544 5325 23760 5461
rect 23760 5325 23764 5461
rect 23540 5321 23764 5325
rect 25541 5462 25765 5466
rect 25541 5326 25545 5462
rect 25545 5326 25761 5462
rect 25761 5326 25765 5462
rect 25541 5322 25765 5326
rect 27541 5461 27765 5465
rect 27541 5325 27545 5461
rect 27545 5325 27761 5461
rect 27761 5325 27765 5461
rect 27541 5321 27765 5325
rect -23089 1643 -22785 1647
rect -23089 1507 -23085 1643
rect -23085 1507 -22789 1643
rect -22789 1507 -22785 1643
rect -23089 1503 -22785 1507
rect -21089 1642 -20785 1646
rect -21089 1506 -21085 1642
rect -21085 1506 -20789 1642
rect -20789 1506 -20785 1642
rect -21089 1502 -20785 1506
rect -19089 1644 -18785 1648
rect -19089 1508 -19085 1644
rect -19085 1508 -18789 1644
rect -18789 1508 -18785 1644
rect -19089 1504 -18785 1508
rect -16607 1655 -16303 1659
rect -16607 1519 -16603 1655
rect -16603 1519 -16307 1655
rect -16307 1519 -16303 1655
rect -16607 1515 -16303 1519
rect -14407 1656 -14103 1660
rect -14407 1520 -14403 1656
rect -14403 1520 -14107 1656
rect -14107 1520 -14103 1656
rect -14407 1516 -14103 1520
rect -12005 1655 -11701 1659
rect -12005 1519 -12001 1655
rect -12001 1519 -11705 1655
rect -11705 1519 -11701 1655
rect -12005 1515 -11701 1519
rect -9406 1653 -9102 1657
rect -9406 1517 -9402 1653
rect -9402 1517 -9106 1653
rect -9106 1517 -9102 1653
rect -9406 1513 -9102 1517
rect -7406 1653 -7102 1657
rect -7406 1517 -7402 1653
rect -7402 1517 -7106 1653
rect -7106 1517 -7102 1653
rect -7406 1513 -7102 1517
rect -5407 1653 -5103 1657
rect -5407 1517 -5403 1653
rect -5403 1517 -5107 1653
rect -5107 1517 -5103 1653
rect -5407 1513 -5103 1517
rect 17929 2317 18153 2321
rect 17929 2181 17933 2317
rect 17933 2181 18149 2317
rect 18149 2181 18153 2317
rect 17929 2177 18153 2181
rect 19929 2317 20153 2321
rect 19929 2181 19933 2317
rect 19933 2181 20149 2317
rect 20149 2181 20153 2317
rect 19929 2177 20153 2181
rect 21928 2317 22152 2321
rect 21928 2181 21932 2317
rect 21932 2181 22148 2317
rect 22148 2181 22152 2317
rect 21928 2177 22152 2181
rect 23283 2314 23507 2318
rect 23283 2178 23287 2314
rect 23287 2178 23503 2314
rect 23503 2178 23507 2314
rect 23283 2174 23507 2178
rect 25281 2315 25505 2319
rect 25281 2179 25285 2315
rect 25285 2179 25501 2315
rect 25501 2179 25505 2315
rect 25281 2175 25505 2179
rect 16684 1514 16968 1788
rect 284 -968 668 -964
rect 284 -1264 288 -968
rect 288 -1264 664 -968
rect 664 -1264 668 -968
rect 284 -1268 668 -1264
rect 15434 -966 15738 -962
rect 15434 -1262 15438 -966
rect 15438 -1262 15734 -966
rect 15734 -1262 15738 -966
rect 15434 -1266 15738 -1262
rect 2245 -1490 2469 -1486
rect 2245 -1626 2249 -1490
rect 2249 -1626 2465 -1490
rect 2465 -1626 2469 -1490
rect 2245 -1630 2469 -1626
rect 4245 -1490 4469 -1486
rect 4245 -1626 4249 -1490
rect 4249 -1626 4465 -1490
rect 4465 -1626 4469 -1490
rect 4245 -1630 4469 -1626
rect 6245 -1490 6469 -1486
rect 6245 -1626 6249 -1490
rect 6249 -1626 6465 -1490
rect 6465 -1626 6469 -1490
rect 6245 -1630 6469 -1626
rect 8472 -1475 8696 -1471
rect 8472 -1691 8476 -1475
rect 8476 -1691 8692 -1475
rect 8692 -1691 8696 -1475
rect 8472 -1695 8696 -1691
rect 10245 -1490 10469 -1486
rect 10245 -1626 10249 -1490
rect 10249 -1626 10465 -1490
rect 10465 -1626 10469 -1490
rect 10245 -1630 10469 -1626
rect 12245 -1490 12469 -1486
rect 12245 -1626 12249 -1490
rect 12249 -1626 12465 -1490
rect 12465 -1626 12469 -1490
rect 12245 -1630 12469 -1626
rect 14245 -1490 14469 -1486
rect 14245 -1626 14249 -1490
rect 14249 -1626 14465 -1490
rect 14465 -1626 14469 -1490
rect 14245 -1630 14469 -1626
<< metal4 >>
rect -812 9088 16212 9458
rect -812 9051 15431 9088
rect -812 8827 -364 9051
rect -140 8827 1636 9051
rect 1860 8827 3636 9051
rect 3860 8827 5636 9051
rect 5860 8827 7636 9051
rect 7860 8827 9636 9051
rect 9860 8827 11636 9051
rect 11860 8827 13636 9051
rect 13860 8864 15431 9051
rect 15655 8864 16212 9088
rect 13860 8827 16212 8864
rect -812 8632 16212 8827
rect -1351 8178 -771 8183
rect 15403 8178 15823 8179
rect -23322 8164 -768 8178
rect -23322 7860 -1333 8164
rect -789 7860 -768 8164
rect -23322 7838 -768 7860
rect 15403 8157 28998 8178
rect 15403 7853 15421 8157
rect 15805 7853 28998 8157
rect -23008 4794 -22688 7838
rect -21008 4827 -20688 7838
rect -19008 4827 -18688 7838
rect -16390 4835 -16070 7838
rect -14390 4839 -14070 7838
rect -12390 4839 -12070 7838
rect -23008 4732 -23004 4794
rect -23007 4650 -23004 4732
rect -22700 4732 -22688 4794
rect -21011 4795 -20685 4827
rect -22700 4650 -22697 4732
rect -23007 4631 -22697 4650
rect -21011 4651 -21000 4795
rect -20696 4651 -20685 4795
rect -21011 4619 -20685 4651
rect -19011 4793 -18688 4827
rect -19011 4649 -19002 4793
rect -18698 4732 -18688 4793
rect -16391 4806 -16070 4835
rect -18698 4649 -18689 4732
rect -19011 4615 -18689 4649
rect -16391 4662 -16384 4806
rect -16080 4718 -16070 4806
rect -14393 4807 -14063 4839
rect -16080 4662 -16073 4718
rect -16391 4633 -16073 4662
rect -14393 4663 -14380 4807
rect -14076 4663 -14063 4807
rect -14393 4631 -14063 4663
rect -12393 4809 -12067 4839
rect -10042 4837 -9722 7838
rect -8042 4837 -7722 7838
rect -6042 4837 -5722 7838
rect 15403 7831 28998 7853
rect 15708 7830 28998 7831
rect 16972 5501 17242 7830
rect 18972 5501 19242 7830
rect 20972 5501 21242 7830
rect 16971 5469 17243 5501
rect 16971 5325 16995 5469
rect 17219 5325 17243 5469
rect 16971 5293 17243 5325
rect 18969 5466 19243 5501
rect 18969 5322 18994 5466
rect 19218 5322 19243 5466
rect 18969 5287 19243 5322
rect 20971 5466 21243 5501
rect 23518 5499 23788 7830
rect 25518 5501 25788 7830
rect 20971 5322 20995 5466
rect 21219 5322 21243 5466
rect 20971 5287 21243 5322
rect 23517 5465 23788 5499
rect 23517 5321 23540 5465
rect 23764 5321 23788 5465
rect 23517 5298 23788 5321
rect 25517 5466 25789 5501
rect 27518 5499 27788 7830
rect 25517 5322 25541 5466
rect 25765 5322 25789 5466
rect 23517 5287 23787 5298
rect 25517 5287 25789 5322
rect 27517 5465 27789 5499
rect 27517 5321 27541 5465
rect 27765 5321 27789 5465
rect 27517 5287 27789 5321
rect -12393 4665 -12382 4809
rect -12078 4665 -12067 4809
rect -12393 4635 -12067 4665
rect -10043 4804 -9721 4837
rect -10043 4660 -10034 4804
rect -9730 4660 -9721 4804
rect -10043 4627 -9721 4660
rect -8043 4802 -7722 4837
rect -8043 4658 -8035 4802
rect -7731 4692 -7722 4802
rect -6043 4802 -5721 4837
rect -7731 4658 -7723 4692
rect -8043 4623 -7723 4658
rect -6043 4658 -6034 4802
rect -5730 4658 -5721 4802
rect -6043 4623 -5721 4658
rect 17901 2321 18181 2343
rect 17901 2177 17929 2321
rect 18153 2177 18181 2321
rect 17901 2155 18181 2177
rect 19901 2321 20181 2343
rect 19901 2177 19929 2321
rect 20153 2177 20181 2321
rect 19901 2155 20181 2177
rect 21899 2321 22181 2343
rect 21899 2177 21928 2321
rect 22152 2177 22181 2321
rect 21899 2155 22181 2177
rect 23253 2318 23537 2339
rect 23253 2174 23283 2318
rect 23507 2174 23537 2318
rect 16683 1788 16969 1789
rect -16632 1681 -16276 1688
rect -14432 1681 -14076 1688
rect -12032 1681 -11676 1688
rect -23117 1647 -22757 1669
rect -23117 1503 -23089 1647
rect -22785 1503 -22757 1647
rect -23117 1481 -22757 1503
rect -21117 1646 -20757 1667
rect -21117 1502 -21089 1646
rect -20785 1502 -20757 1646
rect -21117 1481 -20757 1502
rect -19117 1648 -18757 1669
rect -19117 1504 -19089 1648
rect -18785 1504 -18757 1648
rect -19117 1483 -18757 1504
rect -16635 1659 -16275 1681
rect -16635 1515 -16607 1659
rect -16303 1515 -16275 1659
rect -16635 1493 -16275 1515
rect -14433 1660 -14076 1681
rect -14433 1516 -14407 1660
rect -14103 1516 -14076 1660
rect -14433 1495 -14076 1516
rect -23114 -942 -22758 1481
rect -21114 -942 -20758 1481
rect -19114 -942 -18758 1483
rect -16632 -942 -16276 1493
rect -14432 -942 -14076 1495
rect -12033 1659 -11673 1681
rect -9432 1679 -9076 1688
rect -7432 1679 -7076 1688
rect -5432 1679 -5076 1688
rect -12033 1515 -12005 1659
rect -11701 1515 -11673 1659
rect -12033 1493 -11673 1515
rect -9433 1657 -9075 1679
rect -9433 1513 -9406 1657
rect -9102 1513 -9075 1657
rect -12032 -942 -11676 1493
rect -9433 1491 -9075 1513
rect -7433 1657 -7075 1679
rect -7433 1513 -7406 1657
rect -7102 1513 -7075 1657
rect -7433 1491 -7075 1513
rect -5435 1657 -5075 1679
rect -5435 1513 -5407 1657
rect -5103 1513 -5075 1657
rect 16683 1514 16684 1788
rect 16968 1514 16969 1788
rect 16683 1513 16969 1514
rect -5435 1491 -5075 1513
rect -9432 -942 -9076 1491
rect -7432 -942 -7076 1491
rect -5432 -942 -5076 1491
rect -23322 -946 -1350 -942
rect -23322 -947 696 -946
rect -23322 -964 697 -947
rect -23322 -1268 284 -964
rect 668 -1268 697 -964
rect -23322 -1282 697 -1268
rect 255 -1285 697 -1282
rect 15409 -950 15763 -943
rect 17902 -950 18180 2155
rect 19902 -950 20180 2155
rect 21902 -950 22180 2155
rect 23253 2153 23537 2174
rect 25253 2319 25533 2341
rect 25253 2175 25281 2319
rect 25505 2288 25533 2319
rect 25505 2175 25534 2288
rect 25253 2153 25534 2175
rect 23256 -950 23534 2153
rect 25256 -950 25534 2153
rect 27256 -950 27534 2288
rect 15409 -962 28996 -950
rect 15409 -1266 15434 -962
rect 15738 -1266 28996 -962
rect 15409 -1284 28996 -1266
rect 15409 -1285 15763 -1284
rect 1530 -1471 15894 -1398
rect 1530 -1486 8472 -1471
rect 1530 -1630 2245 -1486
rect 2469 -1630 4245 -1486
rect 4469 -1630 6245 -1486
rect 6469 -1630 8472 -1486
rect 1530 -1695 8472 -1630
rect 8696 -1486 15894 -1471
rect 8696 -1630 10245 -1486
rect 10469 -1630 12245 -1486
rect 12469 -1630 14245 -1486
rect 14469 -1630 15894 -1486
rect 8696 -1695 15894 -1630
rect 1530 -2150 15894 -1695
<< via4 >>
rect 16684 1514 16968 1788
<< metal5 >>
rect 16624 1788 17748 1860
rect 16624 1514 16684 1788
rect 16968 1514 17748 1788
rect 16624 1432 17748 1514
rect 17304 -5146 17748 1432
<< labels >>
rlabel metal1 -17754 3120 -17754 3120 4 Buff_VCO_4/IN
rlabel metal1 22948 3792 22948 3792 4 Buff_VCO_1/IN
rlabel metal1 -10924 3132 -10924 3132 4 Buff_VCO_3/IN
rlabel metal1 -4458 3130 -4458 3130 4 Buff_VCO_2/IN
rlabel metal1 16460 3794 16460 3794 4 Buff_VCO_0/IN
rlabel metal4 7152 8932 7152 8932 4 VP
port 1 se
rlabel metal4 11374 -1581 11374 -1581 4 VN
port 4 se
rlabel metal5 17512 -3998 17512 -3998 1 VCT
port 2 n
rlabel metal3 -3550 -3396 -3550 -3396 1 VB
port 5 n
rlabel metal1 -24636 -3264 -24636 -3264 5 OUT_5
port 9 s
rlabel metal1 -17158 -3270 -17158 -3270 5 OUT_4
port 6 s
rlabel metal1 -10482 -3348 -10482 -3348 5 OUT_3
port 7 s
rlabel metal1 22642 -2778 22642 -2778 5 OUT_1
port 3 s
rlabel metal1 29354 -2726 29354 -2726 5 OUT_2
port 8 s
<< end >>
