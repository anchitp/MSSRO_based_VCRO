magic
tech sky130A
magscale 1 2
timestamp 1636370378
<< error_p >>
rect -845 662 -787 668
rect -845 628 -833 662
rect -845 622 -787 628
<< nmos >>
rect -927 -500 -897 500
rect -831 -500 -801 500
rect -735 -500 -705 500
rect -639 -500 -609 500
rect -543 -500 -513 500
rect -447 -500 -417 500
rect -351 -500 -321 500
rect -255 -500 -225 500
rect -159 -500 -129 500
rect -63 -500 -33 500
rect 33 -500 63 500
rect 129 -500 159 500
rect 225 -500 255 500
rect 321 -500 351 500
rect 417 -500 447 500
rect 513 -500 543 500
rect 609 -500 639 500
rect 705 -500 735 500
rect 801 -500 831 500
rect 897 -500 927 500
<< ndiff >>
rect -989 488 -927 500
rect -989 -488 -977 488
rect -943 -488 -927 488
rect -989 -500 -927 -488
rect -897 488 -831 500
rect -897 -488 -881 488
rect -847 -488 -831 488
rect -897 -500 -831 -488
rect -801 488 -735 500
rect -801 -488 -785 488
rect -751 -488 -735 488
rect -801 -500 -735 -488
rect -705 488 -639 500
rect -705 -488 -689 488
rect -655 -488 -639 488
rect -705 -500 -639 -488
rect -609 488 -543 500
rect -609 -488 -593 488
rect -559 -488 -543 488
rect -609 -500 -543 -488
rect -513 488 -447 500
rect -513 -488 -497 488
rect -463 -488 -447 488
rect -513 -500 -447 -488
rect -417 488 -351 500
rect -417 -488 -401 488
rect -367 -488 -351 488
rect -417 -500 -351 -488
rect -321 488 -255 500
rect -321 -488 -305 488
rect -271 -488 -255 488
rect -321 -500 -255 -488
rect -225 488 -159 500
rect -225 -488 -209 488
rect -175 -488 -159 488
rect -225 -500 -159 -488
rect -129 488 -63 500
rect -129 -488 -113 488
rect -79 -488 -63 488
rect -129 -500 -63 -488
rect -33 488 33 500
rect -33 -488 -17 488
rect 17 -488 33 488
rect -33 -500 33 -488
rect 63 488 129 500
rect 63 -488 79 488
rect 113 -488 129 488
rect 63 -500 129 -488
rect 159 488 225 500
rect 159 -488 175 488
rect 209 -488 225 488
rect 159 -500 225 -488
rect 255 488 321 500
rect 255 -488 271 488
rect 305 -488 321 488
rect 255 -500 321 -488
rect 351 488 417 500
rect 351 -488 367 488
rect 401 -488 417 488
rect 351 -500 417 -488
rect 447 488 513 500
rect 447 -488 463 488
rect 497 -488 513 488
rect 447 -500 513 -488
rect 543 488 609 500
rect 543 -488 559 488
rect 593 -488 609 488
rect 543 -500 609 -488
rect 639 488 705 500
rect 639 -488 655 488
rect 689 -488 705 488
rect 639 -500 705 -488
rect 735 488 801 500
rect 735 -488 751 488
rect 785 -488 801 488
rect 735 -500 801 -488
rect 831 488 897 500
rect 831 -488 847 488
rect 881 -488 897 488
rect 831 -500 897 -488
rect 927 488 989 500
rect 927 -488 943 488
rect 977 -488 989 488
rect 927 -500 989 -488
<< ndiffc >>
rect -977 -488 -943 488
rect -881 -488 -847 488
rect -785 -488 -751 488
rect -689 -488 -655 488
rect -593 -488 -559 488
rect -497 -488 -463 488
rect -401 -488 -367 488
rect -305 -488 -271 488
rect -209 -488 -175 488
rect -113 -488 -79 488
rect -17 -488 17 488
rect 79 -488 113 488
rect 175 -488 209 488
rect 271 -488 305 488
rect 367 -488 401 488
rect 463 -488 497 488
rect 559 -488 593 488
rect 655 -488 689 488
rect 751 -488 785 488
rect 847 -488 881 488
rect 943 -488 977 488
<< poly >>
rect -849 662 -783 678
rect -849 628 -833 662
rect -799 628 -783 662
rect -849 612 -783 628
rect -831 550 -801 612
rect -927 520 927 550
rect -927 500 -897 520
rect -831 500 -801 520
rect -735 500 -705 520
rect -639 500 -609 520
rect -543 500 -513 520
rect -447 500 -417 520
rect -351 500 -321 520
rect -255 500 -225 520
rect -159 500 -129 520
rect -63 500 -33 520
rect 33 500 63 520
rect 129 500 159 520
rect 225 500 255 520
rect 321 500 351 520
rect 417 500 447 520
rect 513 500 543 520
rect 609 500 639 520
rect 705 500 735 520
rect 801 500 831 520
rect 897 500 927 520
rect -927 -526 -897 -500
rect -831 -526 -801 -500
rect -735 -526 -705 -500
rect -639 -526 -609 -500
rect -543 -526 -513 -500
rect -447 -526 -417 -500
rect -351 -526 -321 -500
rect -255 -526 -225 -500
rect -159 -526 -129 -500
rect -63 -526 -33 -500
rect 33 -526 63 -500
rect 129 -526 159 -500
rect 225 -526 255 -500
rect 321 -526 351 -500
rect 417 -526 447 -500
rect 513 -526 543 -500
rect 609 -526 639 -500
rect 705 -526 735 -500
rect 801 -526 831 -500
rect 897 -526 927 -500
<< polycont >>
rect -833 628 -799 662
<< locali >>
rect -849 628 -833 662
rect -799 628 -783 662
rect -881 542 883 576
rect -977 488 -943 504
rect -977 -546 -943 -488
rect -881 488 -847 542
rect -881 -504 -847 -488
rect -785 488 -751 504
rect -785 -546 -751 -488
rect -689 488 -655 542
rect -689 -504 -655 -488
rect -593 488 -559 504
rect -593 -546 -559 -488
rect -497 488 -463 542
rect -497 -504 -463 -488
rect -401 488 -367 504
rect -401 -546 -367 -488
rect -305 488 -271 542
rect -305 -504 -271 -488
rect -209 488 -175 504
rect -209 -546 -175 -488
rect -113 488 -79 542
rect -113 -504 -79 -488
rect -17 488 17 504
rect -17 -546 17 -488
rect 79 488 113 542
rect 79 -504 113 -488
rect 175 488 209 504
rect 175 -546 209 -488
rect 271 488 305 542
rect 271 -504 305 -488
rect 367 488 401 504
rect 367 -546 401 -488
rect 463 488 497 542
rect 463 -504 497 -488
rect 559 488 593 504
rect 559 -546 593 -488
rect 655 488 689 542
rect 655 -504 689 -488
rect 751 488 785 504
rect 751 -546 785 -488
rect 847 488 881 542
rect 847 -504 881 -488
rect 943 488 977 504
rect 943 -546 977 -488
rect -977 -580 977 -546
<< viali >>
rect -833 628 -799 662
rect -977 -488 -943 488
rect -881 -488 -847 488
rect -785 -488 -751 488
rect -689 -488 -655 488
rect -593 -488 -559 488
rect -497 -488 -463 488
rect -401 -488 -367 488
rect -305 -488 -271 488
rect -209 -488 -175 488
rect -113 -488 -79 488
rect -17 -488 17 488
rect 79 -488 113 488
rect 175 -488 209 488
rect 271 -488 305 488
rect 367 -488 401 488
rect 463 -488 497 488
rect 559 -488 593 488
rect 655 -488 689 488
rect 751 -488 785 488
rect 847 -488 881 488
rect 943 -488 977 488
<< metal1 >>
rect -845 662 -787 668
rect -845 628 -833 662
rect -799 628 -787 662
rect -845 622 -787 628
rect -983 488 -937 500
rect -983 -488 -977 488
rect -943 -488 -937 488
rect -983 -500 -937 -488
rect -887 488 -841 500
rect -887 -488 -881 488
rect -847 -488 -841 488
rect -887 -500 -841 -488
rect -791 488 -745 500
rect -791 -488 -785 488
rect -751 -488 -745 488
rect -791 -500 -745 -488
rect -695 488 -649 500
rect -695 -488 -689 488
rect -655 -488 -649 488
rect -695 -500 -649 -488
rect -599 488 -553 500
rect -599 -488 -593 488
rect -559 -488 -553 488
rect -599 -500 -553 -488
rect -503 488 -457 500
rect -503 -488 -497 488
rect -463 -488 -457 488
rect -503 -500 -457 -488
rect -407 488 -361 500
rect -407 -488 -401 488
rect -367 -488 -361 488
rect -407 -500 -361 -488
rect -311 488 -265 500
rect -311 -488 -305 488
rect -271 -488 -265 488
rect -311 -500 -265 -488
rect -215 488 -169 500
rect -215 -488 -209 488
rect -175 -488 -169 488
rect -215 -500 -169 -488
rect -119 488 -73 500
rect -119 -488 -113 488
rect -79 -488 -73 488
rect -119 -500 -73 -488
rect -23 488 23 500
rect -23 -488 -17 488
rect 17 -488 23 488
rect -23 -500 23 -488
rect 73 488 119 500
rect 73 -488 79 488
rect 113 -488 119 488
rect 73 -500 119 -488
rect 169 488 215 500
rect 169 -488 175 488
rect 209 -488 215 488
rect 169 -500 215 -488
rect 265 488 311 500
rect 265 -488 271 488
rect 305 -488 311 488
rect 265 -500 311 -488
rect 361 488 407 500
rect 361 -488 367 488
rect 401 -488 407 488
rect 361 -500 407 -488
rect 457 488 503 500
rect 457 -488 463 488
rect 497 -488 503 488
rect 457 -500 503 -488
rect 553 488 599 500
rect 553 -488 559 488
rect 593 -488 599 488
rect 553 -500 599 -488
rect 649 488 695 500
rect 649 -488 655 488
rect 689 -488 695 488
rect 649 -500 695 -488
rect 745 488 791 500
rect 745 -488 751 488
rect 785 -488 791 488
rect 745 -500 791 -488
rect 841 488 887 500
rect 841 -488 847 488
rect 881 -488 887 488
rect 841 -500 887 -488
rect 937 488 983 500
rect 937 -488 943 488
rect 977 -488 983 488
rect 937 -500 983 -488
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string parameters w 5 l 0.150 m 1 nf 20 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
