* NGSPICE file created from user_analog_project_wrapper_flat.ext - technology: sky130A

.subckt user_analog_project_wrapper_flat gpio_analog[0] gpio_analog[10] gpio_analog[11]
+ gpio_analog[12] gpio_analog[13] gpio_analog[14] gpio_analog[15] gpio_analog[16]
+ gpio_analog[17] gpio_analog[1] gpio_analog[2] gpio_analog[3] gpio_analog[4]
+ gpio_analog[5] gpio_analog[6] gpio_analog[7] gpio_analog[8] gpio_analog[9]
+ gpio_noesd[0] gpio_noesd[10] gpio_noesd[11] gpio_noesd[12] gpio_noesd[13]
+ gpio_noesd[14] gpio_noesd[15] gpio_noesd[16] gpio_noesd[17] gpio_noesd[1]
+ gpio_noesd[2] gpio_noesd[3] gpio_noesd[4] gpio_noesd[5] gpio_noesd[6]
+ gpio_noesd[7] gpio_noesd[8] gpio_noesd[9] io_analog[0] io_analog[10]
+ io_analog[1] io_analog[2] io_analog[3] io_analog[4] io_analog[5]
+ io_analog[6] io_analog[7] io_analog[8] io_analog[9] io_clamp_high[0]
+ io_clamp_high[1] io_clamp_high[2] io_clamp_low[0] io_clamp_low[1] io_clamp_low[2]
+ io_in[0] io_in[10] io_in[11] io_in[12] io_in[13]
+ io_in[14] io_in[15] io_in[16] io_in[17] io_in[18]
+ io_in[19] io_in[1] io_in[20] io_in[21] io_in[22]
+ io_in[23] io_in[24] io_in[25] io_in[26] io_in[2]
+ io_in[3] io_in[4] io_in[5] io_in[6] io_in[7]
+ io_in[8] io_in[9] io_in_3v3[0] io_in_3v3[10] io_in_3v3[11]
+ io_in_3v3[12] io_in_3v3[13] io_in_3v3[14] io_in_3v3[15] io_in_3v3[16]
+ io_in_3v3[17] io_in_3v3[18] io_in_3v3[19] io_in_3v3[1] io_in_3v3[20]
+ io_in_3v3[21] io_in_3v3[22] io_in_3v3[23] io_in_3v3[24] io_in_3v3[25]
+ io_in_3v3[26] io_in_3v3[2] io_in_3v3[3] io_in_3v3[4] io_in_3v3[5]
+ io_in_3v3[6] io_in_3v3[7] io_in_3v3[8] io_in_3v3[9] io_oeb[0]
+ io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14]
+ io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19]
+ io_oeb[1] io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23]
+ io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[2] io_oeb[3]
+ io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8]
+ io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12]
+ io_out[13] io_out[14] io_out[15] io_out[16] io_out[17]
+ io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26]
+ io_out[2] io_out[3] io_out[4] io_out[5] io_out[6]
+ io_out[7] io_out[8] io_out[9] la_data_in[0] la_data_in[100]
+ la_data_in[101] la_data_in[102] la_data_in[103] la_data_in[104] la_data_in[105]
+ la_data_in[106] la_data_in[107] la_data_in[108] la_data_in[109] la_data_in[10]
+ la_data_in[110] la_data_in[111] la_data_in[112] la_data_in[113] la_data_in[114]
+ la_data_in[115] la_data_in[116] la_data_in[117] la_data_in[118] la_data_in[119]
+ la_data_in[11] la_data_in[120] la_data_in[121] la_data_in[122] la_data_in[123]
+ la_data_in[124] la_data_in[125] la_data_in[126] la_data_in[127] la_data_in[12]
+ la_data_in[13] la_data_in[14] la_data_in[15] la_data_in[16] la_data_in[17]
+ la_data_in[18] la_data_in[19] la_data_in[1] la_data_in[20] la_data_in[21]
+ la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25] la_data_in[26]
+ la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30]
+ la_data_in[31] la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35]
+ la_data_in[36] la_data_in[37] la_data_in[38] la_data_in[39] la_data_in[3]
+ la_data_in[40] la_data_in[41] la_data_in[42] la_data_in[43] la_data_in[44]
+ la_data_in[45] la_data_in[46] la_data_in[47] la_data_in[48] la_data_in[49]
+ la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52] la_data_in[53]
+ la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58]
+ la_data_in[59] la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62]
+ la_data_in[63] la_data_in[64] la_data_in[65] la_data_in[66] la_data_in[67]
+ la_data_in[68] la_data_in[69] la_data_in[6] la_data_in[70] la_data_in[71]
+ la_data_in[72] la_data_in[73] la_data_in[74] la_data_in[75] la_data_in[76]
+ la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7] la_data_in[80]
+ la_data_in[81] la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85]
+ la_data_in[86] la_data_in[87] la_data_in[88] la_data_in[89] la_data_in[8]
+ la_data_in[90] la_data_in[91] la_data_in[92] la_data_in[93] la_data_in[94]
+ la_data_in[95] la_data_in[96] la_data_in[97] la_data_in[98] la_data_in[99]
+ la_data_in[9] la_data_out[0] la_data_out[100] la_data_out[101] la_data_out[102]
+ la_data_out[103] la_data_out[104] la_data_out[105] la_data_out[106] la_data_out[107]
+ la_data_out[108] la_data_out[109] la_data_out[10] la_data_out[110] la_data_out[111]
+ la_data_out[112] la_data_out[113] la_data_out[114] la_data_out[115] la_data_out[116]
+ la_data_out[117] la_data_out[118] la_data_out[119] la_data_out[11] la_data_out[120]
+ la_data_out[121] la_data_out[122] la_data_out[123] la_data_out[124] la_data_out[125]
+ la_data_out[126] la_data_out[127] la_data_out[12] la_data_out[13] la_data_out[14]
+ la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19]
+ la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23]
+ la_data_out[24] la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28]
+ la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32]
+ la_data_out[33] la_data_out[34] la_data_out[35] la_data_out[36] la_data_out[37]
+ la_data_out[38] la_data_out[39] la_data_out[3] la_data_out[40] la_data_out[41]
+ la_data_out[42] la_data_out[43] la_data_out[44] la_data_out[45] la_data_out[46]
+ la_data_out[47] la_data_out[48] la_data_out[49] la_data_out[4] la_data_out[50]
+ la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54] la_data_out[55]
+ la_data_out[56] la_data_out[57] la_data_out[58] la_data_out[59] la_data_out[5]
+ la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[64]
+ la_data_out[65] la_data_out[66] la_data_out[67] la_data_out[68] la_data_out[69]
+ la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72] la_data_out[73]
+ la_data_out[74] la_data_out[75] la_data_out[76] la_data_out[77] la_data_out[78]
+ la_data_out[79] la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82]
+ la_data_out[83] la_data_out[84] la_data_out[85] la_data_out[86] la_data_out[87]
+ la_data_out[88] la_data_out[89] la_data_out[8] la_data_out[90] la_data_out[91]
+ la_data_out[92] la_data_out[93] la_data_out[94] la_data_out[95] la_data_out[96]
+ la_data_out[97] la_data_out[98] la_data_out[99] la_data_out[9] la_oenb[0]
+ la_oenb[100] la_oenb[101] la_oenb[102] la_oenb[103] la_oenb[104]
+ la_oenb[105] la_oenb[106] la_oenb[107] la_oenb[108] la_oenb[109]
+ la_oenb[10] la_oenb[110] la_oenb[111] la_oenb[112] la_oenb[113]
+ la_oenb[114] la_oenb[115] la_oenb[116] la_oenb[117] la_oenb[118]
+ la_oenb[119] la_oenb[11] la_oenb[120] la_oenb[121] la_oenb[122]
+ la_oenb[123] la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127]
+ la_oenb[12] la_oenb[13] la_oenb[14] la_oenb[15] la_oenb[16]
+ la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20]
+ la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25]
+ la_oenb[26] la_oenb[27] la_oenb[28] la_oenb[29] la_oenb[2]
+ la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33] la_oenb[34]
+ la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38] la_oenb[39]
+ la_oenb[3] la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43]
+ la_oenb[44] la_oenb[45] la_oenb[46] la_oenb[47] la_oenb[48]
+ la_oenb[49] la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52]
+ la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57]
+ la_oenb[58] la_oenb[59] la_oenb[5] la_oenb[60] la_oenb[61]
+ la_oenb[62] la_oenb[63] la_oenb[64] la_oenb[65] la_oenb[66]
+ la_oenb[67] la_oenb[68] la_oenb[69] la_oenb[6] la_oenb[70]
+ la_oenb[71] la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75]
+ la_oenb[76] la_oenb[77] la_oenb[78] la_oenb[79] la_oenb[7]
+ la_oenb[80] la_oenb[81] la_oenb[82] la_oenb[83] la_oenb[84]
+ la_oenb[85] la_oenb[86] la_oenb[87] la_oenb[88] la_oenb[89]
+ la_oenb[8] la_oenb[90] la_oenb[91] la_oenb[92] la_oenb[93]
+ la_oenb[94] la_oenb[95] la_oenb[96] la_oenb[97] la_oenb[98]
+ la_oenb[99] la_oenb[9] user_clock2 user_irq[0] user_irq[1]
+ user_irq[2] vccd2 vdda1 vdda2 vssa2
+ vssd1 vssd2 wb_clk_i wb_rst_i wbs_ack_o
+ wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13]
+ wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18]
+ wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22]
+ wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27]
+ wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31]
+ wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7]
+ wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10]
+ wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15]
+ wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1]
+ wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24]
+ wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29]
+ wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4]
+ wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9]
+ wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13]
+ wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18]
+ wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22]
+ wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27]
+ wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31]
+ wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7]
+ wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2]
+ wbs_sel_i[3] wbs_stb_i wbs_we_i vssa1 vccd1
X0 esd_3/in vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1 vssa1 vssa1 esd_4/in vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X2 a_481708_644918# a_483446_644892# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3 vssa1 VCO_Flat_0/Buff_VCO_1/IN a_504724_647182# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4 vssa1 vssa1 io_analog[5] vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X5 vccd1 a_471230_648050# esd_5/in vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6 esd_0/in a_500126_647170# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7 vssa1 vssa1 esd_4/in vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X8 vssa1 vssa1 esd_1/in vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X9 vccd1 a_475058_648060# a_473374_648060# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10 a_487694_644902# VCO_Flat_0/Buff_VCO_3/IN VCO_Flat_0/Buff_VCO_2/IN vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X11 io_analog[5] vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X12 vssa1 a_479772_646886# a_493938_644874# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X13 io_analog[4] vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X14 vccd1 a_498236_647184# a_498928_647174# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X15 esd_5/in a_471230_648050# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X16 vssa1 a_468592_648062# a_466908_648062# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X17 vssa1 vssa1 io_analog[7] vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X18 esd_4/in vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X19 esd_1/in vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X20 vccd1 esd_1/in a_493974_650212# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X21 esd_0/in a_500126_647170# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X22 esd_6/in a_506614_647168# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X23 vssa1 a_479772_646886# a_479772_646886# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=200000u
X24 esd_5/in a_471230_648050# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X25 io_analog[4] vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X26 vssa1 vssa1 io_analog[4] vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X27 a_464764_648054# a_466908_648062# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X28 a_500126_647170# a_498928_647174# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X29 a_479772_646886# esd_2/in a_479864_646886# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X30 esd_6/in vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X31 vccd1 vccd1 io_analog[6] vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X32 io_analog[4] vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X33 a_498236_647184# VCO_Flat_0/Buff_VCO_0/IN vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X34 esd_5/in vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X35 vccd1 a_471230_648050# esd_5/in vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X36 a_506614_647168# a_505416_647172# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X37 esd_0/in a_500126_647170# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X38 vssa1 a_498928_647174# a_500126_647170# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X39 vccd1 vccd1 esd_6/in vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X40 io_analog[7] vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X41 vssa1 vssa1 esd_6/in vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X42 a_487730_650240# esd_1/in vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X43 vccd1 a_475058_648060# a_473374_648060# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X44 io_analog[6] vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X45 vssa1 vssa1 esd_3/in vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X46 a_506614_647168# a_505416_647172# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X47 vssa1 vssa1 esd_5/in vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X48 vccd1 a_498236_647184# a_498928_647174# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X49 esd_6/in a_506614_647168# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X50 vssa1 a_498928_647174# a_500126_647170# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X51 a_479772_646886# a_479772_646886# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=200000u
X52 vssa1 VCO_Flat_0/Buff_VCO_3/IN a_468592_648062# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X53 io_analog[5] vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X54 a_464764_648054# a_466908_648062# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X55 a_500126_647170# a_498928_647174# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X56 esd_0/in a_500126_647170# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X57 vccd1 a_479864_646886# a_481744_650256# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X58 esd_3/in a_457934_648038# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X59 vssa1 a_479772_646886# a_490782_644900# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X60 esd_6/in a_506614_647168# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X61 esd_4/in vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X62 vssa1 vssa1 io_analog[6] vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X63 vccd1 a_479864_646886# a_484700_650240# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X64 vccd1 a_473374_648060# a_471230_648050# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X65 a_504724_647182# VCO_Flat_0/Buff_VCO_1/IN vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X66 io_analog[5] vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X67 vccd1 vccd1 io_analog[5] vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X68 io_analog[7] vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X69 esd_4/in vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X70 vccd1 a_504724_647182# a_505416_647172# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X71 esd_0/in a_500126_647170# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X72 vssa1 a_466908_648062# a_464764_648054# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X73 vccd1 vccd1 esd_4/in vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X74 io_analog[6] vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X75 a_475058_648060# VCO_Flat_0/Buff_VCO_2/IN vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X76 vccd1 vccd1 io_analog[4] vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X77 vccd1 a_479864_646886# a_484700_650240# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X78 vccd1 esd_1/in a_490818_650238# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X79 vccd1 a_473374_648060# a_471230_648050# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X80 vccd1 vccd1 esd_4/in vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X81 vccd1 a_479864_646886# a_481744_650256# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X82 VCO_Flat_0/Buff_VCO_0/IN VCO_Flat_0/Buff_VCO_3/IN a_493974_650212# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X83 vccd1 vccd1 esd_0/in vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X84 VCO_Flat_0/Buff_VCO_3/IN VCO_Flat_0/Buff_VCO_1/IN a_484700_650240# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X85 vssa1 a_466908_648062# a_464764_648054# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X86 a_504724_647182# VCO_Flat_0/Buff_VCO_1/IN vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X87 vccd1 vccd1 esd_4/in vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X88 esd_0/in vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X89 vccd1 a_500126_647170# esd_0/in vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X90 vccd1 esd_1/in a_490818_650238# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X91 vssa1 a_483446_644892# a_487694_644902# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X92 VCO_Flat_0/Buff_VCO_3/IN VCO_Flat_0/Buff_VCO_4/IN a_484664_644902# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X93 a_493938_644874# a_479772_646886# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X94 esd_5/in vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X95 VCO_Flat_0/Buff_VCO_3/IN VCO_Flat_0/Buff_VCO_1/IN a_484700_650240# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X96 vccd1 vccd1 esd_5/in vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X97 vssa1 vssa1 esd_0/in vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X98 io_analog[2] vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X99 vccd1 a_506614_647168# esd_6/in vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X100 esd_5/in vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X101 vccd1 a_479864_646886# a_493974_650212# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X102 a_479864_646886# esd_2/in a_479772_646886# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X103 io_analog[2] vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X104 vccd1 a_457934_648038# esd_3/in vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X105 vccd1 a_461762_648050# a_460078_648050# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X106 vccd1 a_500126_647170# esd_0/in vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X107 vssa1 vssa1 esd_0/in vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X108 vccd1 a_506614_647168# esd_6/in vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X109 vssa1 a_479772_646886# a_484664_644902# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X110 a_490782_644900# a_483446_644892# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X111 VCO_Flat_0/Buff_VCO_2/IN VCO_Flat_0/Buff_VCO_3/IN a_487694_644902# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X112 esd_5/in vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X113 esd_5/in a_471230_648050# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X114 esd_5/in a_471230_648050# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X115 vccd1 vccd1 esd_3/in vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X116 io_analog[2] vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X117 vccd1 a_500126_647170# esd_0/in vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X118 io_analog[2] vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X119 a_473374_648060# a_475058_648060# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X120 esd_3/in vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X121 vccd1 vccd1 io_analog[1] vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X122 vccd1 esd_1/in a_484700_650240# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X123 a_490818_650238# VCO_Flat_0/Buff_VCO_4/IN VCO_Flat_0/Buff_VCO_1/IN vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X124 vccd1 a_505416_647172# a_506614_647168# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X125 esd_4/in io_analog[4] vssa1 sky130_fd_pr__res_high_po w=2.85e+06u l=1.3e+06u
X126 a_481744_650256# VCO_Flat_0/Buff_VCO_2/IN VCO_Flat_0/Buff_VCO_4/IN vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X127 a_498928_647174# a_498236_647184# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X128 a_500126_647170# a_498928_647174# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X129 vssa1 a_471230_648050# esd_5/in vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X130 esd_4/in a_464764_648054# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X131 vccd1 vccd1 io_analog[3] vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X132 vssa1 vssa1 esd_1/in vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X133 vccd1 a_466908_648062# a_464764_648054# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X134 vccd1 a_498928_647174# a_500126_647170# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X135 vssa1 a_457934_648038# esd_3/in vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X136 vssa1 a_506614_647168# esd_6/in vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X137 a_490782_644900# VCO_Flat_0/Buff_VCO_2/IN VCO_Flat_0/Buff_VCO_1/IN vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X138 esd_4/in a_464764_648054# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X139 io_analog[1] vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X140 a_498236_647184# VCO_Flat_0/Buff_VCO_0/IN vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X141 a_481708_644918# VCO_Flat_0/Buff_VCO_0/IN VCO_Flat_0/Buff_VCO_4/IN vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X142 a_473374_648060# a_475058_648060# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X143 vccd1 VCO_Flat_0/Buff_VCO_2/IN a_475058_648060# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X144 vccd1 a_498928_647174# a_500126_647170# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X145 vssa1 a_500126_647170# esd_0/in vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X146 a_464764_648054# a_466908_648062# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X147 vssa1 vssa1 io_analog[3] vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X148 vssa1 vssa1 io_analog[1] vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X149 a_484700_650240# a_479864_646886# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X150 a_471230_648050# a_473374_648060# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X151 a_490818_650238# a_479864_646886# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X152 vccd1 vccd1 io_analog[7] vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X153 esd_1/in vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X154 esd_3/in vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X155 a_481744_650256# a_479864_646886# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X156 vccd1 a_505416_647172# a_506614_647168# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X157 vssa1 a_457934_648038# esd_3/in vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X158 a_484700_650240# VCO_Flat_0/Buff_VCO_1/IN VCO_Flat_0/Buff_VCO_3/IN vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X159 a_498928_647174# a_498236_647184# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X160 a_464764_648054# a_466908_648062# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X161 vssa1 vssa1 io_analog[3] vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X162 vssa1 vssa1 io_analog[5] vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X163 vssa1 a_457934_648038# esd_3/in vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X164 vccd1 vccd1 io_analog[7] vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X165 io_analog[3] vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X166 a_490818_650238# a_479864_646886# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X167 a_490818_650238# esd_1/in vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X168 a_487694_644902# a_483446_644892# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X169 a_506614_647168# a_505416_647172# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X170 a_484664_644902# VCO_Flat_0/Buff_VCO_4/IN VCO_Flat_0/Buff_VCO_3/IN vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X171 a_481744_650256# esd_1/in vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X172 a_481708_644918# a_479772_646886# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X173 vssa1 vssa1 esd_1/in vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X174 esd_6/in a_506614_647168# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X175 vccd1 vccd1 esd_3/in vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X176 io_analog[7] vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X177 a_460078_648050# a_461762_648050# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X178 esd_0/in a_500126_647170# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X179 io_analog[4] vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X180 vccd1 esd_1/in a_487730_650240# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X181 esd_6/in a_506614_647168# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X182 a_484664_644902# a_479772_646886# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X183 vccd1 vccd1 io_analog[4] vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X184 vccd1 a_471230_648050# esd_5/in vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X185 a_481708_644918# a_479772_646886# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X186 vssa1 vssa1 esd_4/in vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X187 vssa1 vssa1 esd_1/in vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X188 esd_0/in a_500126_647170# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X189 io_analog[6] vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X190 a_484700_650240# esd_1/in vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X191 a_460078_648050# a_461762_648050# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X192 a_506614_647168# a_505416_647172# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X193 esd_3/in vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X194 VCO_Flat_0/Buff_VCO_4/IN VCO_Flat_0/Buff_VCO_2/IN a_481744_650256# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X195 a_505416_647172# a_504724_647182# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X196 esd_5/in a_471230_648050# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X197 vssa1 a_464764_648054# esd_4/in vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X198 esd_6/in vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X199 vssa1 vssa1 esd_3/in vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X200 a_493974_650212# a_479864_646886# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X201 esd_6/in vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X202 a_500126_647170# a_498928_647174# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X203 a_466908_648062# a_468592_648062# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X204 a_506614_647168# a_505416_647172# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X205 VCO_Flat_0/Buff_VCO_1/IN VCO_Flat_0/Buff_VCO_2/IN a_490782_644900# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X206 esd_6/in vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X207 io_analog[6] vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X208 esd_2/in io_analog[2] vssa1 sky130_fd_pr__res_high_po w=2.85e+06u l=1.3e+06u
X209 VCO_Flat_0/Buff_VCO_4/IN VCO_Flat_0/Buff_VCO_0/IN a_481708_644918# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X210 vssa1 vssa1 esd_6/in vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X211 esd_4/in a_464764_648054# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X212 vccd1 a_471230_648050# esd_5/in vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X213 a_500126_647170# a_498928_647174# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X214 vssa1 vssa1 io_analog[6] vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X215 vssa1 a_464764_648054# esd_4/in vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X216 io_analog[5] vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X217 esd_5/in vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X218 a_466908_648062# a_468592_648062# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X219 vccd1 vccd1 io_analog[7] vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X220 esd_4/in vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X221 vccd1 a_479864_646886# a_490818_650238# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X222 vccd1 a_457934_648038# esd_3/in vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X223 vssa1 vssa1 esd_6/in vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X224 vssa1 vssa1 io_analog[6] vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X225 a_506614_647168# a_505416_647172# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X226 esd_3/in a_457934_648038# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X227 a_493938_644874# a_483446_644892# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X228 vssa1 a_498236_647184# a_498928_647174# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X229 vssa1 a_466908_648062# a_464764_648054# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X230 vssa1 a_464764_648054# esd_4/in vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X231 vccd1 VCO_Flat_0/Buff_VCO_4/IN a_461762_648050# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X232 vssa1 a_460078_648050# a_457934_648038# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X233 vssa1 vssa1 io_analog[6] vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X234 esd_3/in a_457934_648038# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X235 vccd1 a_479864_646886# a_490818_650238# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X236 vssa1 a_505416_647172# a_506614_647168# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X237 esd_3/in io_analog[3] vssa1 sky130_fd_pr__res_high_po w=2.85e+06u l=1.3e+06u
X238 vccd1 esd_1/in a_481744_650256# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X239 vssa1 a_475058_648060# a_473374_648060# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X240 esd_0/in a_500126_647170# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X241 vssa1 a_498236_647184# a_498928_647174# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X242 vssa1 a_466908_648062# a_464764_648054# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X243 vssa1 vssa1 esd_2/in vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X244 vccd1 VCO_Flat_0/Buff_VCO_4/IN a_461762_648050# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X245 vccd1 a_473374_648060# a_471230_648050# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X246 vccd1 vccd1 esd_0/in vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X247 vssa1 vssa1 io_analog[2] vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X248 vccd1 a_479864_646886# a_490818_650238# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X249 vccd1 vccd1 esd_2/in vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X250 vssa1 a_479772_646886# a_484664_644902# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X251 esd_6/in a_506614_647168# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X252 vccd1 vccd1 esd_0/in vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X253 vccd1 vccd1 io_analog[2] vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X254 vssa1 a_498236_647184# a_498928_647174# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X255 VCO_Flat_0/Buff_VCO_3/IN VCO_Flat_0/Buff_VCO_1/IN vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X256 esd_0/in vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X257 vssa1 a_479772_646886# a_481708_644918# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X258 vssa1 a_505416_647172# a_506614_647168# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X259 io_analog[4] vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X260 vssa1 vssa1 esd_2/in vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X261 esd_0/in vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X262 vccd1 vccd1 esd_2/in vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X263 io_analog[2] vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X264 vssa1 a_505416_647172# a_506614_647168# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X265 esd_0/in vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X266 vccd1 a_461762_648050# a_460078_648050# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X267 vssa1 a_479772_646886# a_481708_644918# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X268 vccd1 vccd1 esd_5/in vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X269 io_analog[2] vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X270 io_analog[1] vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X271 vssa1 a_504724_647182# a_505416_647172# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X272 vccd1 vccd1 io_analog[1] vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X273 vccd1 a_479864_646886# a_493974_650212# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X274 esd_0/in vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X275 vssa1 vssa1 esd_0/in vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X276 vccd1 esd_1/in a_484700_650240# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X277 vccd1 a_461762_648050# a_460078_648050# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X278 a_490782_644900# a_483446_644892# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X279 vccd1 vccd1 esd_3/in vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X280 vccd1 vccd1 io_analog[1] vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X281 vccd1 a_464764_648054# esd_4/in vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X282 a_481708_644918# VCO_Flat_0/Buff_VCO_0/IN VCO_Flat_0/Buff_VCO_4/IN vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X283 vssa1 a_471230_648050# esd_5/in vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X284 vssa1 vssa1 io_analog[1] vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X285 esd_5/in a_471230_648050# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X286 io_analog[3] vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X287 io_analog[1] vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X288 vccd1 a_500126_647170# esd_0/in vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X289 esd_4/in a_464764_648054# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X290 vccd1 a_468592_648062# a_466908_648062# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X291 io_analog[4] vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X292 vccd1 esd_1/in a_484700_650240# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X293 vccd1 a_464764_648054# esd_4/in vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X294 vccd1 vccd1 io_analog[3] vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X295 vccd1 a_505416_647172# a_506614_647168# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X296 esd_4/in a_464764_648054# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X297 esd_0/in io_analog[6] vssa1 sky130_fd_pr__res_high_po w=2.85e+06u l=1.3e+06u
X298 vccd1 a_479864_646886# a_479864_646886# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=200000u
X299 vssa1 a_471230_648050# esd_5/in vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X300 io_analog[3] vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X301 io_analog[4] vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X302 esd_3/in vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X303 io_analog[1] vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X304 a_461762_648050# VCO_Flat_0/Buff_VCO_4/IN vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X305 a_457934_648038# a_460078_648050# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X306 vssa1 a_457934_648038# esd_3/in vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X307 esd_3/in vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X308 esd_2/in vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X309 a_490818_650238# a_479864_646886# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X310 vccd1 a_464764_648054# esd_4/in vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X311 vssa1 a_483446_644892# a_493938_644874# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X312 vssa1 a_500126_647170# esd_0/in vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X313 a_473374_648060# a_475058_648060# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X314 a_457934_648038# a_460078_648050# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X315 esd_2/in vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X316 esd_1/in vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X317 vssa1 vssa1 io_analog[3] vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X318 a_498928_647174# a_498236_647184# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X319 vssa1 vssa1 esd_2/in vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X320 a_481744_650256# a_479864_646886# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X321 a_490818_650238# a_479864_646886# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X322 esd_3/in a_457934_648038# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X323 vccd1 vccd1 esd_2/in vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X324 io_analog[5] vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X325 vssa1 a_483446_644892# a_493938_644874# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X326 vssa1 a_506614_647168# esd_6/in vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X327 esd_1/in vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X328 a_506614_647168# a_505416_647172# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X329 a_498928_647174# a_498236_647184# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X330 esd_4/in vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X331 vssa1 vssa1 esd_1/in vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X332 a_479864_646886# a_479864_646886# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=200000u
X333 a_487694_644902# a_479772_646886# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X334 a_481708_644918# a_479772_646886# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X335 io_analog[5] vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X336 vssa1 vssa1 io_analog[5] vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X337 vccd1 vccd1 io_analog[4] vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X338 vssa1 vssa1 io_analog[7] vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X339 esd_4/in vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X340 vssa1 vssa1 esd_4/in vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X341 a_481708_644918# a_479772_646886# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X342 a_506614_647168# a_505416_647172# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X343 vssa1 vssa1 io_analog[4] vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X344 vssa1 vssa1 esd_1/in vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X345 a_505416_647172# a_504724_647182# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X346 vccd1 vccd1 esd_6/in vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X347 vssa1 vssa1 esd_4/in vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X348 esd_1/in vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X349 a_493974_650212# a_479864_646886# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X350 esd_3/in vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
R0 vccd1 io_clamp_high[1] sky130_fd_pr__res_generic_m3 w=1.08e+07u l=1.29e+06u
X351 vccd1 vccd1 io_analog[4] vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X352 vssa1 vssa1 esd_4/in vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X353 vssa1 a_483446_644892# a_490782_644900# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X354 vssa1 a_483446_644892# a_490782_644900# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X355 a_475058_648060# VCO_Flat_0/Buff_VCO_2/IN vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X356 esd_6/in vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X357 esd_4/in a_464764_648054# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X358 vccd1 a_471230_648050# esd_5/in vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X359 vccd1 vccd1 esd_6/in vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X360 io_analog[6] vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X361 esd_0/in a_500126_647170# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X362 esd_1/in io_analog[1] vssa1 sky130_fd_pr__res_high_po w=2.85e+06u l=1.3e+06u
X363 esd_5/in vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X364 a_466908_648062# a_468592_648062# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X365 esd_6/in vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X366 vssa1 vssa1 esd_5/in vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X367 esd_5/in vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X368 a_504724_647182# VCO_Flat_0/Buff_VCO_1/IN vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X369 vccd1 vccd1 io_analog[7] vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X370 esd_6/in a_506614_647168# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X371 esd_6/in vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X372 vssa1 vssa1 io_analog[6] vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X373 a_493974_650212# a_479864_646886# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X374 esd_4/in a_464764_648054# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X375 vssa1 a_460078_648050# a_457934_648038# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X376 esd_5/in vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X377 a_466908_648062# a_468592_648062# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X378 vssa1 vssa1 esd_6/in vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X379 esd_4/in a_464764_648054# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X380 io_analog[7] vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X381 vccd1 a_479864_646886# a_487730_650240# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X382 a_487694_644902# a_483446_644892# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X383 a_493938_644874# a_483446_644892# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X384 vssa1 a_475058_648060# a_473374_648060# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X385 vssa1 a_460078_648050# a_457934_648038# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X386 io_analog[6] vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X387 a_504724_647182# VCO_Flat_0/Buff_VCO_1/IN vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X388 io_analog[5] vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X389 vccd1 a_457934_648038# esd_3/in vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X390 a_493938_644874# a_479772_646886# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X391 vccd1 a_479864_646886# a_481744_650256# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X392 a_493938_644874# VCO_Flat_0/Buff_VCO_1/IN VCO_Flat_0/Buff_VCO_0/IN vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X393 vccd1 vccd1 esd_4/in vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X394 esd_4/in vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X395 a_493938_644874# a_483446_644892# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X396 esd_6/in a_506614_647168# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X397 vssa1 a_464764_648054# esd_4/in vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X398 vccd1 vccd1 esd_0/in vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X399 io_analog[4] vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X400 vssa1 a_483446_644892# a_484664_644902# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X401 a_460078_648050# a_461762_648050# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X402 a_479864_646886# a_479864_646886# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=200000u
X403 vssa1 a_460078_648050# a_457934_648038# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X404 vssa1 a_479772_646886# a_487694_644902# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X405 esd_0/in vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X406 io_analog[2] vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X407 vccd1 a_479864_646886# a_479864_646886# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=200000u
X408 vccd1 vccd1 io_analog[4] vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X409 io_analog[2] vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X410 vssa1 a_505416_647172# a_506614_647168# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X411 vccd1 vccd1 esd_0/in vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X412 esd_5/in vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X413 vssa1 vssa1 io_analog[2] vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X414 vccd1 vccd1 io_analog[2] vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X415 vssa1 vssa1 esd_0/in vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X416 vssa1 a_479772_646886# a_487694_644902# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X417 vccd1 vccd1 esd_5/in vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X418 a_493974_650212# esd_1/in vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X419 io_analog[1] vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X420 vssa1 vssa1 io_analog[2] vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X421 a_490782_644900# a_483446_644892# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X422 vssa1 VCO_Flat_0/Buff_VCO_2/IN a_475058_648060# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X423 esd_5/in vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X424 esd_0/in vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X425 vccd1 a_466908_648062# a_464764_648054# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X426 vccd1 vccd1 io_analog[2] vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X427 vccd1 VCO_Flat_0/Buff_VCO_3/IN a_468592_648062# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X428 vssa1 a_479772_646886# a_487694_644902# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X429 vssa1 a_473374_648060# a_471230_648050# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X430 io_analog[2] vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X431 vccd1 a_500126_647170# esd_0/in vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X432 vssa1 VCO_Flat_0/Buff_VCO_0/IN a_498236_647184# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X433 vccd1 vccd1 esd_5/in vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X434 vccd1 vccd1 io_analog[3] vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X435 vccd1 vccd1 esd_3/in vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X436 io_analog[5] vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X437 io_analog[2] vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X438 vssa1 a_473374_648060# a_471230_648050# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X439 vccd1 VCO_Flat_0/Buff_VCO_1/IN a_504724_647182# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X440 vccd1 a_506614_647168# esd_6/in vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X441 vccd1 a_479864_646886# a_493974_650212# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X442 vccd1 vccd1 esd_3/in vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X443 io_analog[3] vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X444 vssa1 vssa1 io_analog[4] vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X445 vssa1 vssa1 esd_3/in vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X446 vccd1 a_464764_648054# esd_4/in vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X447 esd_5/in a_471230_648050# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X448 a_487730_650240# a_479864_646886# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X449 vccd1 VCO_Flat_0/Buff_VCO_1/IN a_504724_647182# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X450 vssa1 a_483446_644892# a_487694_644902# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X451 io_analog[7] vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X452 esd_3/in vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X453 esd_2/in vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X454 vssa1 vssa1 io_analog[1] vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X455 esd_3/in a_457934_648038# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X456 vssa1 a_479772_646886# a_493938_644874# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X457 VCO_Flat_0/Buff_VCO_0/IN VCO_Flat_0/Buff_VCO_1/IN a_493938_644874# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X458 esd_2/in vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X459 vssa1 vssa1 io_analog[3] vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X460 esd_2/in vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X461 vssa1 a_483446_644892# a_493938_644874# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X462 esd_4/in a_464764_648054# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X463 vssa1 a_461762_648050# a_460078_648050# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X464 esd_6/in io_analog[7] vssa1 sky130_fd_pr__res_high_po w=2.85e+06u l=1.3e+06u
X465 a_484664_644902# a_483446_644892# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X466 io_analog[7] vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X467 esd_2/in vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X468 a_487730_650240# a_479864_646886# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X469 a_457934_648038# a_460078_648050# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X470 a_487694_644902# a_479772_646886# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X471 vccd1 vccd1 esd_1/in vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X472 a_484664_644902# a_483446_644892# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X473 io_analog[5] vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X474 a_473374_648060# a_475058_648060# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X475 esd_1/in vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X476 a_487730_650240# a_479864_646886# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X477 vssa1 vssa1 io_analog[7] vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X478 esd_4/in vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X479 esd_1/in vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X480 a_487694_644902# a_479772_646886# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X481 vccd1 esd_1/in a_493974_650212# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X482 vccd1 esd_1/in a_493974_650212# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X483 vccd1 a_460078_648050# a_457934_648038# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X484 esd_3/in vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X485 a_475058_648060# VCO_Flat_0/Buff_VCO_2/IN vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X486 a_464764_648054# a_466908_648062# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X487 vssa1 a_468592_648062# a_466908_648062# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X488 vssa1 vssa1 io_analog[7] vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X489 vccd1 a_460078_648050# a_457934_648038# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X490 a_468592_648062# VCO_Flat_0/Buff_VCO_3/IN vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X491 a_487694_644902# a_479772_646886# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X492 vccd1 vccd1 esd_6/in vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X493 a_498236_647184# VCO_Flat_0/Buff_VCO_0/IN vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X494 vccd1 a_479864_646886# a_479864_646886# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=200000u
X495 vccd1 vccd1 esd_6/in vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X496 io_analog[4] vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X497 vssa1 vssa1 esd_3/in vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X498 a_506614_647168# a_505416_647172# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X499 a_471230_648050# a_473374_648060# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X500 vssa1 VCO_Flat_0/Buff_VCO_4/IN a_461762_648050# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X501 vccd1 vccd1 esd_6/in vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X502 vccd1 vccd1 io_analog[6] vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X503 esd_3/in a_457934_648038# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X504 vssa1 a_479772_646886# a_490782_644900# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X505 io_analog[4] vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X506 io_analog[6] vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X507 vccd1 vccd1 io_analog[5] vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X508 a_471230_648050# a_473374_648060# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X509 io_analog[7] vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X510 io_analog[6] vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X511 vssa1 vssa1 esd_5/in vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X512 a_493938_644874# VCO_Flat_0/Buff_VCO_1/IN VCO_Flat_0/Buff_VCO_0/IN vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X513 esd_6/in vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X514 a_471230_648050# a_473374_648060# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X515 vccd1 vccd1 io_analog[5] vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X516 esd_4/in vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X517 esd_6/in vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X518 vssa1 a_464764_648054# esd_4/in vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X519 a_460078_648050# a_461762_648050# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X520 vssa1 a_483446_644892# a_484664_644902# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X521 vccd1 vccd1 esd_4/in vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X522 esd_6/in vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X523 io_analog[6] vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X524 vccd1 a_479864_646886# a_487730_650240# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X525 VCO_Flat_0/Buff_VCO_2/IN VCO_Flat_0/Buff_VCO_0/IN vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X526 vssa1 a_483446_644892# a_484664_644902# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X527 esd_0/in vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X528 vccd1 a_479864_646886# a_487730_650240# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X529 esd_4/in a_464764_648054# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X530 vssa1 vssa1 io_analog[7] vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X531 vssa1 a_483446_644892# a_481708_644918# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
R1 vssa1 io_clamp_low[1] sky130_fd_pr__res_generic_m3 w=1.084e+07u l=1.29e+06u
X532 vccd1 a_457934_648038# esd_3/in vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X533 VCO_Flat_0/Buff_VCO_2/IN VCO_Flat_0/Buff_VCO_0/IN a_487730_650240# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X534 vssa1 a_479772_646886# a_484664_644902# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X535 a_493974_650212# esd_1/in vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X536 a_457934_648038# a_460078_648050# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X537 vssa1 a_483446_644892# a_481708_644918# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X538 esd_5/in a_471230_648050# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X539 esd_0/in vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X540 esd_2/in vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X541 vssa1 a_479772_646886# a_487694_644902# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X542 a_466908_648062# a_468592_648062# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X543 io_analog[2] vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X544 a_457934_648038# a_460078_648050# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X545 a_473374_648060# a_475058_648060# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X546 VCO_Flat_0/Buff_VCO_2/IN VCO_Flat_0/Buff_VCO_3/IN a_487694_644902# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X547 esd_2/in vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X548 esd_5/in vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X549 io_analog[2] vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X550 vccd1 a_457934_648038# esd_3/in vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X551 VCO_Flat_0/Buff_VCO_2/IN VCO_Flat_0/Buff_VCO_0/IN a_487730_650240# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X552 a_498928_647174# a_498236_647184# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X553 vssa1 vssa1 io_analog[2] vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X554 vssa1 a_473374_648060# a_471230_648050# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X555 vssa1 a_471230_648050# esd_5/in vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X556 a_466908_648062# a_468592_648062# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X557 a_461762_648050# VCO_Flat_0/Buff_VCO_4/IN vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X558 vssa1 vssa1 esd_0/in vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X559 vccd1 vccd1 io_analog[2] vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X560 vssa1 vssa1 io_analog[2] vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X561 a_490782_644900# a_479772_646886# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X562 io_analog[1] vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X563 vssa1 vssa1 esd_0/in vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X564 a_457934_648038# a_460078_648050# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X565 a_481744_650256# VCO_Flat_0/Buff_VCO_2/IN VCO_Flat_0/Buff_VCO_4/IN vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X566 vssa1 a_457934_648038# esd_3/in vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X567 vccd1 vccd1 io_analog[2] vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X568 io_analog[1] vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X569 esd_0/in vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X570 a_498928_647174# a_498236_647184# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X571 vssa1 a_500126_647170# esd_0/in vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X572 a_500126_647170# a_498928_647174# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X573 vssa1 a_473374_648060# a_471230_648050# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X574 vssa1 vssa1 io_analog[4] vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X575 vccd1 esd_1/in a_487730_650240# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X576 esd_3/in vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X577 io_analog[1] vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X578 a_490782_644900# a_479772_646886# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X579 vssa1 a_506614_647168# esd_6/in vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X580 vccd1 vccd1 io_analog[3] vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X581 vssa1 vssa1 io_analog[1] vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X582 a_479772_646886# a_479772_646886# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=200000u
X583 vssa1 a_473374_648060# a_471230_648050# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X584 vssa1 a_479772_646886# a_479772_646886# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=200000u
X585 vssa1 vssa1 io_analog[4] vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X586 a_490782_644900# a_479772_646886# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X587 vssa1 a_500126_647170# esd_0/in vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X588 io_analog[3] vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X589 vssa1 vssa1 esd_3/in vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X590 esd_2/in vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X591 vssa1 vssa1 io_analog[1] vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X592 a_484700_650240# a_479864_646886# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X593 a_471230_648050# a_473374_648060# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X594 vssa1 a_457934_648038# esd_3/in vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X595 esd_2/in vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X596 io_analog[3] vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X597 vccd1 vccd1 esd_1/in vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X598 a_487730_650240# a_479864_646886# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X599 vccd1 a_464764_648054# esd_4/in vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X600 a_505416_647172# a_504724_647182# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X601 a_481708_644918# a_483446_644892# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X602 vssa1 vssa1 io_analog[3] vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X603 a_487730_650240# VCO_Flat_0/Buff_VCO_0/IN VCO_Flat_0/Buff_VCO_2/IN vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X604 esd_3/in a_457934_648038# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X605 a_484664_644902# a_479772_646886# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X606 io_analog[3] vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X607 a_481708_644918# a_483446_644892# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X608 vssa1 VCO_Flat_0/Buff_VCO_1/IN a_504724_647182# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X609 a_484664_644902# a_483446_644892# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X610 vssa1 a_461762_648050# a_460078_648050# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X611 esd_0/in a_500126_647170# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X612 vccd1 a_460078_648050# a_457934_648038# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X613 vccd1 a_475058_648060# a_473374_648060# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X614 a_484664_644902# a_479772_646886# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X615 a_487694_644902# VCO_Flat_0/Buff_VCO_3/IN VCO_Flat_0/Buff_VCO_2/IN vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X616 vssa1 a_479772_646886# a_493938_644874# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X617 esd_1/in vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X618 esd_3/in a_457934_648038# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X619 vccd1 a_498236_647184# a_498928_647174# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X620 vssa1 a_468592_648062# a_466908_648062# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X621 esd_5/in a_471230_648050# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X622 vssa1 VCO_Flat_0/Buff_VCO_4/IN a_461762_648050# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X623 io_analog[5] vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X624 a_479772_646886# esd_2/in a_479864_646886# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X625 io_analog[4] vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X626 vssa1 vssa1 esd_4/in vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X627 esd_4/in vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X628 io_analog[4] vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X629 esd_1/in vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X630 esd_3/in a_457934_648038# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X631 vccd1 a_460078_648050# a_457934_648038# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X632 VCO_Flat_0/Buff_VCO_4/IN VCO_Flat_0/Buff_VCO_2/IN a_481744_650256# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X633 esd_3/in a_457934_648038# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X634 esd_6/in vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X635 vccd1 vccd1 io_analog[6] vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X636 vccd1 a_471230_648050# esd_5/in vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X637 vssa1 vssa1 io_analog[4] vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X638 vssa1 a_498928_647174# a_500126_647170# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X639 a_487730_650240# esd_1/in vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X640 vccd1 a_475058_648060# a_473374_648060# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X641 VCO_Flat_0/Buff_VCO_4/IN VCO_Flat_0/Buff_VCO_0/IN a_481708_644918# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X642 vccd1 vccd1 esd_6/in vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X643 esd_5/in vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X644 VCO_Flat_0/Buff_VCO_1/IN VCO_Flat_0/Buff_VCO_4/IN a_490818_650238# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X645 vssa1 a_479772_646886# a_490782_644900# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X646 vccd1 vccd1 io_analog[7] vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X647 vccd1 a_498236_647184# a_498928_647174# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X648 esd_6/in a_506614_647168# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X649 vssa1 a_498928_647174# a_500126_647170# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X650 io_analog[7] vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X651 vccd1 vccd1 io_analog[6] vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X652 vssa1 vssa1 esd_6/in vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X653 a_471230_648050# a_473374_648060# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X654 vssa1 vssa1 esd_5/in vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X655 a_464764_648054# a_466908_648062# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X656 vccd1 vccd1 io_analog[6] vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X657 vssa1 a_479772_646886# a_490782_644900# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X658 esd_0/in a_500126_647170# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X659 vccd1 vccd1 io_analog[5] vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X660 esd_6/in vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X661 esd_5/in vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X662 vccd1 a_473374_648060# a_471230_648050# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X663 esd_3/in a_457934_648038# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X664 esd_6/in a_506614_647168# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X665 vccd1 VCO_Flat_0/Buff_VCO_0/IN a_498236_647184# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X666 vssa1 vssa1 esd_6/in vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X667 io_analog[6] vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X668 esd_0/in a_500126_647170# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X669 vssa1 a_498928_647174# a_500126_647170# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X670 vssa1 a_466908_648062# a_464764_648054# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X671 vssa1 vssa1 esd_5/in vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X672 vccd1 a_504724_647182# a_505416_647172# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X673 vccd1 a_479864_646886# a_484700_650240# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X674 vccd1 a_473374_648060# a_471230_648050# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X675 esd_6/in vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X676 io_analog[5] vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X677 vssa1 vssa1 io_analog[7] vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X678 vccd1 a_504724_647182# a_505416_647172# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X679 esd_0/in a_500126_647170# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X680 vssa1 a_483446_644892# a_481708_644918# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X681 a_504724_647182# VCO_Flat_0/Buff_VCO_1/IN vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X682 vccd1 vccd1 esd_4/in vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X683 io_analog[4] vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X684 vssa1 vssa1 esd_2/in vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X685 vccd1 esd_1/in a_490818_650238# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X686 vccd1 a_473374_648060# a_471230_648050# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X687 a_473374_648060# a_475058_648060# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X688 vssa1 a_479772_646886# a_484664_644902# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X689 vssa1 a_483446_644892# a_487694_644902# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X690 vssa1 a_479772_646886# a_479772_646886# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=200000u
X691 esd_0/in vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X692 a_493938_644874# a_479772_646886# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X693 vccd1 vccd1 esd_2/in vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X694 vccd1 a_457934_648038# esd_3/in vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X695 vccd1 a_506614_647168# esd_6/in vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X696 vssa1 a_483446_644892# a_481708_644918# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X697 esd_5/in vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X698 vssa1 vssa1 esd_2/in vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X699 a_479864_646886# esd_2/in a_479772_646886# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X700 vccd1 a_457934_648038# esd_3/in vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X701 vccd1 a_461762_648050# a_460078_648050# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X702 vccd1 vccd1 esd_5/in vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X703 vccd1 vccd1 esd_2/in vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X704 vssa1 vssa1 esd_0/in vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X705 a_487730_650240# esd_1/in vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X706 vccd1 a_506614_647168# esd_6/in vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X707 io_analog[1] vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X708 esd_0/in vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X709 esd_5/in a_471230_648050# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X710 a_500126_647170# a_498928_647174# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X711 esd_5/in vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X712 vccd1 a_500126_647170# esd_0/in vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X713 vssa1 VCO_Flat_0/Buff_VCO_3/IN a_468592_648062# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X714 vccd1 vccd1 io_analog[1] vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X715 io_analog[2] vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X716 a_473374_648060# a_475058_648060# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X717 vccd1 vccd1 io_analog[5] vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X718 vssa1 vssa1 esd_0/in vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X719 a_490818_650238# VCO_Flat_0/Buff_VCO_4/IN VCO_Flat_0/Buff_VCO_1/IN vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X720 vccd1 a_505416_647172# a_506614_647168# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X721 io_analog[2] vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X722 a_498928_647174# a_498236_647184# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X723 vssa1 a_506614_647168# esd_6/in vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X724 a_500126_647170# a_498928_647174# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X725 vssa1 a_471230_648050# esd_5/in vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X726 esd_4/in a_464764_648054# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X727 esd_3/in vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X728 vccd1 vccd1 io_analog[1] vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X729 io_analog[1] vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X730 vccd1 a_466908_648062# a_464764_648054# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X731 vccd1 a_498928_647174# a_500126_647170# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X732 io_analog[3] vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X733 vccd1 vccd1 io_analog[3] vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X734 vssa1 a_457934_648038# esd_3/in vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X735 vssa1 a_506614_647168# esd_6/in vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X736 a_490782_644900# VCO_Flat_0/Buff_VCO_2/IN VCO_Flat_0/Buff_VCO_1/IN vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X737 a_498236_647184# VCO_Flat_0/Buff_VCO_0/IN vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X738 vccd1 vccd1 io_analog[3] vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X739 vssa1 vssa1 esd_3/in vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X740 vccd1 a_466908_648062# a_464764_648054# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X741 vccd1 a_498928_647174# a_500126_647170# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X742 vccd1 a_505416_647172# a_506614_647168# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X743 vssa1 a_500126_647170# esd_0/in vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X744 a_500126_647170# a_498928_647174# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X745 a_464764_648054# a_466908_648062# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X746 vssa1 vssa1 io_analog[3] vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X747 a_505416_647172# a_504724_647182# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X748 io_analog[4] vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X749 a_484700_650240# a_479864_646886# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X750 vccd1 esd_1/in a_487730_650240# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X751 a_471230_648050# a_473374_648060# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X752 vssa1 vssa1 esd_2/in vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X753 vccd1 vccd1 io_analog[3] vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X754 a_505416_647172# a_504724_647182# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X755 vssa1 a_506614_647168# esd_6/in vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X756 vssa1 a_500126_647170# esd_0/in vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X757 a_498928_647174# a_498236_647184# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X758 a_464764_648054# a_466908_648062# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X759 vccd1 vccd1 io_analog[7] vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X760 vccd1 vccd1 esd_2/in vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X761 esd_1/in vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X762 vssa1 vssa1 esd_3/in vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X763 io_analog[3] vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X764 vssa1 a_479772_646886# a_479772_646886# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=200000u
X765 vssa1 vssa1 io_analog[5] vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X766 a_490818_650238# esd_1/in vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X767 a_471230_648050# a_473374_648060# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X768 a_487694_644902# a_483446_644892# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X769 a_479772_646886# a_479772_646886# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=200000u
X770 io_analog[7] vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X771 vccd1 vccd1 esd_1/in vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X772 a_481744_650256# esd_1/in vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X773 vssa1 a_479772_646886# a_493938_644874# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X774 io_analog[7] vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X775 a_464764_648054# a_466908_648062# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X776 esd_1/in vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X777 vccd1 vccd1 esd_1/in vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X778 vccd1 VCO_Flat_0/Buff_VCO_2/IN a_475058_648060# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X779 esd_6/in a_506614_647168# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X780 a_471230_648050# a_473374_648060# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
R2 vssa1 io_clamp_low[2] sky130_fd_pr__res_generic_m3 w=1.085e+07u l=1.29e+06u
X781 esd_3/in vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X782 vssa1 vssa1 io_analog[5] vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X783 esd_4/in vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X784 a_493974_650212# VCO_Flat_0/Buff_VCO_3/IN VCO_Flat_0/Buff_VCO_0/IN vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X785 esd_6/in a_506614_647168# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X786 VCO_Flat_0/Buff_VCO_4/IN VCO_Flat_0/Buff_VCO_2/IN vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X787 io_analog[7] vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X788 vssa1 vssa1 esd_4/in vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X789 vccd1 a_471230_648050# esd_5/in vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X790 vssa1 vssa1 esd_1/in vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X791 esd_0/in a_500126_647170# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X792 vssa1 a_483446_644892# a_490782_644900# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X793 a_468592_648062# VCO_Flat_0/Buff_VCO_3/IN vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X794 vccd1 vccd1 io_analog[4] vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X795 vccd1 a_475058_648060# a_473374_648060# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X796 esd_1/in vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X797 a_460078_648050# a_461762_648050# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X798 VCO_Flat_0/Buff_VCO_1/IN VCO_Flat_0/Buff_VCO_4/IN a_490818_650238# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X799 a_506614_647168# a_505416_647172# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X800 vssa1 a_479772_646886# a_493938_644874# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X801 esd_6/in a_506614_647168# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X802 esd_5/in a_471230_648050# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X803 esd_6/in vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X804 esd_0/in a_500126_647170# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X805 io_analog[6] vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X806 a_464764_648054# a_466908_648062# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X807 a_500126_647170# a_498928_647174# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X808 a_479772_646886# esd_2/in a_479864_646886# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X809 esd_3/in vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X810 a_484700_650240# esd_1/in vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X811 a_460078_648050# a_461762_648050# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X812 VCO_Flat_0/Buff_VCO_1/IN VCO_Flat_0/Buff_VCO_2/IN a_490782_644900# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X813 vccd1 VCO_Flat_0/Buff_VCO_0/IN a_498236_647184# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X814 esd_5/in a_471230_648050# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X815 esd_6/in vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X816 vccd1 vccd1 io_analog[6] vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X817 a_506614_647168# a_505416_647172# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X818 vssa1 vssa1 esd_6/in vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X819 a_464764_648054# a_466908_648062# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X820 a_500126_647170# a_498928_647174# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X821 vssa1 a_498928_647174# a_500126_647170# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X822 vssa1 a_466908_648062# a_464764_648054# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X823 io_analog[6] vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X824 esd_5/in vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X825 vssa1 vssa1 esd_6/in vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X826 io_analog[5] vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X827 vssa1 vssa1 esd_6/in vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X828 a_484700_650240# esd_1/in vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X829 a_506614_647168# a_505416_647172# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X830 a_487694_644902# a_483446_644892# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X831 esd_6/in a_506614_647168# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X832 esd_0/in a_500126_647170# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X833 esd_5/in a_471230_648050# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X834 vssa1 a_464764_648054# esd_4/in vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X835 vccd1 vccd1 io_analog[7] vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X836 esd_4/in vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X837 vssa1 vssa1 io_analog[6] vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X838 vccd1 vccd1 io_analog[5] vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X839 a_464764_648054# a_466908_648062# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X840 a_500126_647170# a_498928_647174# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X841 esd_3/in a_457934_648038# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X842 VCO_Flat_0/Buff_VCO_0/IN VCO_Flat_0/Buff_VCO_3/IN vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X843 vccd1 vccd1 esd_4/in vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X844 io_analog[6] vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X845 vccd1 a_479864_646886# a_484700_650240# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X846 vccd1 a_473374_648060# a_471230_648050# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X847 vssa1 a_483446_644892# a_487694_644902# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
R3 vccd1 io_clamp_high[0] sky130_fd_pr__res_generic_m3 w=1.081e+07u l=1.29e+06u
X848 vccd1 vccd1 io_analog[4] vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X849 esd_4/in vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X850 io_analog[7] vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X851 a_475058_648060# VCO_Flat_0/Buff_VCO_2/IN vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X852 vccd1 a_504724_647182# a_505416_647172# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X853 esd_0/in a_500126_647170# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X854 vssa1 a_466908_648062# a_464764_648054# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X855 vccd1 vccd1 esd_0/in vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X856 vccd1 a_479864_646886# a_484700_650240# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X857 vccd1 a_473374_648060# a_471230_648050# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X858 vccd1 a_479864_646886# a_490818_650238# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X859 vccd1 esd_1/in a_490818_650238# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X860 VCO_Flat_0/Buff_VCO_0/IN VCO_Flat_0/Buff_VCO_3/IN a_493974_650212# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X861 vccd1 esd_1/in a_481744_650256# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X862 esd_0/in vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X863 vccd1 a_506614_647168# esd_6/in vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X864 vssa1 a_498236_647184# a_498928_647174# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X865 vssa1 a_505416_647172# a_506614_647168# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X866 vccd1 a_500126_647170# esd_0/in vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X867 vssa1 VCO_Flat_0/Buff_VCO_3/IN a_468592_648062# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X868 esd_0/in vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X869 io_analog[2] vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X870 vccd1 esd_1/in a_481744_650256# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X871 a_493938_644874# a_479772_646886# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X872 vssa1 a_479772_646886# a_481708_644918# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X873 io_analog[5] vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X874 io_analog[2] vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X875 vssa1 vssa1 io_analog[2] vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X876 vccd1 a_506614_647168# esd_6/in vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X877 vssa1 a_471230_648050# esd_5/in vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X878 vccd1 vccd1 io_analog[1] vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X879 io_analog[2] vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X880 vccd1 a_479864_646886# a_493974_650212# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X881 vccd1 a_500126_647170# esd_0/in vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X882 vssa1 a_504724_647182# a_505416_647172# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X883 vccd1 vccd1 esd_5/in vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X884 vccd1 vccd1 io_analog[2] vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X885 io_analog[2] vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X886 io_analog[2] vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X887 vccd1 a_461762_648050# a_460078_648050# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X888 a_490782_644900# a_483446_644892# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X889 esd_0/in vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X890 vssa1 a_504724_647182# a_505416_647172# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X891 io_analog[2] vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X892 vccd1 a_479864_646886# a_493974_650212# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X893 vccd1 a_464764_648054# esd_4/in vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X894 esd_5/in a_471230_648050# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X895 vccd1 a_498928_647174# a_500126_647170# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X896 vccd1 a_505416_647172# a_506614_647168# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X897 vccd1 vccd1 io_analog[1] vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X898 vssa1 a_471230_648050# esd_5/in vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X899 vccd1 vccd1 esd_3/in vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X900 vccd1 a_468592_648062# a_466908_648062# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X901 vccd1 a_500126_647170# esd_0/in vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X902 vccd1 esd_1/in a_484700_650240# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X903 vccd1 a_505416_647172# a_506614_647168# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X904 vssa1 a_483446_644892# a_487694_644902# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X905 io_analog[4] vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X906 vssa1 a_471230_648050# esd_5/in vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X907 esd_4/in a_464764_648054# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X908 io_analog[3] vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X909 io_analog[1] vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X910 vccd1 a_464764_648054# esd_4/in vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X911 a_457934_648038# a_460078_648050# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X912 vccd1 a_466908_648062# a_464764_648054# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X913 vccd1 a_498928_647174# a_500126_647170# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X914 io_analog[7] vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X915 io_analog[1] vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X916 vccd1 a_468592_648062# a_466908_648062# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X917 vssa1 a_457934_648038# esd_3/in vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X918 esd_4/in a_464764_648054# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X919 io_analog[3] vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X920 a_484664_644902# a_483446_644892# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X921 a_487730_650240# a_479864_646886# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X922 a_473374_648060# a_475058_648060# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X923 a_457934_648038# a_460078_648050# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X924 vccd1 vccd1 io_analog[7] vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X925 vssa1 vssa1 esd_2/in vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X926 vccd1 VCO_Flat_0/Buff_VCO_2/IN a_475058_648060# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X927 a_464764_648054# a_466908_648062# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X928 esd_1/in vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X929 esd_3/in vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X930 vccd1 vccd1 esd_2/in vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X931 vssa1 vssa1 io_analog[3] vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X932 a_481744_650256# esd_1/in vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X933 a_490818_650238# a_479864_646886# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X934 esd_1/in vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X935 a_481744_650256# a_479864_646886# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X936 a_481744_650256# a_479864_646886# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X937 a_484700_650240# VCO_Flat_0/Buff_VCO_1/IN VCO_Flat_0/Buff_VCO_3/IN vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X938 vssa1 a_506614_647168# esd_6/in vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X939 vssa1 vssa1 esd_2/in vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X940 a_498928_647174# a_498236_647184# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X941 io_analog[3] vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X942 a_506614_647168# a_505416_647172# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X943 vccd1 vccd1 esd_2/in vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X944 vssa1 vssa1 io_analog[5] vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X945 vssa1 a_457934_648038# esd_3/in vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X946 vssa1 vssa1 esd_1/in vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X947 a_490818_650238# esd_1/in vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X948 a_506614_647168# a_505416_647172# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X949 a_484664_644902# VCO_Flat_0/Buff_VCO_4/IN VCO_Flat_0/Buff_VCO_3/IN vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X950 a_481744_650256# esd_1/in vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X951 a_481708_644918# a_479772_646886# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X952 vccd1 vccd1 io_analog[4] vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X953 a_505416_647172# a_504724_647182# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X954 a_493974_650212# a_479864_646886# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X955 a_460078_648050# a_461762_648050# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X956 vssa1 vssa1 esd_4/in vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X957 vssa1 a_483446_644892# a_490782_644900# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X958 a_505416_647172# a_504724_647182# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X959 io_analog[4] vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X960 vccd1 a_471230_648050# esd_5/in vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X961 io_analog[6] vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X962 esd_0/in a_500126_647170# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X963 a_484700_650240# esd_1/in vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X964 a_493974_650212# a_479864_646886# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X965 io_analog[6] vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X966 vccd1 a_471230_648050# esd_5/in vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X967 a_487694_644902# a_483446_644892# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X968 vssa1 a_464764_648054# esd_4/in vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X969 esd_5/in vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X970 esd_6/in a_506614_647168# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X971 a_505416_647172# a_504724_647182# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X972 esd_5/in a_471230_648050# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X973 vccd1 vccd1 io_analog[5] vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X974 vssa1 vssa1 esd_5/in vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X975 a_493974_650212# a_479864_646886# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X976 esd_4/in a_464764_648054# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X977 vssa1 a_460078_648050# a_457934_648038# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X978 esd_6/in vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X979 io_analog[7] vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X980 esd_6/in vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X981 vssa1 vssa1 io_analog[6] vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X982 a_466908_648062# a_468592_648062# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X983 vssa1 a_464764_648054# esd_4/in vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X984 io_analog[5] vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X985 esd_4/in a_464764_648054# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X986 esd_5/in vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X987 vccd1 a_471230_648050# esd_5/in vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X988 a_500126_647170# a_498928_647174# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X989 vssa1 a_475058_648060# a_473374_648060# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X990 esd_4/in vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X991 vssa1 vssa1 esd_6/in vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X992 vssa1 vssa1 io_analog[5] vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X993 a_504724_647182# VCO_Flat_0/Buff_VCO_1/IN vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X994 vssa1 vssa1 io_analog[7] vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X995 io_analog[5] vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X996 io_analog[7] vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X997 vssa1 vssa1 io_analog[6] vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X998 vccd1 a_479864_646886# a_481744_650256# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X999 vccd1 a_479864_646886# a_490818_650238# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1000 vccd1 a_457934_648038# esd_3/in vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1001 esd_4/in a_464764_648054# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1002 esd_4/in vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1003 esd_3/in a_457934_648038# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1004 a_493938_644874# a_483446_644892# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1005 esd_6/in a_506614_647168# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1006 vssa1 a_475058_648060# a_473374_648060# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1007 vssa1 a_464764_648054# esd_4/in vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1008 vssa1 vssa1 io_analog[6] vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1009 vssa1 a_498236_647184# a_498928_647174# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1010 vccd1 VCO_Flat_0/Buff_VCO_4/IN a_461762_648050# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1011 vssa1 a_460078_648050# a_457934_648038# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1012 esd_2/in vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1013 esd_3/in a_457934_648038# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1014 esd_2/in vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1015 vccd1 esd_1/in a_481744_650256# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1016 vssa1 a_479772_646886# a_481708_644918# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1017 vssa1 a_505416_647172# a_506614_647168# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1018 vssa1 a_475058_648060# a_473374_648060# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1019 vssa1 a_460078_648050# a_457934_648038# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1020 vccd1 vccd1 io_analog[4] vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1021 vssa1 vssa1 io_analog[2] vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1022 vccd1 a_479864_646886# a_490818_650238# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1023 vssa1 a_479772_646886# a_487694_644902# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1024 vccd1 vccd1 esd_0/in vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1025 vccd1 vccd1 io_analog[2] vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1026 vssa1 vssa1 io_analog[2] vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1027 vccd1 a_479864_646886# a_481744_650256# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1028 a_493974_650212# esd_1/in vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1029 io_analog[1] vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1030 vssa1 VCO_Flat_0/Buff_VCO_2/IN a_475058_648060# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1031 vccd1 vccd1 io_analog[2] vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1032 vssa1 a_504724_647182# a_505416_647172# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1033 VCO_Flat_0/Buff_VCO_3/IN VCO_Flat_0/Buff_VCO_4/IN a_484664_644902# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1034 vccd1 vccd1 esd_5/in vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1035 io_analog[1] vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1036 vssa1 a_479772_646886# a_481708_644918# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1037 esd_0/in vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1038 vccd1 VCO_Flat_0/Buff_VCO_3/IN a_468592_648062# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1039 vccd1 vccd1 esd_5/in vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1040 vccd1 a_479864_646886# a_479864_646886# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=200000u
X1041 vccd1 vccd1 io_analog[1] vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1042 a_479864_646886# a_479864_646886# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=200000u
X1043 vssa1 a_479772_646886# a_481708_644918# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1044 vssa1 a_505416_647172# a_506614_647168# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1045 vccd1 vccd1 esd_3/in vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1046 vccd1 vccd1 esd_5/in vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1047 vccd1 a_506614_647168# esd_6/in vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1048 vssa1 a_504724_647182# a_505416_647172# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1049 vccd1 a_479864_646886# a_493974_650212# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1050 esd_5/in a_471230_648050# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1051 io_analog[3] vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1052 io_analog[1] vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1053 vccd1 a_468592_648062# a_466908_648062# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1054 a_490782_644900# a_483446_644892# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1055 vccd1 vccd1 esd_3/in vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1056 vccd1 a_464764_648054# esd_4/in vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1057 vssa1 vssa1 io_analog[1] vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1058 esd_5/in a_471230_648050# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1059 io_analog[3] vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1060 vssa1 vssa1 io_analog[4] vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1061 esd_2/in vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1062 vccd1 a_468592_648062# a_466908_648062# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1063 vccd1 a_500126_647170# esd_0/in vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1064 esd_3/in a_457934_648038# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1065 esd_2/in vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1066 vssa1 vssa1 io_analog[1] vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1067 a_481744_650256# a_479864_646886# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1068 vccd1 a_464764_648054# esd_4/in vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1069 VCO_Flat_0/Buff_VCO_0/IN VCO_Flat_0/Buff_VCO_1/IN a_493938_644874# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1070 esd_3/in vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1071 vssa1 a_483446_644892# a_493938_644874# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1072 esd_4/in a_464764_648054# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1073 io_analog[3] vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1074 vssa1 vssa1 io_analog[3] vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1075 vssa1 a_461762_648050# a_460078_648050# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1076 esd_2/in vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1077 a_461762_648050# VCO_Flat_0/Buff_VCO_4/IN vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1078 a_457934_648038# a_460078_648050# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1079 esd_2/in vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1080 vssa1 vssa1 io_analog[3] vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1081 vccd1 vccd1 esd_1/in vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1082 esd_5/in io_analog[5] vssa1 sky130_fd_pr__res_high_po w=2.85e+06u l=1.3e+06u
X1083 esd_3/in a_457934_648038# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1084 a_484664_644902# a_483446_644892# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1085 vssa1 a_483446_644892# a_493938_644874# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1086 vssa1 a_500126_647170# esd_0/in vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1087 a_473374_648060# a_475058_648060# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1088 a_457934_648038# a_460078_648050# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1089 vssa1 a_461762_648050# a_460078_648050# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1090 vccd1 vccd1 io_analog[7] vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1091 esd_1/in vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1092 io_analog[5] vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1093 vssa1 vssa1 io_analog[3] vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1094 a_490818_650238# a_479864_646886# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1095 esd_3/in a_457934_648038# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1096 a_487694_644902# a_479772_646886# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1097 vssa1 vssa1 io_analog[7] vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1098 esd_4/in vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1099 a_481744_650256# a_479864_646886# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1100 vccd1 a_460078_648050# a_457934_648038# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1101 esd_1/in vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1102 vssa1 vssa1 io_analog[5] vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1103 a_506614_647168# a_505416_647172# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1104 vssa1 vssa1 esd_4/in vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1105 a_487694_644902# a_479772_646886# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1106 io_analog[7] vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1107 vssa1 vssa1 io_analog[4] vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1108 vssa1 vssa1 esd_1/in vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1109 vccd1 a_506614_647168# esd_6/in vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1110 esd_4/in vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1111 vccd1 vccd1 esd_6/in vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1112 esd_1/in vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1113 vssa1 vssa1 esd_1/in vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1114 a_481708_644918# a_479772_646886# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1115 a_506614_647168# a_505416_647172# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1116 vccd1 vccd1 esd_3/in vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1117 io_analog[4] vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1118 esd_3/in vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1119 esd_6/in a_506614_647168# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1120 vssa1 a_479772_646886# a_490782_644900# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1121 vssa1 a_483446_644892# a_490782_644900# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1122 vccd1 vccd1 io_analog[6] vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1123 io_analog[7] vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1124 vssa1 a_506614_647168# esd_6/in vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1125 a_471230_648050# a_473374_648060# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1126 esd_0/in a_500126_647170# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1127 io_analog[6] vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1128 esd_6/in vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1129 io_analog[5] vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1130 esd_4/in a_464764_648054# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1131 vccd1 vccd1 io_analog[5] vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1132 io_analog[6] vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1133 a_479864_646886# a_479864_646886# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=200000u
X1134 vssa1 vssa1 esd_5/in vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1135 a_460078_648050# a_461762_648050# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1136 vccd1 vccd1 esd_4/in vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1137 vccd1 vccd1 io_analog[5] vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1138 esd_6/in vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1139 vssa1 vssa1 io_analog[6] vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1140 vccd1 vccd1 esd_4/in vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1141 vssa1 a_483446_644892# a_484664_644902# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1142 io_analog[6] vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1143 esd_4/in a_464764_648054# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
R4 vssa1 io_clamp_low[0] sky130_fd_pr__res_generic_m3 w=1.082e+07u l=1.29e+06u
X1144 vssa1 a_460078_648050# a_457934_648038# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1145 io_analog[5] vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1146 vccd1 a_479864_646886# a_487730_650240# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1147 a_493938_644874# a_483446_644892# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1148 esd_4/in vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1149 a_460078_648050# a_461762_648050# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1150 vccd1 vccd1 esd_0/in vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1151 io_analog[4] vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1152 vccd1 a_457934_648038# esd_3/in vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1153 vccd1 vccd1 io_analog[4] vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1154 vssa1 vssa1 io_analog[7] vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1155 vccd1 a_479864_646886# a_481744_650256# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1156 a_457934_648038# a_460078_648050# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1157 a_493938_644874# a_483446_644892# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1158 vssa1 a_464764_648054# esd_4/in vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1159 a_460078_648050# a_461762_648050# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1160 vccd1 vccd1 esd_0/in vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1161 vssa1 a_483446_644892# a_484664_644902# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1162 esd_6/in a_506614_647168# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1163 vssa1 a_479772_646886# a_487694_644902# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1164 esd_5/in vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1165 vssa1 vssa1 esd_0/in vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1166 a_483446_644892# esd_1/in vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=150000u
X1167 vssa1 a_471230_648050# esd_5/in vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1168 a_466908_648062# a_468592_648062# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1169 a_461762_648050# VCO_Flat_0/Buff_VCO_4/IN vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1170 vccd1 vccd1 esd_5/in vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1171 vssa1 vssa1 io_analog[2] vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1172 esd_0/in vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1173 vccd1 vccd1 io_analog[2] vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1174 vccd1 vccd1 esd_1/in vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1175 a_457934_648038# a_460078_648050# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1176 a_490782_644900# a_483446_644892# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1177 vssa1 VCO_Flat_0/Buff_VCO_2/IN a_475058_648060# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1178 io_analog[1] vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1179 vssa1 a_473374_648060# a_471230_648050# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1180 a_498236_647184# VCO_Flat_0/Buff_VCO_0/IN vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1181 vccd1 vccd1 io_analog[3] vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1182 vccd1 vccd1 io_analog[1] vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1183 a_490782_644900# a_479772_646886# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1184 vssa1 vssa1 io_analog[4] vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1185 vssa1 vssa1 io_analog[1] vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1186 vssa1 a_473374_648060# a_471230_648050# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1187 a_464764_648054# a_466908_648062# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1188 esd_3/in vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1189 vccd1 a_506614_647168# esd_6/in vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1190 vccd1 vccd1 io_analog[3] vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1191 a_490782_644900# a_479772_646886# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1192 esd_2/in vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1193 vssa1 vssa1 io_analog[1] vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1194 io_analog[3] vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1195 vssa1 vssa1 esd_3/in vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1196 a_487730_650240# a_479864_646886# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1197 a_479772_646886# esd_2/in a_479864_646886# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1198 esd_2/in vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1199 vccd1 vccd1 esd_1/in vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1200 vccd1 VCO_Flat_0/Buff_VCO_3/IN a_468592_648062# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1201 io_analog[7] vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1202 vssa1 vssa1 io_analog[5] vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1203 io_analog[3] vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1204 vccd1 a_460078_648050# a_457934_648038# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1205 a_484664_644902# a_483446_644892# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1206 a_481708_644918# a_483446_644892# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1207 esd_4/in a_464764_648054# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1208 vssa1 a_461762_648050# a_460078_648050# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1209 io_analog[7] vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1210 io_analog[3] vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1211 io_analog[5] vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1212 a_484664_644902# a_479772_646886# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1213 vccd1 vccd1 esd_1/in vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1214 vssa1 vssa1 io_analog[7] vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1215 esd_4/in vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1216 esd_1/in vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1217 esd_5/in a_471230_648050# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1218 vssa1 a_468592_648062# a_466908_648062# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1219 vssa1 VCO_Flat_0/Buff_VCO_4/IN a_461762_648050# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1220 io_analog[5] vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1221 a_481708_644918# a_483446_644892# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1222 esd_3/in vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1223 esd_1/in vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1224 vccd1 vccd1 esd_3/in vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1225 esd_4/in vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1226 esd_3/in a_457934_648038# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1227 vccd1 a_460078_648050# a_457934_648038# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1228 vccd1 esd_1/in a_493974_650212# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1229 vccd1 vssa1 a_483446_644892# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X1230 vssa1 a_498928_647174# a_500126_647170# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1231 a_471230_648050# a_473374_648060# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1232 vssa1 a_468592_648062# a_466908_648062# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1233 vccd1 vccd1 esd_6/in vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1234 vccd1 a_460078_648050# a_457934_648038# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1235 vccd1 vccd1 io_analog[6] vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1236 vssa1 vssa1 io_analog[4] vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1237 vccd1 a_498236_647184# a_498928_647174# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1238 esd_6/in a_506614_647168# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1239 a_471230_648050# a_473374_648060# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1240 esd_5/in a_471230_648050# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1241 vssa1 a_466908_648062# a_464764_648054# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1242 vccd1 vccd1 esd_6/in vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1243 vccd1 vccd1 io_analog[6] vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1244 vssa1 a_479772_646886# a_490782_644900# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1245 vccd1 vccd1 io_analog[5] vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1246 esd_3/in a_457934_648038# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1247 esd_6/in a_506614_647168# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1248 vccd1 vccd1 io_analog[6] vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1249 vssa1 vssa1 esd_5/in vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1250 a_498236_647184# VCO_Flat_0/Buff_VCO_0/IN vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1251 io_analog[6] vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1252 esd_0/in a_500126_647170# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1253 a_479864_646886# esd_2/in a_479772_646886# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1254 vssa1 vssa1 esd_5/in vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1255 vccd1 a_479864_646886# a_484700_650240# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1256 io_analog[6] vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1257 a_487730_650240# esd_1/in vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1258 vssa1 vssa1 esd_5/in vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1259 a_468592_648062# VCO_Flat_0/Buff_VCO_3/IN vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1260 vccd1 a_504724_647182# a_505416_647172# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1261 io_analog[4] vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1262 esd_6/in vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1263 io_analog[7] vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1264 esd_0/in vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1265 vccd1 a_479864_646886# a_487730_650240# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1266 vssa1 a_479772_646886# a_484664_644902# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1267 vccd1 vccd1 esd_4/in vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1268 a_493938_644874# a_479772_646886# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1269 a_493938_644874# a_479772_646886# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
R5 vccd1 io_clamp_high[2] sky130_fd_pr__res_generic_m3 w=1.08e+07u l=1.29e+06u
X1270 vccd1 a_479864_646886# a_487730_650240# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1271 a_466908_648062# a_468592_648062# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1272 esd_0/in vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1273 vssa1 a_483446_644892# a_481708_644918# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1274 esd_2/in vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1275 vccd1 a_457934_648038# esd_3/in vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1276 a_457934_648038# a_460078_648050# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1277 vssa1 a_479772_646886# a_484664_644902# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1278 esd_0/in vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1279 vccd1 vccd1 esd_0/in vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1280 a_493974_650212# esd_1/in vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1281 a_483446_644892# vssa1 vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X1282 esd_2/in vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1283 vssa1 vssa1 io_analog[2] vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1284 esd_5/in a_471230_648050# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1285 a_500126_647170# a_498928_647174# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1286 a_466908_648062# a_468592_648062# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1287 vccd1 vccd1 io_analog[2] vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1288 vccd1 vccd1 io_analog[1] vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1289 a_457934_648038# a_460078_648050# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1290 a_473374_648060# a_475058_648060# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1291 io_analog[1] vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1292 esd_5/in vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1293 a_498928_647174# a_498236_647184# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1294 a_479772_646886# a_479772_646886# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=200000u
X1295 vssa1 a_471230_648050# esd_5/in vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1296 vssa1 vssa1 esd_0/in vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1297 vccd1 a_466908_648062# a_464764_648054# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1298 vccd1 a_466908_648062# a_464764_648054# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1299 vccd1 a_498928_647174# a_500126_647170# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1300 a_479864_646886# esd_2/in a_479772_646886# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1301 io_analog[1] vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1302 a_490782_644900# a_479772_646886# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1303 esd_3/in vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1304 io_analog[1] vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1305 vssa1 a_457934_648038# esd_3/in vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1306 vssa1 VCO_Flat_0/Buff_VCO_0/IN a_498236_647184# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1307 io_analog[1] vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1308 vccd1 a_466908_648062# a_464764_648054# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1309 vssa1 a_500126_647170# esd_0/in vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1310 a_500126_647170# a_498928_647174# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1311 esd_3/in vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1312 vssa1 vssa1 io_analog[1] vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1313 a_484700_650240# a_479864_646886# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1314 vccd1 esd_1/in a_487730_650240# vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1315 vccd1 vccd1 io_analog[3] vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1316 vssa1 vssa1 esd_3/in vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1317 a_505416_647172# a_504724_647182# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1318 vssa1 a_506614_647168# esd_6/in vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1319 vssa1 a_500126_647170# esd_0/in vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1320 a_500126_647170# a_498928_647174# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1321 io_analog[4] vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1322 vssa1 vssa1 esd_2/in vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1323 vssa1 a_473374_648060# a_471230_648050# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1324 a_468592_648062# VCO_Flat_0/Buff_VCO_3/IN vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1325 vccd1 vccd1 esd_2/in vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1326 io_analog[3] vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1327 vccd1 vccd1 esd_1/in vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1328 vssa1 vssa1 esd_3/in vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1329 a_484700_650240# a_479864_646886# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1330 a_471230_648050# a_473374_648060# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1331 a_484664_644902# a_479772_646886# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1332 a_487694_644902# a_483446_644892# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1333 vssa1 a_506614_647168# esd_6/in vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1334 VCO_Flat_0/Buff_VCO_1/IN VCO_Flat_0/Buff_VCO_4/IN vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1335 vssa1 a_479772_646886# a_493938_644874# vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1336 io_analog[3] vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1337 vccd1 a_464764_648054# esd_4/in vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1338 vssa1 a_500126_647170# esd_0/in vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1339 vccd1 vccd1 io_analog[7] vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1340 vssa1 vssa1 esd_2/in vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1341 a_505416_647172# a_504724_647182# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1342 a_481708_644918# a_483446_644892# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1343 vccd1 vccd1 esd_2/in vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1344 vccd1 vccd1 esd_1/in vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1345 a_484700_650240# a_479864_646886# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1346 a_490818_650238# esd_1/in vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1347 a_471230_648050# a_473374_648060# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1348 esd_3/in a_457934_648038# vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1349 a_487730_650240# VCO_Flat_0/Buff_VCO_0/IN VCO_Flat_0/Buff_VCO_2/IN vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1350 a_493974_650212# VCO_Flat_0/Buff_VCO_3/IN VCO_Flat_0/Buff_VCO_0/IN vccd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1351 esd_1/in vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1352 vssa1 vssa1 io_analog[5] vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1353 a_484664_644902# a_479772_646886# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
C0 io_analog[2] vccd1 26.70fF
C1 a_466908_648062# a_468592_648062# 1.00fF
C2 vccd1 a_490818_650238# 34.67fF
C3 a_490782_644900# a_483446_644892# 0.45fF
C4 VCO_Flat_0/Buff_VCO_0/IN a_487730_650240# 0.17fF
C5 a_484700_650240# vccd1 34.66fF
C6 esd_4/in VCO_Flat_0/Buff_VCO_4/IN 1.58fF
C7 VCO_Flat_0/Buff_VCO_2/IN a_475058_648060# 0.40fF
C8 a_466908_648062# VCO_Flat_0/Buff_VCO_4/IN 0.99fF
C9 a_457934_648038# a_460078_648050# 0.82fF
C10 VCO_Flat_0/Buff_VCO_3/IN a_493974_650212# 0.17fF
C11 a_481744_650256# VCO_Flat_0/Buff_VCO_4/IN 6.48fF
C12 a_479864_646886# a_493974_650212# 0.02fF
C13 VCO_Flat_0/Buff_VCO_2/IN VCO_Flat_0/Buff_VCO_0/IN 2.96fF
C14 a_481708_644918# a_483446_644892# 0.45fF
C15 VCO_Flat_0/Buff_VCO_4/IN esd_5/in 1.10fF
C16 a_479864_646886# a_479772_646886# 13.59fF
C17 a_481708_644918# VCO_Flat_0/Buff_VCO_0/IN 0.02fF
C18 io_analog[4] io_clamp_low[0] 3.96fF
C19 VCO_Flat_0/Buff_VCO_2/IN VCO_Flat_0/Buff_VCO_4/IN 3.68fF
C20 a_471230_648050# esd_5/in 2.28fF
C21 a_490782_644900# a_487694_644902# 0.25fF
C22 io_clamp_low[1] io_clamp_high[1] 0.81fF
C23 a_481708_644918# VCO_Flat_0/Buff_VCO_4/IN 6.58fF
C24 a_505416_647172# a_506614_647168# 0.82fF
C25 VCO_Flat_0/Buff_VCO_2/IN a_487694_644902# 6.58fF
C26 a_479772_646886# esd_2/in 0.28fF
C27 esd_1/in VCO_Flat_0/Buff_VCO_1/IN 0.44fF
C28 a_457934_648038# esd_3/in 2.28fF
C29 a_498928_647174# vccd1 17.68fF
C30 a_464764_648054# esd_4/in 2.28fF
C31 a_464764_648054# a_466908_648062# 0.82fF
C32 io_analog[3] vccd1 26.68fF
C33 a_498236_647184# VCO_Flat_0/Buff_VCO_0/IN 0.40fF
C34 a_479864_646886# esd_1/in 1.17fF
C35 vccd1 VCO_Flat_0/Buff_VCO_1/IN 0.33fF
C36 VCO_Flat_0/Buff_VCO_0/IN a_483446_644892# 0.06fF
C37 VCO_Flat_0/Buff_VCO_3/IN vccd1 1.23fF
C38 m3_173410_700370# io_clamp_low[2] 0.00fF
C39 a_479864_646886# vccd1 23.05fF
C40 VCO_Flat_0/Buff_VCO_1/IN a_504724_647182# 0.40fF
C41 a_475058_648060# VCO_Flat_0/Buff_VCO_4/IN 0.47fF
C42 esd_1/in esd_2/in 1.17fF
C43 a_468592_648062# VCO_Flat_0/Buff_VCO_4/IN 0.61fF
C44 vccd1 io_analog[7] 26.76fF
C45 VCO_Flat_0/Buff_VCO_0/IN VCO_Flat_0/Buff_VCO_4/IN 4.75fF
C46 vccd1 esd_2/in 56.36fF
C47 a_473374_648060# vccd1 17.71fF
C48 a_483446_644892# a_487694_644902# 0.45fF
C49 a_490782_644900# a_479772_646886# 0.51fF
C50 VCO_Flat_0/Buff_VCO_3/IN a_484664_644902# 6.59fF
C51 io_analog[5] io_clamp_low[1] 3.96fF
C52 vccd1 a_500126_647170# 27.24fF
C53 VCO_Flat_0/Buff_VCO_1/IN a_490818_650238# 6.49fF
C54 esd_6/in esd_1/in 0.74fF
C55 a_460078_648050# vccd1 17.69fF
C56 a_484700_650240# VCO_Flat_0/Buff_VCO_1/IN 0.16fF
C57 a_479864_646886# a_490818_650238# 0.02fF
C58 a_471230_648050# VCO_Flat_0/Buff_VCO_4/IN 1.15fF
C59 VCO_Flat_0/Buff_VCO_2/IN a_479772_646886# 0.10fF
C60 a_493938_644874# VCO_Flat_0/Buff_VCO_1/IN 0.02fF
C61 VCO_Flat_0/Buff_VCO_3/IN a_484700_650240# 6.48fF
C62 a_479864_646886# a_484700_650240# 0.02fF
C63 esd_6/in vccd1 52.65fF
C64 vccd1 io_analog[6] 26.87fF
C65 a_479772_646886# a_481708_644918# 0.51fF
C66 a_506614_647168# vccd1 27.23fF
C67 a_460078_648050# a_461762_648050# 1.00fF
C68 esd_4/in vccd1 52.65fF
C69 a_466908_648062# vccd1 17.70fF
C70 io_analog[2] esd_2/in 0.50fF
C71 vccd1 a_487730_650240# 34.66fF
C72 a_481744_650256# vccd1 34.72fF
C73 vccd1 esd_5/in 53.10fF
C74 a_464764_648054# VCO_Flat_0/Buff_VCO_4/IN 1.51fF
C75 vccd1 esd_3/in 52.65fF
C76 io_analog[4] vccd1 26.68fF
C77 VCO_Flat_0/Buff_VCO_2/IN vccd1 0.06fF
C78 io_clamp_low[2] io_analog[6] 3.81fF
C79 a_493974_650212# VCO_Flat_0/Buff_VCO_0/IN 6.48fF
C80 a_479772_646886# a_483446_644892# 4.73fF
C81 io_analog[1] esd_1/in 0.50fF
C82 io_analog[5] esd_5/in 0.50fF
C83 io_analog[1] vccd1 26.75fF
C84 vccd1 m3_170914_700368# 0.00fF
C85 VCO_Flat_0/Buff_VCO_3/IN VCO_Flat_0/Buff_VCO_1/IN 0.74fF
C86 a_479864_646886# VCO_Flat_0/Buff_VCO_3/IN 0.08fF
C87 esd_0/in esd_1/in 0.74fF
C88 a_490782_644900# a_493938_644874# 0.20fF
C89 esd_1/in a_483446_644892# 0.17fF
C90 a_498236_647184# vccd1 9.22fF
C91 a_481708_644918# a_484664_644902# 0.84fF
C92 a_479772_646886# a_487694_644902# 0.51fF
C93 esd_1/in VCO_Flat_0/Buff_VCO_0/IN 0.18fF
C94 esd_0/in vccd1 52.65fF
C95 a_483446_644892# vccd1 5.82fF
C96 vccd1 a_475058_648060# 9.21fF
C97 a_468592_648062# vccd1 9.21fF
C98 a_498928_647174# a_500126_647170# 0.82fF
C99 m3_324320_700392# m3_326806_700392# 0.05fF
C100 VCO_Flat_0/Buff_VCO_0/IN vccd1 0.14fF
C101 a_479864_646886# esd_2/in 0.53fF
C102 vccd1 VCO_Flat_0/Buff_VCO_4/IN 1.58fF
C103 io_clamp_low[2] io_clamp_high[2] 0.85fF
C104 a_471230_648050# vccd1 27.24fF
C105 a_483446_644892# a_484664_644902# 0.45fF
C106 io_analog[4] io_clamp_high[0] 3.96fF
C107 a_461762_648050# VCO_Flat_0/Buff_VCO_4/IN 0.40fF
C108 a_457934_648038# vccd1 27.23fF
C109 a_479864_646886# a_487730_650240# 0.02fF
C110 a_490782_644900# VCO_Flat_0/Buff_VCO_1/IN 6.60fF
C111 a_493938_644874# a_483446_644892# 0.77fF
C112 esd_6/in io_analog[7] 0.50fF
C113 a_479864_646886# a_481744_650256# 0.07fF
C114 io_analog[3] esd_3/in 0.50fF
C115 a_484664_644902# VCO_Flat_0/Buff_VCO_4/IN 0.02fF
C116 m3_170914_700368# m3_173410_700370# 0.05fF
C117 esd_6/in esd_2/in 0.85fF
C118 a_493938_644874# VCO_Flat_0/Buff_VCO_0/IN 6.81fF
C119 VCO_Flat_0/Buff_VCO_3/IN esd_5/in 0.02fF
C120 a_505416_647172# vccd1 17.69fF
C121 VCO_Flat_0/Buff_VCO_2/IN VCO_Flat_0/Buff_VCO_1/IN 1.42fF
C122 VCO_Flat_0/Buff_VCO_4/IN a_490818_650238# 0.17fF
C123 VCO_Flat_0/Buff_VCO_3/IN VCO_Flat_0/Buff_VCO_2/IN 0.72fF
C124 a_464764_648054# vccd1 27.24fF
C125 a_484664_644902# a_487694_644902# 0.31fF
C126 a_505416_647172# a_504724_647182# 1.04fF
C127 a_493974_650212# esd_1/in 0.01fF
C128 a_493974_650212# vccd1 34.68fF
C129 a_506614_647168# esd_6/in 1.73fF
C130 VCO_Flat_0/Buff_VCO_2/IN esd_2/in 0.45fF
C131 a_498236_647184# a_498928_647174# 1.00fF
C132 io_clamp_low[0] io_clamp_high[0] 0.85fF
C133 esd_0/in VCO_Flat_0/Buff_VCO_1/IN 0.23fF
C134 io_analog[5] io_clamp_high[1] 3.96fF
C135 a_483446_644892# VCO_Flat_0/Buff_VCO_1/IN 0.06fF
C136 a_468592_648062# VCO_Flat_0/Buff_VCO_3/IN 0.40fF
C137 VCO_Flat_0/Buff_VCO_0/IN VCO_Flat_0/Buff_VCO_1/IN 1.94fF
C138 VCO_Flat_0/Buff_VCO_3/IN VCO_Flat_0/Buff_VCO_0/IN 1.72fF
C139 io_analog[4] esd_4/in 0.50fF
C140 esd_1/in vccd1 36.97fF
C141 VCO_Flat_0/Buff_VCO_2/IN a_487730_650240# 6.48fF
C142 VCO_Flat_0/Buff_VCO_1/IN VCO_Flat_0/Buff_VCO_4/IN 1.94fF
C143 a_479772_646886# a_484664_644902# 0.51fF
C144 VCO_Flat_0/Buff_VCO_2/IN a_481744_650256# 0.16fF
C145 VCO_Flat_0/Buff_VCO_3/IN VCO_Flat_0/Buff_VCO_4/IN 5.50fF
C146 m3_222608_700522# m3_225118_700522# 0.05fF
C147 esd_0/in esd_2/in 0.84fF
C148 a_490782_644900# VCO_Flat_0/Buff_VCO_2/IN 0.02fF
C149 a_479864_646886# VCO_Flat_0/Buff_VCO_4/IN 0.10fF
C150 a_473374_648060# a_475058_648060# 1.00fF
C151 esd_0/in a_500126_647170# 2.28fF
C152 a_493938_644874# a_479772_646886# 0.45fF
C153 VCO_Flat_0/Buff_VCO_3/IN a_487694_644902# 0.02fF
C154 vccd1 a_504724_647182# 9.23fF
C155 io_analog[5] vccd1 27.14fF
C156 vccd1 a_461762_648050# 9.21fF
C157 io_clamp_high[2] io_analog[6] 3.81fF
C158 VCO_Flat_0/Buff_VCO_4/IN esd_2/in 0.20fF
C159 a_473374_648060# VCO_Flat_0/Buff_VCO_4/IN 0.76fF
C160 esd_0/in io_analog[6] 0.50fF
C161 a_471230_648050# a_473374_648060# 0.82fF
C162 io_in_3v3[0] vssa1 0.61fF
C163 io_oeb[26] vssa1 0.61fF
C164 io_in[0] vssa1 0.61fF
C165 io_out[26] vssa1 0.61fF
C166 io_out[0] vssa1 0.61fF
C167 io_in[26] vssa1 0.61fF
C168 io_oeb[0] vssa1 0.61fF
C169 io_in_3v3[26] vssa1 0.61fF
C170 io_in_3v3[1] vssa1 0.61fF
C171 io_oeb[25] vssa1 0.61fF
C172 io_in[1] vssa1 0.61fF
C173 io_out[25] vssa1 0.61fF
C174 io_out[1] vssa1 0.61fF
C175 io_in[25] vssa1 0.61fF
C176 io_oeb[1] vssa1 0.61fF
C177 io_in_3v3[25] vssa1 0.61fF
C178 io_in_3v3[2] vssa1 0.61fF
C179 io_oeb[24] vssa1 0.61fF
C180 io_in[2] vssa1 0.61fF
C181 io_out[24] vssa1 0.61fF
C182 io_out[2] vssa1 0.61fF
C183 io_in[24] vssa1 0.61fF
C184 io_oeb[2] vssa1 0.61fF
C185 io_in_3v3[24] vssa1 0.61fF
C186 io_in_3v3[3] vssa1 0.61fF
C187 gpio_noesd[17] vssa1 0.61fF
C188 io_in[3] vssa1 0.61fF
C189 gpio_analog[17] vssa1 0.61fF
C190 io_out[3] vssa1 0.61fF
C191 io_oeb[3] vssa1 0.61fF
C192 io_in_3v3[4] vssa1 0.61fF
C193 io_in[4] vssa1 0.61fF
C194 io_out[4] vssa1 0.61fF
C195 io_oeb[4] vssa1 0.61fF
C196 io_oeb[23] vssa1 0.61fF
C197 io_out[23] vssa1 0.61fF
C198 io_in[23] vssa1 0.61fF
C199 io_in_3v3[23] vssa1 0.61fF
C200 gpio_noesd[16] vssa1 0.61fF
C201 gpio_analog[16] vssa1 0.61fF
C202 io_in_3v3[5] vssa1 0.61fF
C203 io_in[5] vssa1 0.61fF
C204 io_out[5] vssa1 0.61fF
C205 io_oeb[5] vssa1 0.61fF
C206 io_oeb[22] vssa1 0.61fF
C207 io_out[22] vssa1 0.61fF
C208 io_in[22] vssa1 0.61fF
C209 io_in_3v3[22] vssa1 0.61fF
C210 gpio_noesd[15] vssa1 0.61fF
C211 gpio_analog[15] vssa1 0.61fF
C212 io_in_3v3[6] vssa1 0.61fF
C213 io_in[6] vssa1 0.61fF
C214 io_out[6] vssa1 0.61fF
C215 io_oeb[6] vssa1 0.61fF
C216 io_oeb[21] vssa1 0.61fF
C217 io_out[21] vssa1 0.61fF
C218 io_in[21] vssa1 0.61fF
C219 io_in_3v3[21] vssa1 0.61fF
C220 gpio_noesd[14] vssa1 0.61fF
C221 gpio_analog[14] vssa1 0.61fF
C222 vssd2 vssa1 13.04fF
C223 vssd1 vssa1 13.04fF
C224 vdda2 vssa1 13.04fF
C225 vdda1 vssa1 26.08fF
C226 io_oeb[20] vssa1 0.61fF
C227 io_out[20] vssa1 0.61fF
C228 io_in[20] vssa1 0.61fF
C229 io_in_3v3[20] vssa1 0.61fF
C230 gpio_noesd[13] vssa1 0.61fF
C231 gpio_analog[13] vssa1 0.61fF
C232 gpio_analog[0] vssa1 0.61fF
C233 gpio_noesd[0] vssa1 0.61fF
C234 io_in_3v3[7] vssa1 0.61fF
C235 io_in[7] vssa1 0.61fF
C236 io_out[7] vssa1 0.61fF
C237 io_oeb[7] vssa1 0.61fF
C238 io_oeb[19] vssa1 0.61fF
C239 io_out[19] vssa1 0.61fF
C240 io_in[19] vssa1 0.61fF
C241 io_in_3v3[19] vssa1 0.61fF
C242 gpio_noesd[12] vssa1 0.61fF
C243 gpio_analog[12] vssa1 0.61fF
C244 gpio_analog[1] vssa1 0.61fF
C245 gpio_noesd[1] vssa1 0.61fF
C246 io_in_3v3[8] vssa1 0.61fF
C247 io_in[8] vssa1 0.61fF
C248 io_out[8] vssa1 0.61fF
C249 io_oeb[8] vssa1 0.61fF
C250 io_oeb[18] vssa1 0.61fF
C251 io_out[18] vssa1 0.61fF
C252 io_in[18] vssa1 0.61fF
C253 io_in_3v3[18] vssa1 0.61fF
C254 gpio_noesd[11] vssa1 0.61fF
C255 gpio_analog[11] vssa1 0.61fF
C256 gpio_analog[2] vssa1 0.61fF
C257 gpio_noesd[2] vssa1 0.61fF
C258 io_in_3v3[9] vssa1 0.61fF
C259 io_in[9] vssa1 0.61fF
C260 io_out[9] vssa1 0.61fF
C261 io_oeb[9] vssa1 0.61fF
C262 io_oeb[17] vssa1 0.61fF
C263 io_out[17] vssa1 0.61fF
C264 io_in[17] vssa1 0.61fF
C265 io_in_3v3[17] vssa1 0.61fF
C266 gpio_noesd[10] vssa1 0.61fF
C267 gpio_analog[10] vssa1 0.61fF
C268 gpio_analog[3] vssa1 0.61fF
C269 gpio_noesd[3] vssa1 0.61fF
C270 io_in_3v3[10] vssa1 0.61fF
C271 io_in[10] vssa1 0.61fF
C272 io_out[10] vssa1 0.61fF
C273 io_oeb[10] vssa1 0.61fF
C274 io_oeb[16] vssa1 0.61fF
C275 io_out[16] vssa1 0.61fF
C276 io_in[16] vssa1 0.61fF
C277 io_in_3v3[16] vssa1 0.61fF
C278 gpio_noesd[9] vssa1 0.61fF
C279 gpio_analog[9] vssa1 0.61fF
C280 gpio_analog[4] vssa1 0.61fF
C281 gpio_noesd[4] vssa1 0.61fF
C282 io_in_3v3[11] vssa1 0.61fF
C283 io_in[11] vssa1 0.61fF
C284 io_out[11] vssa1 0.61fF
C285 io_oeb[11] vssa1 0.61fF
C286 io_oeb[15] vssa1 0.61fF
C287 io_out[15] vssa1 0.61fF
C288 io_in[15] vssa1 0.61fF
C289 io_in_3v3[15] vssa1 0.61fF
C290 gpio_noesd[8] vssa1 0.61fF
C291 gpio_analog[8] vssa1 0.61fF
C292 gpio_analog[5] vssa1 0.61fF
C293 gpio_noesd[5] vssa1 0.61fF
C294 io_in_3v3[12] vssa1 0.61fF
C295 io_in[12] vssa1 0.61fF
C296 io_out[12] vssa1 0.61fF
C297 io_oeb[12] vssa1 0.61fF
C298 io_oeb[14] vssa1 0.61fF
C299 io_out[14] vssa1 0.61fF
C300 io_in[14] vssa1 0.61fF
C301 io_in_3v3[14] vssa1 0.61fF
C302 gpio_noesd[7] vssa1 0.61fF
C303 gpio_analog[7] vssa1 0.61fF
C304 vssa2 vssa1 13.04fF
C305 gpio_analog[6] vssa1 0.61fF
C306 gpio_noesd[6] vssa1 0.61fF
C307 io_in_3v3[13] vssa1 0.61fF
C308 io_in[13] vssa1 0.61fF
C309 io_out[13] vssa1 0.61fF
C310 io_oeb[13] vssa1 0.61fF
C311 vccd2 vssa1 13.04fF
C312 io_analog[0] vssa1 6.83fF
C313 io_analog[10] vssa1 6.83fF
C314 io_clamp_high[0] vssa1 4.88fF
C315 io_clamp_low[0] vssa1 4.88fF
C316 io_clamp_high[1] vssa1 4.74fF
C317 io_clamp_low[1] vssa1 4.74fF
C318 io_clamp_high[2] vssa1 4.90fF
C319 io_clamp_low[2] vssa1 4.91fF
C320 io_analog[8] vssa1 6.83fF
C321 io_analog[9] vssa1 6.83fF
C322 user_irq[2] vssa1 0.63fF
C323 user_irq[1] vssa1 0.63fF
C324 user_irq[0] vssa1 0.63fF
C325 user_clock2 vssa1 0.63fF
C326 la_oenb[127] vssa1 0.63fF
C327 la_data_out[127] vssa1 0.63fF
C328 la_data_in[127] vssa1 0.63fF
C329 la_oenb[126] vssa1 0.63fF
C330 la_data_out[126] vssa1 0.63fF
C331 la_data_in[126] vssa1 0.63fF
C332 la_oenb[125] vssa1 0.63fF
C333 la_data_out[125] vssa1 0.63fF
C334 la_data_in[125] vssa1 0.63fF
C335 la_oenb[124] vssa1 0.63fF
C336 la_data_out[124] vssa1 0.63fF
C337 la_data_in[124] vssa1 0.63fF
C338 la_oenb[123] vssa1 0.63fF
C339 la_data_out[123] vssa1 0.63fF
C340 la_data_in[123] vssa1 0.63fF
C341 la_oenb[122] vssa1 0.63fF
C342 la_data_out[122] vssa1 0.63fF
C343 la_data_in[122] vssa1 0.63fF
C344 la_oenb[121] vssa1 0.63fF
C345 la_data_out[121] vssa1 0.63fF
C346 la_data_in[121] vssa1 0.63fF
C347 la_oenb[120] vssa1 0.63fF
C348 la_data_out[120] vssa1 0.63fF
C349 la_data_in[120] vssa1 0.63fF
C350 la_oenb[119] vssa1 0.63fF
C351 la_data_out[119] vssa1 0.63fF
C352 la_data_in[119] vssa1 0.63fF
C353 la_oenb[118] vssa1 0.63fF
C354 la_data_out[118] vssa1 0.63fF
C355 la_data_in[118] vssa1 0.63fF
C356 la_oenb[117] vssa1 0.63fF
C357 la_data_out[117] vssa1 0.63fF
C358 la_data_in[117] vssa1 0.63fF
C359 la_oenb[116] vssa1 0.63fF
C360 la_data_out[116] vssa1 0.63fF
C361 la_data_in[116] vssa1 0.63fF
C362 la_oenb[115] vssa1 0.63fF
C363 la_data_out[115] vssa1 0.63fF
C364 la_data_in[115] vssa1 0.63fF
C365 la_oenb[114] vssa1 0.63fF
C366 la_data_out[114] vssa1 0.63fF
C367 la_data_in[114] vssa1 0.63fF
C368 la_oenb[113] vssa1 0.63fF
C369 la_data_out[113] vssa1 0.63fF
C370 la_data_in[113] vssa1 0.63fF
C371 la_oenb[112] vssa1 0.63fF
C372 la_data_out[112] vssa1 0.63fF
C373 la_data_in[112] vssa1 0.63fF
C374 la_oenb[111] vssa1 0.63fF
C375 la_data_out[111] vssa1 0.63fF
C376 la_data_in[111] vssa1 0.63fF
C377 la_oenb[110] vssa1 0.63fF
C378 la_data_out[110] vssa1 0.63fF
C379 la_data_in[110] vssa1 0.63fF
C380 la_oenb[109] vssa1 0.63fF
C381 la_data_out[109] vssa1 0.63fF
C382 la_data_in[109] vssa1 0.63fF
C383 la_oenb[108] vssa1 0.63fF
C384 la_data_out[108] vssa1 0.63fF
C385 la_data_in[108] vssa1 0.63fF
C386 la_oenb[107] vssa1 0.63fF
C387 la_data_out[107] vssa1 0.63fF
C388 la_data_in[107] vssa1 0.63fF
C389 la_oenb[106] vssa1 0.63fF
C390 la_data_out[106] vssa1 0.63fF
C391 la_data_in[106] vssa1 0.63fF
C392 la_oenb[105] vssa1 0.63fF
C393 la_data_out[105] vssa1 0.63fF
C394 la_data_in[105] vssa1 0.63fF
C395 la_oenb[104] vssa1 0.63fF
C396 la_data_out[104] vssa1 0.63fF
C397 la_data_in[104] vssa1 0.63fF
C398 la_oenb[103] vssa1 0.63fF
C399 la_data_out[103] vssa1 0.63fF
C400 la_data_in[103] vssa1 0.63fF
C401 la_oenb[102] vssa1 0.63fF
C402 la_data_out[102] vssa1 0.63fF
C403 la_data_in[102] vssa1 0.63fF
C404 la_oenb[101] vssa1 0.63fF
C405 la_data_out[101] vssa1 0.63fF
C406 la_data_in[101] vssa1 0.63fF
C407 la_oenb[100] vssa1 0.63fF
C408 la_data_out[100] vssa1 0.63fF
C409 la_data_in[100] vssa1 0.63fF
C410 la_oenb[99] vssa1 0.63fF
C411 la_data_out[99] vssa1 0.63fF
C412 la_data_in[99] vssa1 0.63fF
C413 la_oenb[98] vssa1 0.63fF
C414 la_data_out[98] vssa1 0.63fF
C415 la_data_in[98] vssa1 0.63fF
C416 la_oenb[97] vssa1 0.63fF
C417 la_data_out[97] vssa1 0.63fF
C418 la_data_in[97] vssa1 0.63fF
C419 la_oenb[96] vssa1 0.63fF
C420 la_data_out[96] vssa1 0.63fF
C421 la_data_in[96] vssa1 0.63fF
C422 la_oenb[95] vssa1 0.63fF
C423 la_data_out[95] vssa1 0.63fF
C424 la_data_in[95] vssa1 0.63fF
C425 la_oenb[94] vssa1 0.63fF
C426 la_data_out[94] vssa1 0.63fF
C427 la_data_in[94] vssa1 0.63fF
C428 la_oenb[93] vssa1 0.63fF
C429 la_data_out[93] vssa1 0.63fF
C430 la_data_in[93] vssa1 0.63fF
C431 la_oenb[92] vssa1 0.63fF
C432 la_data_out[92] vssa1 0.63fF
C433 la_data_in[92] vssa1 0.63fF
C434 la_oenb[91] vssa1 0.63fF
C435 la_data_out[91] vssa1 0.63fF
C436 la_data_in[91] vssa1 0.63fF
C437 la_oenb[90] vssa1 0.63fF
C438 la_data_out[90] vssa1 0.63fF
C439 la_data_in[90] vssa1 0.63fF
C440 la_oenb[89] vssa1 0.63fF
C441 la_data_out[89] vssa1 0.63fF
C442 la_data_in[89] vssa1 0.63fF
C443 la_oenb[88] vssa1 0.63fF
C444 la_data_out[88] vssa1 0.63fF
C445 la_data_in[88] vssa1 0.63fF
C446 la_oenb[87] vssa1 0.63fF
C447 la_data_out[87] vssa1 0.63fF
C448 la_data_in[87] vssa1 0.63fF
C449 la_oenb[86] vssa1 0.63fF
C450 la_data_out[86] vssa1 0.63fF
C451 la_data_in[86] vssa1 0.63fF
C452 la_oenb[85] vssa1 0.63fF
C453 la_data_out[85] vssa1 0.63fF
C454 la_data_in[85] vssa1 0.63fF
C455 la_oenb[84] vssa1 0.63fF
C456 la_data_out[84] vssa1 0.63fF
C457 la_data_in[84] vssa1 0.63fF
C458 la_oenb[83] vssa1 0.63fF
C459 la_data_out[83] vssa1 0.63fF
C460 la_data_in[83] vssa1 0.63fF
C461 la_oenb[82] vssa1 0.63fF
C462 la_data_out[82] vssa1 0.63fF
C463 la_data_in[82] vssa1 0.63fF
C464 la_oenb[81] vssa1 0.63fF
C465 la_data_out[81] vssa1 0.63fF
C466 la_data_in[81] vssa1 0.63fF
C467 la_oenb[80] vssa1 0.63fF
C468 la_data_out[80] vssa1 0.63fF
C469 la_data_in[80] vssa1 0.63fF
C470 la_oenb[79] vssa1 0.63fF
C471 la_data_out[79] vssa1 0.63fF
C472 la_data_in[79] vssa1 0.63fF
C473 la_oenb[78] vssa1 0.63fF
C474 la_data_out[78] vssa1 0.63fF
C475 la_data_in[78] vssa1 0.63fF
C476 la_oenb[77] vssa1 0.63fF
C477 la_data_out[77] vssa1 0.63fF
C478 la_data_in[77] vssa1 0.63fF
C479 la_oenb[76] vssa1 0.63fF
C480 la_data_out[76] vssa1 0.63fF
C481 la_data_in[76] vssa1 0.63fF
C482 la_oenb[75] vssa1 0.63fF
C483 la_data_out[75] vssa1 0.63fF
C484 la_data_in[75] vssa1 0.63fF
C485 la_oenb[74] vssa1 0.63fF
C486 la_data_out[74] vssa1 0.63fF
C487 la_data_in[74] vssa1 0.63fF
C488 la_oenb[73] vssa1 0.63fF
C489 la_data_out[73] vssa1 0.63fF
C490 la_data_in[73] vssa1 0.63fF
C491 la_oenb[72] vssa1 0.63fF
C492 la_data_out[72] vssa1 0.63fF
C493 la_data_in[72] vssa1 0.63fF
C494 la_oenb[71] vssa1 0.63fF
C495 la_data_out[71] vssa1 0.63fF
C496 la_data_in[71] vssa1 0.63fF
C497 la_oenb[70] vssa1 0.63fF
C498 la_data_out[70] vssa1 0.63fF
C499 la_data_in[70] vssa1 0.63fF
C500 la_oenb[69] vssa1 0.63fF
C501 la_data_out[69] vssa1 0.63fF
C502 la_data_in[69] vssa1 0.63fF
C503 la_oenb[68] vssa1 0.63fF
C504 la_data_out[68] vssa1 0.63fF
C505 la_data_in[68] vssa1 0.63fF
C506 la_oenb[67] vssa1 0.63fF
C507 la_data_out[67] vssa1 0.63fF
C508 la_data_in[67] vssa1 0.63fF
C509 la_oenb[66] vssa1 0.63fF
C510 la_data_out[66] vssa1 0.63fF
C511 la_data_in[66] vssa1 0.63fF
C512 la_oenb[65] vssa1 0.63fF
C513 la_data_out[65] vssa1 0.63fF
C514 la_data_in[65] vssa1 0.63fF
C515 la_oenb[64] vssa1 0.63fF
C516 la_data_out[64] vssa1 0.63fF
C517 la_data_in[64] vssa1 0.63fF
C518 la_oenb[63] vssa1 0.63fF
C519 la_data_out[63] vssa1 0.63fF
C520 la_data_in[63] vssa1 0.63fF
C521 la_oenb[62] vssa1 0.63fF
C522 la_data_out[62] vssa1 0.63fF
C523 la_data_in[62] vssa1 0.63fF
C524 la_oenb[61] vssa1 0.63fF
C525 la_data_out[61] vssa1 0.63fF
C526 la_data_in[61] vssa1 0.63fF
C527 la_oenb[60] vssa1 0.63fF
C528 la_data_out[60] vssa1 0.63fF
C529 la_data_in[60] vssa1 0.63fF
C530 la_oenb[59] vssa1 0.63fF
C531 la_data_out[59] vssa1 0.63fF
C532 la_data_in[59] vssa1 0.63fF
C533 la_oenb[58] vssa1 0.63fF
C534 la_data_out[58] vssa1 0.63fF
C535 la_data_in[58] vssa1 0.63fF
C536 la_oenb[57] vssa1 0.63fF
C537 la_data_out[57] vssa1 0.63fF
C538 la_data_in[57] vssa1 0.63fF
C539 la_oenb[56] vssa1 0.63fF
C540 la_data_out[56] vssa1 0.63fF
C541 la_data_in[56] vssa1 0.63fF
C542 la_oenb[55] vssa1 0.63fF
C543 la_data_out[55] vssa1 0.63fF
C544 la_data_in[55] vssa1 0.63fF
C545 la_oenb[54] vssa1 0.63fF
C546 la_data_out[54] vssa1 0.63fF
C547 la_data_in[54] vssa1 0.63fF
C548 la_oenb[53] vssa1 0.63fF
C549 la_data_out[53] vssa1 0.63fF
C550 la_data_in[53] vssa1 0.63fF
C551 la_oenb[52] vssa1 0.63fF
C552 la_data_out[52] vssa1 0.63fF
C553 la_data_in[52] vssa1 0.63fF
C554 la_oenb[51] vssa1 0.63fF
C555 la_data_out[51] vssa1 0.63fF
C556 la_data_in[51] vssa1 0.63fF
C557 la_oenb[50] vssa1 0.63fF
C558 la_data_out[50] vssa1 0.63fF
C559 la_data_in[50] vssa1 0.63fF
C560 la_oenb[49] vssa1 0.63fF
C561 la_data_out[49] vssa1 0.63fF
C562 la_data_in[49] vssa1 0.63fF
C563 la_oenb[48] vssa1 0.63fF
C564 la_data_out[48] vssa1 0.63fF
C565 la_data_in[48] vssa1 0.63fF
C566 la_oenb[47] vssa1 0.63fF
C567 la_data_out[47] vssa1 0.63fF
C568 la_data_in[47] vssa1 0.63fF
C569 la_oenb[46] vssa1 0.63fF
C570 la_data_out[46] vssa1 0.63fF
C571 la_data_in[46] vssa1 0.63fF
C572 la_oenb[45] vssa1 0.63fF
C573 la_data_out[45] vssa1 0.63fF
C574 la_data_in[45] vssa1 0.63fF
C575 la_oenb[44] vssa1 0.63fF
C576 la_data_out[44] vssa1 0.63fF
C577 la_data_in[44] vssa1 0.63fF
C578 la_oenb[43] vssa1 0.63fF
C579 la_data_out[43] vssa1 0.63fF
C580 la_data_in[43] vssa1 0.63fF
C581 la_oenb[42] vssa1 0.63fF
C582 la_data_out[42] vssa1 0.63fF
C583 la_data_in[42] vssa1 0.63fF
C584 la_oenb[41] vssa1 0.63fF
C585 la_data_out[41] vssa1 0.63fF
C586 la_data_in[41] vssa1 0.63fF
C587 la_oenb[40] vssa1 0.63fF
C588 la_data_out[40] vssa1 0.63fF
C589 la_data_in[40] vssa1 0.63fF
C590 la_oenb[39] vssa1 0.63fF
C591 la_data_out[39] vssa1 0.63fF
C592 la_data_in[39] vssa1 0.63fF
C593 la_oenb[38] vssa1 0.63fF
C594 la_data_out[38] vssa1 0.63fF
C595 la_data_in[38] vssa1 0.63fF
C596 la_oenb[37] vssa1 0.63fF
C597 la_data_out[37] vssa1 0.63fF
C598 la_data_in[37] vssa1 0.63fF
C599 la_oenb[36] vssa1 0.63fF
C600 la_data_out[36] vssa1 0.63fF
C601 la_data_in[36] vssa1 0.63fF
C602 la_oenb[35] vssa1 0.63fF
C603 la_data_out[35] vssa1 0.63fF
C604 la_data_in[35] vssa1 0.63fF
C605 la_oenb[34] vssa1 0.63fF
C606 la_data_out[34] vssa1 0.63fF
C607 la_data_in[34] vssa1 0.63fF
C608 la_oenb[33] vssa1 0.63fF
C609 la_data_out[33] vssa1 0.63fF
C610 la_data_in[33] vssa1 0.63fF
C611 la_oenb[32] vssa1 0.63fF
C612 la_data_out[32] vssa1 0.63fF
C613 la_data_in[32] vssa1 0.63fF
C614 la_oenb[31] vssa1 0.63fF
C615 la_data_out[31] vssa1 0.63fF
C616 la_data_in[31] vssa1 0.63fF
C617 la_oenb[30] vssa1 0.63fF
C618 la_data_out[30] vssa1 0.63fF
C619 la_data_in[30] vssa1 0.63fF
C620 la_oenb[29] vssa1 0.63fF
C621 la_data_out[29] vssa1 0.63fF
C622 la_data_in[29] vssa1 0.63fF
C623 la_oenb[28] vssa1 0.63fF
C624 la_data_out[28] vssa1 0.63fF
C625 la_data_in[28] vssa1 0.63fF
C626 la_oenb[27] vssa1 0.63fF
C627 la_data_out[27] vssa1 0.63fF
C628 la_data_in[27] vssa1 0.63fF
C629 la_oenb[26] vssa1 0.63fF
C630 la_data_out[26] vssa1 0.63fF
C631 la_data_in[26] vssa1 0.63fF
C632 la_oenb[25] vssa1 0.63fF
C633 la_data_out[25] vssa1 0.63fF
C634 la_data_in[25] vssa1 0.63fF
C635 la_oenb[24] vssa1 0.63fF
C636 la_data_out[24] vssa1 0.63fF
C637 la_data_in[24] vssa1 0.63fF
C638 la_oenb[23] vssa1 0.63fF
C639 la_data_out[23] vssa1 0.63fF
C640 la_data_in[23] vssa1 0.63fF
C641 la_oenb[22] vssa1 0.63fF
C642 la_data_out[22] vssa1 0.63fF
C643 la_data_in[22] vssa1 0.63fF
C644 la_oenb[21] vssa1 0.63fF
C645 la_data_out[21] vssa1 0.63fF
C646 la_data_in[21] vssa1 0.63fF
C647 la_oenb[20] vssa1 0.63fF
C648 la_data_out[20] vssa1 0.63fF
C649 la_data_in[20] vssa1 0.63fF
C650 la_oenb[19] vssa1 0.63fF
C651 la_data_out[19] vssa1 0.63fF
C652 la_data_in[19] vssa1 0.63fF
C653 la_oenb[18] vssa1 0.63fF
C654 la_data_out[18] vssa1 0.63fF
C655 la_data_in[18] vssa1 0.63fF
C656 la_oenb[17] vssa1 0.63fF
C657 la_data_out[17] vssa1 0.63fF
C658 la_data_in[17] vssa1 0.63fF
C659 la_oenb[16] vssa1 0.63fF
C660 la_data_out[16] vssa1 0.63fF
C661 la_data_in[16] vssa1 0.63fF
C662 la_oenb[15] vssa1 0.63fF
C663 la_data_out[15] vssa1 0.63fF
C664 la_data_in[15] vssa1 0.63fF
C665 la_oenb[14] vssa1 0.63fF
C666 la_data_out[14] vssa1 0.63fF
C667 la_data_in[14] vssa1 0.63fF
C668 la_oenb[13] vssa1 0.63fF
C669 la_data_out[13] vssa1 0.63fF
C670 la_data_in[13] vssa1 0.63fF
C671 la_oenb[12] vssa1 0.63fF
C672 la_data_out[12] vssa1 0.63fF
C673 la_data_in[12] vssa1 0.63fF
C674 la_oenb[11] vssa1 0.63fF
C675 la_data_out[11] vssa1 0.63fF
C676 la_data_in[11] vssa1 0.63fF
C677 la_oenb[10] vssa1 0.63fF
C678 la_data_out[10] vssa1 0.63fF
C679 la_data_in[10] vssa1 0.63fF
C680 la_oenb[9] vssa1 0.63fF
C681 la_data_out[9] vssa1 0.63fF
C682 la_data_in[9] vssa1 0.63fF
C683 la_oenb[8] vssa1 0.63fF
C684 la_data_out[8] vssa1 0.63fF
C685 la_data_in[8] vssa1 0.63fF
C686 la_oenb[7] vssa1 0.63fF
C687 la_data_out[7] vssa1 0.63fF
C688 la_data_in[7] vssa1 0.63fF
C689 la_oenb[6] vssa1 0.63fF
C690 la_data_out[6] vssa1 0.63fF
C691 la_data_in[6] vssa1 0.63fF
C692 la_oenb[5] vssa1 0.63fF
C693 la_data_out[5] vssa1 0.63fF
C694 la_data_in[5] vssa1 0.63fF
C695 la_oenb[4] vssa1 0.63fF
C696 la_data_out[4] vssa1 0.63fF
C697 la_data_in[4] vssa1 0.63fF
C698 la_oenb[3] vssa1 0.63fF
C699 la_data_out[3] vssa1 0.63fF
C700 la_data_in[3] vssa1 0.63fF
C701 la_oenb[2] vssa1 0.63fF
C702 la_data_out[2] vssa1 0.63fF
C703 la_data_in[2] vssa1 0.63fF
C704 la_oenb[1] vssa1 0.63fF
C705 la_data_out[1] vssa1 0.63fF
C706 la_data_in[1] vssa1 0.63fF
C707 la_oenb[0] vssa1 0.63fF
C708 la_data_out[0] vssa1 0.63fF
C709 la_data_in[0] vssa1 0.63fF
C710 wbs_dat_o[31] vssa1 0.63fF
C711 wbs_dat_i[31] vssa1 0.63fF
C712 wbs_adr_i[31] vssa1 0.63fF
C713 wbs_dat_o[30] vssa1 0.63fF
C714 wbs_dat_i[30] vssa1 0.63fF
C715 wbs_adr_i[30] vssa1 0.63fF
C716 wbs_dat_o[29] vssa1 0.63fF
C717 wbs_dat_i[29] vssa1 0.63fF
C718 wbs_adr_i[29] vssa1 0.63fF
C719 wbs_dat_o[28] vssa1 0.63fF
C720 wbs_dat_i[28] vssa1 0.63fF
C721 wbs_adr_i[28] vssa1 0.63fF
C722 wbs_dat_o[27] vssa1 0.63fF
C723 wbs_dat_i[27] vssa1 0.63fF
C724 wbs_adr_i[27] vssa1 0.63fF
C725 wbs_dat_o[26] vssa1 0.63fF
C726 wbs_dat_i[26] vssa1 0.63fF
C727 wbs_adr_i[26] vssa1 0.63fF
C728 wbs_dat_o[25] vssa1 0.63fF
C729 wbs_dat_i[25] vssa1 0.63fF
C730 wbs_adr_i[25] vssa1 0.63fF
C731 wbs_dat_o[24] vssa1 0.63fF
C732 wbs_dat_i[24] vssa1 0.63fF
C733 wbs_adr_i[24] vssa1 0.63fF
C734 wbs_dat_o[23] vssa1 0.63fF
C735 wbs_dat_i[23] vssa1 0.63fF
C736 wbs_adr_i[23] vssa1 0.63fF
C737 wbs_dat_o[22] vssa1 0.63fF
C738 wbs_dat_i[22] vssa1 0.63fF
C739 wbs_adr_i[22] vssa1 0.63fF
C740 wbs_dat_o[21] vssa1 0.63fF
C741 wbs_dat_i[21] vssa1 0.63fF
C742 wbs_adr_i[21] vssa1 0.63fF
C743 wbs_dat_o[20] vssa1 0.63fF
C744 wbs_dat_i[20] vssa1 0.63fF
C745 wbs_adr_i[20] vssa1 0.63fF
C746 wbs_dat_o[19] vssa1 0.63fF
C747 wbs_dat_i[19] vssa1 0.63fF
C748 wbs_adr_i[19] vssa1 0.63fF
C749 wbs_dat_o[18] vssa1 0.63fF
C750 wbs_dat_i[18] vssa1 0.63fF
C751 wbs_adr_i[18] vssa1 0.63fF
C752 wbs_dat_o[17] vssa1 0.63fF
C753 wbs_dat_i[17] vssa1 0.63fF
C754 wbs_adr_i[17] vssa1 0.63fF
C755 wbs_dat_o[16] vssa1 0.63fF
C756 wbs_dat_i[16] vssa1 0.63fF
C757 wbs_adr_i[16] vssa1 0.63fF
C758 wbs_dat_o[15] vssa1 0.63fF
C759 wbs_dat_i[15] vssa1 0.63fF
C760 wbs_adr_i[15] vssa1 0.63fF
C761 wbs_dat_o[14] vssa1 0.63fF
C762 wbs_dat_i[14] vssa1 0.63fF
C763 wbs_adr_i[14] vssa1 0.63fF
C764 wbs_dat_o[13] vssa1 0.63fF
C765 wbs_dat_i[13] vssa1 0.63fF
C766 wbs_adr_i[13] vssa1 0.63fF
C767 wbs_dat_o[12] vssa1 0.63fF
C768 wbs_dat_i[12] vssa1 0.63fF
C769 wbs_adr_i[12] vssa1 0.63fF
C770 wbs_dat_o[11] vssa1 0.63fF
C771 wbs_dat_i[11] vssa1 0.63fF
C772 wbs_adr_i[11] vssa1 0.63fF
C773 wbs_dat_o[10] vssa1 0.63fF
C774 wbs_dat_i[10] vssa1 0.63fF
C775 wbs_adr_i[10] vssa1 0.63fF
C776 wbs_dat_o[9] vssa1 0.63fF
C777 wbs_dat_i[9] vssa1 0.63fF
C778 wbs_adr_i[9] vssa1 0.63fF
C779 wbs_dat_o[8] vssa1 0.63fF
C780 wbs_dat_i[8] vssa1 0.63fF
C781 wbs_adr_i[8] vssa1 0.63fF
C782 wbs_dat_o[7] vssa1 0.63fF
C783 wbs_dat_i[7] vssa1 0.63fF
C784 wbs_adr_i[7] vssa1 0.63fF
C785 wbs_dat_o[6] vssa1 0.63fF
C786 wbs_dat_i[6] vssa1 0.63fF
C787 wbs_adr_i[6] vssa1 0.63fF
C788 wbs_dat_o[5] vssa1 0.63fF
C789 wbs_dat_i[5] vssa1 0.63fF
C790 wbs_adr_i[5] vssa1 0.63fF
C791 wbs_dat_o[4] vssa1 0.63fF
C792 wbs_dat_i[4] vssa1 0.63fF
C793 wbs_adr_i[4] vssa1 0.63fF
C794 wbs_sel_i[3] vssa1 0.63fF
C795 wbs_dat_o[3] vssa1 0.63fF
C796 wbs_dat_i[3] vssa1 0.63fF
C797 wbs_adr_i[3] vssa1 0.63fF
C798 wbs_sel_i[2] vssa1 0.63fF
C799 wbs_dat_o[2] vssa1 0.63fF
C800 wbs_dat_i[2] vssa1 0.63fF
C801 wbs_adr_i[2] vssa1 0.63fF
C802 wbs_sel_i[1] vssa1 0.63fF
C803 wbs_dat_o[1] vssa1 0.63fF
C804 wbs_dat_i[1] vssa1 0.63fF
C805 wbs_adr_i[1] vssa1 0.63fF
C806 wbs_sel_i[0] vssa1 0.63fF
C807 wbs_dat_o[0] vssa1 0.63fF
C808 wbs_dat_i[0] vssa1 0.63fF
C809 wbs_adr_i[0] vssa1 0.63fF
C810 wbs_we_i vssa1 0.63fF
C811 wbs_stb_i vssa1 0.63fF
C812 wbs_cyc_i vssa1 0.63fF
C813 wbs_ack_o vssa1 0.63fF
C814 wb_rst_i vssa1 0.63fF
C815 wb_clk_i vssa1 0.63fF
C816 m3_326806_700392# vssa1 0.27fF $ **FLOATING
C817 m3_324320_700392# vssa1 0.27fF $ **FLOATING
C818 m3_225118_700522# vssa1 0.27fF $ **FLOATING
C819 m3_222608_700522# vssa1 0.27fF $ **FLOATING
C820 m3_173410_700370# vssa1 0.27fF $ **FLOATING
C821 m3_170914_700368# vssa1 0.27fF $ **FLOATING
C822 a_493938_644874# vssa1 43.58fF
C823 a_490782_644900# vssa1 42.98fF
C824 a_487694_644902# vssa1 43.39fF
C825 a_484664_644902# vssa1 43.98fF
C826 a_481708_644918# vssa1 44.10fF
C827 a_479772_646886# vssa1 35.70fF
C828 a_506614_647168# vssa1 33.83fF
C829 a_505416_647172# vssa1 22.63fF
C830 a_504724_647182# vssa1 12.41fF
C831 a_500126_647170# vssa1 33.86fF
C832 a_498928_647174# vssa1 22.60fF
C833 a_498236_647184# vssa1 12.39fF
C834 a_483446_644892# vssa1 21.83fF
C835 VCO_Flat_0/Buff_VCO_0/IN vssa1 12.42fF
C836 VCO_Flat_0/Buff_VCO_1/IN vssa1 16.05fF
C837 a_475058_648060# vssa1 12.40fF
C838 a_473374_648060# vssa1 22.58fF
C839 a_471230_648050# vssa1 33.87fF
C840 VCO_Flat_0/Buff_VCO_3/IN vssa1 18.42fF
C841 a_468592_648062# vssa1 12.39fF
C842 a_466908_648062# vssa1 22.59fF
C843 a_464764_648054# vssa1 33.85fF
C844 VCO_Flat_0/Buff_VCO_4/IN vssa1 15.80fF
C845 a_461762_648050# vssa1 12.39fF
C846 a_460078_648050# vssa1 22.61fF
C847 a_457934_648038# vssa1 33.90fF
C848 VCO_Flat_0/Buff_VCO_2/IN vssa1 13.45fF
C849 a_493974_650212# vssa1 2.48fF
C850 a_490818_650238# vssa1 2.48fF
C851 a_487730_650240# vssa1 2.48fF
C852 a_484700_650240# vssa1 2.48fF
C853 a_481744_650256# vssa1 2.47fF
C854 a_479864_646886# vssa1 15.32fF
C855 esd_1/in vssa1 171.63fF
C856 io_analog[1] vssa1 47.87fF
C857 esd_2/in vssa1 246.98fF
C858 io_analog[2] vssa1 47.79fF
C859 esd_3/in vssa1 147.76fF
C860 io_analog[3] vssa1 47.61fF
C861 esd_4/in vssa1 228.91fF
C862 io_analog[4] vssa1 62.55fF
C863 esd_5/in vssa1 337.52fF
C864 io_analog[5] vssa1 62.55fF
C865 esd_0/in vssa1 421.01fF
C866 io_analog[6] vssa1 62.80fF
C867 esd_6/in vssa1 484.76fF
C868 io_analog[7] vssa1 47.62fF
C869 vccd1 vssa1 2520.64fF
.ends

