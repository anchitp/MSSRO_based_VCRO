magic
tech sky130A
magscale 1 2
timestamp 1636295761
<< error_p >>
rect -705 536 -617 562
rect -705 528 701 536
rect 785 528 869 562
rect -741 492 737 500
rect -907 -392 -785 -358
rect -907 -492 -373 -392
rect -907 -500 749 -492
rect -907 -526 -373 -500
rect -785 -528 -373 -526
rect -785 -536 743 -528
rect -785 -600 -459 -536
rect 785 -600 911 -360
rect -739 -646 -627 -600
rect -701 -667 -643 -661
rect -701 -701 -689 -667
rect -701 -707 -643 -701
rect -627 -720 -571 -646
<< nwell >>
rect -785 528 -705 562
rect 701 528 785 562
rect -785 -526 785 528
rect -785 -600 -739 -526
rect -627 -528 785 -526
rect -627 -600 -561 -528
rect 743 -600 785 -528
rect -739 -720 -627 -646
<< pmos >>
rect -687 -500 -657 500
rect -591 -500 -561 500
rect -495 -500 -465 500
rect -399 -500 -369 500
rect -303 -500 -273 500
rect -207 -500 -177 500
rect -111 -500 -81 500
rect -15 -500 15 500
rect 81 -500 111 500
rect 177 -500 207 500
rect 273 -500 303 500
rect 369 -500 399 500
rect 465 -500 495 500
rect 561 -500 591 500
rect 657 -500 687 500
<< pdiff >>
rect -749 488 -687 500
rect -749 -488 -737 488
rect -703 -488 -687 488
rect -749 -500 -687 -488
rect -657 488 -591 500
rect -657 -488 -641 488
rect -607 -488 -591 488
rect -657 -500 -591 -488
rect -561 488 -495 500
rect -561 -488 -545 488
rect -511 -488 -495 488
rect -561 -500 -495 -488
rect -465 488 -399 500
rect -465 -488 -449 488
rect -415 -488 -399 488
rect -465 -500 -399 -488
rect -369 488 -303 500
rect -369 -488 -353 488
rect -319 -488 -303 488
rect -369 -500 -303 -488
rect -273 488 -207 500
rect -273 -488 -257 488
rect -223 -488 -207 488
rect -273 -500 -207 -488
rect -177 488 -111 500
rect -177 -488 -161 488
rect -127 -488 -111 488
rect -177 -500 -111 -488
rect -81 488 -15 500
rect -81 -488 -65 488
rect -31 -488 -15 488
rect -81 -500 -15 -488
rect 15 488 81 500
rect 15 -488 31 488
rect 65 -488 81 488
rect 15 -500 81 -488
rect 111 488 177 500
rect 111 -488 127 488
rect 161 -488 177 488
rect 111 -500 177 -488
rect 207 488 273 500
rect 207 -488 223 488
rect 257 -488 273 488
rect 207 -500 273 -488
rect 303 488 369 500
rect 303 -488 319 488
rect 353 -488 369 488
rect 303 -500 369 -488
rect 399 488 465 500
rect 399 -488 415 488
rect 449 -488 465 488
rect 399 -500 465 -488
rect 495 488 561 500
rect 495 -488 511 488
rect 545 -488 561 488
rect 495 -500 561 -488
rect 591 488 657 500
rect 591 -488 607 488
rect 641 -488 657 488
rect 591 -500 657 -488
rect 687 488 749 500
rect 687 -488 703 488
rect 737 -488 749 488
rect 687 -500 749 -488
<< pdiffc >>
rect -737 -488 -703 488
rect -641 -488 -607 488
rect -545 -488 -511 488
rect -449 -488 -415 488
rect -353 -488 -319 488
rect -257 -488 -223 488
rect -161 -488 -127 488
rect -65 -488 -31 488
rect 31 -488 65 488
rect 127 -488 161 488
rect 223 -488 257 488
rect 319 -488 353 488
rect 415 -488 449 488
rect 511 -488 545 488
rect 607 -488 641 488
rect 703 -488 737 488
<< poly >>
rect -687 500 -657 526
rect -591 500 -561 528
rect -495 500 -465 526
rect -399 500 -369 528
rect -303 500 -273 526
rect -207 500 -177 528
rect -111 500 -81 526
rect -15 500 15 528
rect 81 500 111 526
rect 177 500 207 528
rect 273 500 303 526
rect 369 500 399 528
rect 465 500 495 526
rect 561 500 591 528
rect 657 500 687 526
rect -687 -518 -657 -500
rect -591 -518 -561 -500
rect -495 -518 -465 -500
rect -399 -518 -369 -500
rect -303 -518 -273 -500
rect -207 -518 -177 -500
rect -111 -518 -81 -500
rect -15 -518 15 -500
rect 81 -518 111 -500
rect 177 -518 207 -500
rect 273 -518 303 -500
rect 369 -518 399 -500
rect 465 -518 495 -500
rect 561 -518 591 -500
rect 657 -518 687 -500
rect -687 -548 687 -518
rect -687 -651 -657 -548
rect -705 -667 -639 -651
rect -705 -701 -689 -667
rect -655 -701 -639 -667
rect -705 -717 -639 -701
<< polycont >>
rect -689 -701 -655 -667
<< locali >>
rect -737 546 641 580
rect -737 488 -703 546
rect -737 -504 -703 -488
rect -641 488 -607 504
rect -641 -562 -607 -488
rect -545 488 -511 546
rect -545 -504 -511 -488
rect -449 488 -415 504
rect -449 -562 -415 -488
rect -353 488 -319 546
rect -353 -504 -319 -488
rect -257 488 -223 504
rect -257 -562 -223 -488
rect -161 488 -127 546
rect -161 -504 -127 -488
rect -65 488 -31 504
rect -65 -562 -31 -488
rect 31 488 65 546
rect 31 -504 65 -488
rect 127 488 161 504
rect 127 -562 161 -488
rect 223 488 257 546
rect 223 -504 257 -488
rect 319 488 353 504
rect 319 -562 353 -488
rect 415 488 449 546
rect 415 -504 449 -488
rect 511 488 545 504
rect 511 -562 545 -488
rect 607 488 641 546
rect 607 -504 641 -488
rect 703 488 737 504
rect 703 -562 737 -488
rect -641 -596 737 -562
rect -705 -701 -689 -667
rect -655 -701 -639 -667
<< viali >>
rect -737 -488 -703 488
rect -641 -488 -607 488
rect -545 -488 -511 488
rect -449 -488 -415 488
rect -353 -488 -319 488
rect -257 -488 -223 488
rect -161 -488 -127 488
rect -65 -488 -31 488
rect 31 -488 65 488
rect 127 -488 161 488
rect 223 -488 257 488
rect 319 -488 353 488
rect 415 -488 449 488
rect 511 -488 545 488
rect 607 -488 641 488
rect 703 -488 737 488
rect -689 -701 -655 -667
<< metal1 >>
rect -743 488 -697 500
rect -743 -488 -737 488
rect -703 -488 -697 488
rect -743 -500 -697 -488
rect -647 488 -601 500
rect -647 -488 -641 488
rect -607 -488 -601 488
rect -647 -500 -601 -488
rect -551 488 -505 500
rect -551 -488 -545 488
rect -511 -488 -505 488
rect -551 -500 -505 -488
rect -455 488 -409 500
rect -455 -488 -449 488
rect -415 -488 -409 488
rect -455 -500 -409 -488
rect -359 488 -313 500
rect -359 -488 -353 488
rect -319 -488 -313 488
rect -359 -500 -313 -488
rect -263 488 -217 500
rect -263 -488 -257 488
rect -223 -488 -217 488
rect -263 -500 -217 -488
rect -167 488 -121 500
rect -167 -488 -161 488
rect -127 -488 -121 488
rect -167 -500 -121 -488
rect -71 488 -25 500
rect -71 -488 -65 488
rect -31 -488 -25 488
rect -71 -500 -25 -488
rect 25 488 71 500
rect 25 -488 31 488
rect 65 -488 71 488
rect 25 -500 71 -488
rect 121 488 167 500
rect 121 -488 127 488
rect 161 -488 167 488
rect 121 -500 167 -488
rect 217 488 263 500
rect 217 -488 223 488
rect 257 -488 263 488
rect 217 -500 263 -488
rect 313 488 359 500
rect 313 -488 319 488
rect 353 -488 359 488
rect 313 -500 359 -488
rect 409 488 455 500
rect 409 -488 415 488
rect 449 -488 455 488
rect 409 -500 455 -488
rect 505 488 551 500
rect 505 -488 511 488
rect 545 -488 551 488
rect 505 -500 551 -488
rect 601 488 647 500
rect 601 -488 607 488
rect 641 -488 647 488
rect 601 -500 647 -488
rect 697 488 743 500
rect 697 -488 703 488
rect 737 -488 743 488
rect 697 -500 743 -488
rect -701 -667 -643 -661
rect -701 -701 -689 -667
rect -655 -701 -643 -667
rect -701 -707 -643 -701
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string parameters w 5 l 0.15 m 1 nf 15 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
